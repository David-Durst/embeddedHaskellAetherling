// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  output [7:0] O
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x205_TREADY(dontcare), // @[:@1298.4]
    .io_in_x205_TDATA(I_0), // @[:@1298.4]
    .io_in_x205_TID(8'h0),
    .io_in_x205_TDEST(8'h0),
    .io_in_x206_TVALID(valid_down), // @[:@1298.4]
    .io_in_x206_TDATA(O), // @[:@1298.4]
    .io_in_x206_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x213_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh3e); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh3e); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 284:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x326_outr_UnitPipe_sm( // @[:@2390.2]
  input   clock, // @[:@2391.4]
  input   reset, // @[:@2392.4]
  input   io_enable, // @[:@2393.4]
  output  io_done, // @[:@2393.4]
  input   io_parentAck, // @[:@2393.4]
  input   io_doneIn_0, // @[:@2393.4]
  output  io_enableOut_0, // @[:@2393.4]
  output  io_childAck_0, // @[:@2393.4]
  input   io_ctrCopyDone_0 // @[:@2393.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2396.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2399.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2416.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2533.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2431.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2432.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2433.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2434.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2435.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2438.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2440.4]
  wire  _T_126; // @[package.scala 96:25:@2452.4 package.scala 96:25:@2453.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2455.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2456.4]
  wire  _T_138; // @[package.scala 96:25:@2466.4 package.scala 96:25:@2467.4]
  wire  _T_156; // @[package.scala 96:25:@2484.4 package.scala 96:25:@2485.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2487.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2488.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2502.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2504.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2506.4]
  reg  _T_186; // @[package.scala 48:56:@2512.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2514.4]
  reg  _T_200; // @[package.scala 48:56:@2530.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2396.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2399.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2416.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2447.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2461.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2479.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2516.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2533.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2431.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2432.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2433.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2434.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2435.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2438.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2440.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2452.4 package.scala 96:25:@2453.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2455.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2456.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2466.4 package.scala 96:25:@2467.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2484.4 package.scala 96:25:@2485.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2487.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2488.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2502.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2504.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2506.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2514.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2540.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2510.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2501.4]
  assign active_0_clock = clock; // @[:@2397.4]
  assign active_0_reset = reset; // @[:@2398.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2442.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2446.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2404.4]
  assign done_0_clock = clock; // @[:@2400.4]
  assign done_0_reset = reset; // @[:@2401.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2492.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2414.4 Controllers.scala 170:32:@2499.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2405.4]
  assign iterDone_0_clock = clock; // @[:@2417.4]
  assign iterDone_0_reset = reset; // @[:@2418.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2460.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2428.4 Controllers.scala 168:36:@2476.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2419.4]
  assign RetimeWrapper_clock = clock; // @[:@2448.4]
  assign RetimeWrapper_reset = reset; // @[:@2449.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2451.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2450.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2462.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2463.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2465.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2464.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2480.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2481.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2483.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2482.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2517.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2518.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2520.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2519.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2534.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2535.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2537.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2536.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2661.2]
  input         clock, // @[:@2662.4]
  input         reset, // @[:@2663.4]
  input         io_input_reset, // @[:@2664.4]
  input         io_input_enable, // @[:@2664.4]
  output [12:0] io_output_count_0, // @[:@2664.4]
  output        io_output_oobs_0, // @[:@2664.4]
  output        io_output_done, // @[:@2664.4]
  output        io_output_saturated // @[:@2664.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@2677.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@2677.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@2677.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@2693.4]
  wire  _T_36; // @[Counter.scala 264:45:@2696.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@2721.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@2722.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@2723.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@2724.4]
  wire  _T_57; // @[Counter.scala 293:18:@2726.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@2734.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@2737.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@2738.4]
  wire  _T_75; // @[Counter.scala 322:102:@2742.4]
  wire  _T_77; // @[Counter.scala 322:130:@2743.4]
  FF bases_0 ( // @[Counter.scala 261:53:@2677.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@2693.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@2696.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@2721.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2722.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2723.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@2724.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh780); // @[Counter.scala 293:18:@2726.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@2734.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@2737.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@2738.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 322:102:@2742.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh780); // @[Counter.scala 322:130:@2743.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@2741.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@2745.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@2747.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh780); // @[Counter.scala 340:25:@2750.4]
  assign bases_0_clock = clock; // @[:@2678.4]
  assign bases_0_reset = reset; // @[:@2679.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@2740.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@2719.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@2720.4]
  assign SRFF_clock = clock; // @[:@2694.4]
  assign SRFF_reset = reset; // @[:@2695.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@2698.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@2700.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@2701.4]
endmodule
module SingleCounter_2( // @[:@2790.2]
  input         clock, // @[:@2791.4]
  input         reset, // @[:@2792.4]
  input         io_setup_saturate, // @[:@2793.4]
  input         io_input_reset, // @[:@2793.4]
  input         io_input_enable, // @[:@2793.4]
  output [12:0] io_output_count_0, // @[:@2793.4]
  output        io_output_oobs_0, // @[:@2793.4]
  output        io_output_done // @[:@2793.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@2806.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@2806.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@2806.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@2822.4]
  wire  _T_36; // @[Counter.scala 264:45:@2825.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@2850.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@2851.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@2852.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@2853.4]
  wire  _T_57; // @[Counter.scala 293:18:@2855.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@2863.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@2865.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@2866.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@2867.4]
  wire  _T_75; // @[Counter.scala 322:102:@2871.4]
  wire  _T_77; // @[Counter.scala 322:130:@2872.4]
  FF bases_0 ( // @[Counter.scala 261:53:@2806.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@2822.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@2825.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@2850.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2851.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2852.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@2853.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh400); // @[Counter.scala 293:18:@2855.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@2863.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 299:85:@2865.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@2866.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@2867.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 322:102:@2871.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh400); // @[Counter.scala 322:130:@2872.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@2870.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@2874.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@2876.4]
  assign bases_0_clock = clock; // @[:@2807.4]
  assign bases_0_reset = reset; // @[:@2808.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@2869.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@2848.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@2849.4]
  assign SRFF_clock = clock; // @[:@2823.4]
  assign SRFF_reset = reset; // @[:@2824.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@2827.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@2829.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@2830.4]
endmodule
module x213_ctrchain( // @[:@2881.2]
  input         clock, // @[:@2882.4]
  input         reset, // @[:@2883.4]
  input         io_input_reset, // @[:@2884.4]
  input         io_input_enable, // @[:@2884.4]
  output [31:0] io_output_counts_1, // @[:@2884.4]
  output [31:0] io_output_counts_0, // @[:@2884.4]
  output        io_output_oobs_0, // @[:@2884.4]
  output        io_output_oobs_1, // @[:@2884.4]
  output        io_output_done // @[:@2884.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@2886.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@2889.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@2889.4]
  wire  isDone; // @[Counter.scala 541:51:@2906.4]
  reg  wasDone; // @[Counter.scala 542:24:@2907.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@2915.4]
  wire  _T_66; // @[Counter.scala 546:80:@2916.4]
  reg  doneLatch; // @[Counter.scala 550:26:@2921.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@2922.4]
  wire  _T_74; // @[Counter.scala 551:19:@2923.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@2886.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@2889.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@2906.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@2915.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@2916.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@2922.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@2923.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@2928.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@2925.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@2927.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@2930.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@2918.4]
  assign ctrs_0_clock = clock; // @[:@2887.4]
  assign ctrs_0_reset = reset; // @[:@2888.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@2895.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@2902.4]
  assign ctrs_1_clock = clock; // @[:@2890.4]
  assign ctrs_1_reset = reset; // @[:@2891.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@2905.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@2899.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@2900.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2970.2]
  input   clock, // @[:@2971.4]
  input   reset, // @[:@2972.4]
  input   io_flow, // @[:@2973.4]
  input   io_in, // @[:@2973.4]
  output  io_out // @[:@2973.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(62)) sr ( // @[RetimeShiftRegister.scala 15:20:@2975.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2988.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2987.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2986.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2985.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2984.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2982.4]
endmodule
module RetimeWrapper_16( // @[:@3098.2]
  input   clock, // @[:@3099.4]
  input   reset, // @[:@3100.4]
  input   io_flow, // @[:@3101.4]
  input   io_in, // @[:@3101.4]
  output  io_out // @[:@3101.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(61)) sr ( // @[RetimeShiftRegister.scala 15:20:@3103.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3116.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3115.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3114.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3113.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3112.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3110.4]
endmodule
module x325_inr_Foreach_SAMPLER_BOX_sm( // @[:@3118.2]
  input   clock, // @[:@3119.4]
  input   reset, // @[:@3120.4]
  input   io_enable, // @[:@3121.4]
  output  io_done, // @[:@3121.4]
  output  io_doneLatch, // @[:@3121.4]
  input   io_ctrDone, // @[:@3121.4]
  output  io_datapathEn, // @[:@3121.4]
  output  io_ctrInc, // @[:@3121.4]
  output  io_ctrRst, // @[:@3121.4]
  input   io_parentAck, // @[:@3121.4]
  input   io_backpressure, // @[:@3121.4]
  input   io_break // @[:@3121.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3123.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3123.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3126.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3126.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3218.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3131.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3132.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3133.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3134.4]
  wire  _T_100; // @[package.scala 100:49:@3151.4]
  reg  _T_103; // @[package.scala 48:56:@3152.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3165.4 package.scala 96:25:@3166.4]
  wire  _T_110; // @[package.scala 100:49:@3167.4]
  reg  _T_113; // @[package.scala 48:56:@3168.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3170.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3175.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3176.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3179.4]
  wire  _T_124; // @[package.scala 96:25:@3187.4 package.scala 96:25:@3188.4]
  wire  _T_126; // @[package.scala 100:49:@3189.4]
  reg  _T_129; // @[package.scala 48:56:@3190.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3212.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3214.4]
  reg  _T_153; // @[package.scala 48:56:@3215.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3223.4 package.scala 96:25:@3224.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3225.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3226.4]
  SRFF active ( // @[Controllers.scala 261:22:@3123.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3126.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3160.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3182.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3194.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3202.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3218.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3131.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3132.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3133.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3134.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3151.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3165.4 package.scala 96:25:@3166.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3167.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3170.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3175.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3176.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3179.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3187.4 package.scala 96:25:@3188.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3189.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3214.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3223.4 package.scala 96:25:@3224.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3225.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3226.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3193.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3228.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3178.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3181.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3173.4]
  assign active_clock = clock; // @[:@3124.4]
  assign active_reset = reset; // @[:@3125.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3136.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3140.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3141.4]
  assign done_clock = clock; // @[:@3127.4]
  assign done_reset = reset; // @[:@3128.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3156.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3149.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3150.4]
  assign RetimeWrapper_clock = clock; // @[:@3161.4]
  assign RetimeWrapper_reset = reset; // @[:@3162.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3164.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3163.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3183.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3184.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3186.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3185.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3195.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3196.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3198.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3197.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3203.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3204.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3206.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3205.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3219.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3220.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3222.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3221.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3335.2]
  input  [31:0] io_a, // @[:@3338.4]
  output [31:0] io_b // @[:@3338.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3351.4]
endmodule
module _( // @[:@3353.2]
  input  [31:0] io_b, // @[:@3356.4]
  output [31:0] io_result // @[:@3356.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3361.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3361.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3361.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3374.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3369.4]
endmodule
module SRAM( // @[:@3433.2]
  input        clock, // @[:@3434.4]
  input  [8:0] io_raddr, // @[:@3436.4]
  input        io_wen, // @[:@3436.4]
  input  [8:0] io_waddr, // @[:@3436.4]
  input  [7:0] io_wdata, // @[:@3436.4]
  output [7:0] io_rdata, // @[:@3436.4]
  input        io_backpressure // @[:@3436.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 143:23:@3438.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 143:23:@3438.4]
  wire [8:0] SRAMVerilogSim_waddr; // @[SRAM.scala 143:23:@3438.4]
  wire [8:0] SRAMVerilogSim_raddr; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 143:23:@3438.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(342), .AWIDTH(9)) SRAMVerilogSim ( // @[SRAM.scala 143:23:@3438.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 153:16:@3458.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 148:20:@3452.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 149:27:@3453.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 146:18:@3450.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 151:22:@3455.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 150:22:@3454.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 147:20:@3451.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 145:20:@3449.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 144:18:@3448.4]
endmodule
module RetimeWrapper_20( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_flow, // @[:@3475.4]
  input  [8:0] io_in, // @[:@3475.4]
  output [8:0] io_out // @[:@3475.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3477.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3490.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3489.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@3488.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3487.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3486.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3484.4]
endmodule
module Mem1D_4( // @[:@3492.2]
  input        clock, // @[:@3493.4]
  input        reset, // @[:@3494.4]
  input  [8:0] io_r_ofs_0, // @[:@3495.4]
  input        io_r_backpressure, // @[:@3495.4]
  input  [8:0] io_w_ofs_0, // @[:@3495.4]
  input  [7:0] io_w_data_0, // @[:@3495.4]
  input        io_w_en_0, // @[:@3495.4]
  output [7:0] io_output // @[:@3495.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_wdata; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3502.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3502.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3502.4]
  wire  wInBound; // @[MemPrimitives.scala 554:32:@3497.4]
  SRAM SRAM ( // @[MemPrimitives.scala 567:21:@3499.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_20 RetimeWrapper ( // @[package.scala 93:22:@3502.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h156; // @[MemPrimitives.scala 554:32:@3497.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 574:17:@3515.4]
  assign SRAM_clock = clock; // @[:@3500.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 568:37:@3509.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 571:22:@3512.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 570:22:@3510.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 572:22:@3513.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 573:30:@3514.4]
  assign RetimeWrapper_clock = clock; // @[:@3503.4]
  assign RetimeWrapper_reset = reset; // @[:@3504.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3506.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3505.4]
endmodule
module StickySelects( // @[:@4617.2]
  input   clock, // @[:@4618.4]
  input   reset, // @[:@4619.4]
  input   io_ins_0, // @[:@4620.4]
  input   io_ins_1, // @[:@4620.4]
  input   io_ins_2, // @[:@4620.4]
  input   io_ins_3, // @[:@4620.4]
  input   io_ins_4, // @[:@4620.4]
  input   io_ins_5, // @[:@4620.4]
  input   io_ins_6, // @[:@4620.4]
  input   io_ins_7, // @[:@4620.4]
  input   io_ins_8, // @[:@4620.4]
  output  io_outs_0, // @[:@4620.4]
  output  io_outs_1, // @[:@4620.4]
  output  io_outs_2, // @[:@4620.4]
  output  io_outs_3, // @[:@4620.4]
  output  io_outs_4, // @[:@4620.4]
  output  io_outs_5, // @[:@4620.4]
  output  io_outs_6, // @[:@4620.4]
  output  io_outs_7, // @[:@4620.4]
  output  io_outs_8 // @[:@4620.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4622.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4623.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4624.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@4625.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@4626.4]
  wire  _T_24; // @[StickySelects.scala 22:54:@4627.4]
  wire  _T_25; // @[StickySelects.scala 22:54:@4628.4]
  wire  _T_26; // @[StickySelects.scala 22:54:@4629.4]
  wire  _T_28; // @[StickySelects.scala 24:52:@4630.4]
  wire  _T_29; // @[StickySelects.scala 24:21:@4631.4]
  reg  _T_32; // @[StickySelects.scala 21:22:@4633.4]
  reg [31:0] _RAND_1;
  wire  _T_33; // @[StickySelects.scala 22:54:@4634.4]
  wire  _T_34; // @[StickySelects.scala 22:54:@4635.4]
  wire  _T_35; // @[StickySelects.scala 22:54:@4636.4]
  wire  _T_36; // @[StickySelects.scala 22:54:@4637.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@4638.4]
  wire  _T_38; // @[StickySelects.scala 22:54:@4639.4]
  wire  _T_39; // @[StickySelects.scala 22:54:@4640.4]
  wire  _T_41; // @[StickySelects.scala 24:52:@4641.4]
  wire  _T_42; // @[StickySelects.scala 24:21:@4642.4]
  reg  _T_45; // @[StickySelects.scala 21:22:@4644.4]
  reg [31:0] _RAND_2;
  wire  _T_46; // @[StickySelects.scala 22:54:@4645.4]
  wire  _T_47; // @[StickySelects.scala 22:54:@4646.4]
  wire  _T_48; // @[StickySelects.scala 22:54:@4647.4]
  wire  _T_49; // @[StickySelects.scala 22:54:@4648.4]
  wire  _T_50; // @[StickySelects.scala 22:54:@4649.4]
  wire  _T_51; // @[StickySelects.scala 22:54:@4650.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@4651.4]
  wire  _T_54; // @[StickySelects.scala 24:52:@4652.4]
  wire  _T_55; // @[StickySelects.scala 24:21:@4653.4]
  reg  _T_58; // @[StickySelects.scala 21:22:@4655.4]
  reg [31:0] _RAND_3;
  wire  _T_60; // @[StickySelects.scala 22:54:@4657.4]
  wire  _T_61; // @[StickySelects.scala 22:54:@4658.4]
  wire  _T_62; // @[StickySelects.scala 22:54:@4659.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@4660.4]
  wire  _T_64; // @[StickySelects.scala 22:54:@4661.4]
  wire  _T_65; // @[StickySelects.scala 22:54:@4662.4]
  wire  _T_67; // @[StickySelects.scala 24:52:@4663.4]
  wire  _T_68; // @[StickySelects.scala 24:21:@4664.4]
  reg  _T_71; // @[StickySelects.scala 21:22:@4666.4]
  reg [31:0] _RAND_4;
  wire  _T_74; // @[StickySelects.scala 22:54:@4669.4]
  wire  _T_75; // @[StickySelects.scala 22:54:@4670.4]
  wire  _T_76; // @[StickySelects.scala 22:54:@4671.4]
  wire  _T_77; // @[StickySelects.scala 22:54:@4672.4]
  wire  _T_78; // @[StickySelects.scala 22:54:@4673.4]
  wire  _T_80; // @[StickySelects.scala 24:52:@4674.4]
  wire  _T_81; // @[StickySelects.scala 24:21:@4675.4]
  reg  _T_84; // @[StickySelects.scala 21:22:@4677.4]
  reg [31:0] _RAND_5;
  wire  _T_88; // @[StickySelects.scala 22:54:@4681.4]
  wire  _T_89; // @[StickySelects.scala 22:54:@4682.4]
  wire  _T_90; // @[StickySelects.scala 22:54:@4683.4]
  wire  _T_91; // @[StickySelects.scala 22:54:@4684.4]
  wire  _T_93; // @[StickySelects.scala 24:52:@4685.4]
  wire  _T_94; // @[StickySelects.scala 24:21:@4686.4]
  reg  _T_97; // @[StickySelects.scala 21:22:@4688.4]
  reg [31:0] _RAND_6;
  wire  _T_102; // @[StickySelects.scala 22:54:@4693.4]
  wire  _T_103; // @[StickySelects.scala 22:54:@4694.4]
  wire  _T_104; // @[StickySelects.scala 22:54:@4695.4]
  wire  _T_106; // @[StickySelects.scala 24:52:@4696.4]
  wire  _T_107; // @[StickySelects.scala 24:21:@4697.4]
  reg  _T_110; // @[StickySelects.scala 21:22:@4699.4]
  reg [31:0] _RAND_7;
  wire  _T_116; // @[StickySelects.scala 22:54:@4705.4]
  wire  _T_117; // @[StickySelects.scala 22:54:@4706.4]
  wire  _T_119; // @[StickySelects.scala 24:52:@4707.4]
  wire  _T_120; // @[StickySelects.scala 24:21:@4708.4]
  reg  _T_123; // @[StickySelects.scala 21:22:@4710.4]
  reg [31:0] _RAND_8;
  wire  _T_130; // @[StickySelects.scala 22:54:@4717.4]
  wire  _T_132; // @[StickySelects.scala 24:52:@4718.4]
  wire  _T_133; // @[StickySelects.scala 24:21:@4719.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4623.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4624.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@4625.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@4626.4]
  assign _T_24 = _T_23 | io_ins_6; // @[StickySelects.scala 22:54:@4627.4]
  assign _T_25 = _T_24 | io_ins_7; // @[StickySelects.scala 22:54:@4628.4]
  assign _T_26 = _T_25 | io_ins_8; // @[StickySelects.scala 22:54:@4629.4]
  assign _T_28 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4630.4]
  assign _T_29 = _T_26 ? 1'h0 : _T_28; // @[StickySelects.scala 24:21:@4631.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4634.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 22:54:@4635.4]
  assign _T_35 = _T_34 | io_ins_4; // @[StickySelects.scala 22:54:@4636.4]
  assign _T_36 = _T_35 | io_ins_5; // @[StickySelects.scala 22:54:@4637.4]
  assign _T_37 = _T_36 | io_ins_6; // @[StickySelects.scala 22:54:@4638.4]
  assign _T_38 = _T_37 | io_ins_7; // @[StickySelects.scala 22:54:@4639.4]
  assign _T_39 = _T_38 | io_ins_8; // @[StickySelects.scala 22:54:@4640.4]
  assign _T_41 = io_ins_1 | _T_32; // @[StickySelects.scala 24:52:@4641.4]
  assign _T_42 = _T_39 ? 1'h0 : _T_41; // @[StickySelects.scala 24:21:@4642.4]
  assign _T_46 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4645.4]
  assign _T_47 = _T_46 | io_ins_3; // @[StickySelects.scala 22:54:@4646.4]
  assign _T_48 = _T_47 | io_ins_4; // @[StickySelects.scala 22:54:@4647.4]
  assign _T_49 = _T_48 | io_ins_5; // @[StickySelects.scala 22:54:@4648.4]
  assign _T_50 = _T_49 | io_ins_6; // @[StickySelects.scala 22:54:@4649.4]
  assign _T_51 = _T_50 | io_ins_7; // @[StickySelects.scala 22:54:@4650.4]
  assign _T_52 = _T_51 | io_ins_8; // @[StickySelects.scala 22:54:@4651.4]
  assign _T_54 = io_ins_2 | _T_45; // @[StickySelects.scala 24:52:@4652.4]
  assign _T_55 = _T_52 ? 1'h0 : _T_54; // @[StickySelects.scala 24:21:@4653.4]
  assign _T_60 = _T_46 | io_ins_2; // @[StickySelects.scala 22:54:@4657.4]
  assign _T_61 = _T_60 | io_ins_4; // @[StickySelects.scala 22:54:@4658.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 22:54:@4659.4]
  assign _T_63 = _T_62 | io_ins_6; // @[StickySelects.scala 22:54:@4660.4]
  assign _T_64 = _T_63 | io_ins_7; // @[StickySelects.scala 22:54:@4661.4]
  assign _T_65 = _T_64 | io_ins_8; // @[StickySelects.scala 22:54:@4662.4]
  assign _T_67 = io_ins_3 | _T_58; // @[StickySelects.scala 24:52:@4663.4]
  assign _T_68 = _T_65 ? 1'h0 : _T_67; // @[StickySelects.scala 24:21:@4664.4]
  assign _T_74 = _T_60 | io_ins_3; // @[StickySelects.scala 22:54:@4669.4]
  assign _T_75 = _T_74 | io_ins_5; // @[StickySelects.scala 22:54:@4670.4]
  assign _T_76 = _T_75 | io_ins_6; // @[StickySelects.scala 22:54:@4671.4]
  assign _T_77 = _T_76 | io_ins_7; // @[StickySelects.scala 22:54:@4672.4]
  assign _T_78 = _T_77 | io_ins_8; // @[StickySelects.scala 22:54:@4673.4]
  assign _T_80 = io_ins_4 | _T_71; // @[StickySelects.scala 24:52:@4674.4]
  assign _T_81 = _T_78 ? 1'h0 : _T_80; // @[StickySelects.scala 24:21:@4675.4]
  assign _T_88 = _T_74 | io_ins_4; // @[StickySelects.scala 22:54:@4681.4]
  assign _T_89 = _T_88 | io_ins_6; // @[StickySelects.scala 22:54:@4682.4]
  assign _T_90 = _T_89 | io_ins_7; // @[StickySelects.scala 22:54:@4683.4]
  assign _T_91 = _T_90 | io_ins_8; // @[StickySelects.scala 22:54:@4684.4]
  assign _T_93 = io_ins_5 | _T_84; // @[StickySelects.scala 24:52:@4685.4]
  assign _T_94 = _T_91 ? 1'h0 : _T_93; // @[StickySelects.scala 24:21:@4686.4]
  assign _T_102 = _T_88 | io_ins_5; // @[StickySelects.scala 22:54:@4693.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 22:54:@4694.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 22:54:@4695.4]
  assign _T_106 = io_ins_6 | _T_97; // @[StickySelects.scala 24:52:@4696.4]
  assign _T_107 = _T_104 ? 1'h0 : _T_106; // @[StickySelects.scala 24:21:@4697.4]
  assign _T_116 = _T_102 | io_ins_6; // @[StickySelects.scala 22:54:@4705.4]
  assign _T_117 = _T_116 | io_ins_8; // @[StickySelects.scala 22:54:@4706.4]
  assign _T_119 = io_ins_7 | _T_110; // @[StickySelects.scala 24:52:@4707.4]
  assign _T_120 = _T_117 ? 1'h0 : _T_119; // @[StickySelects.scala 24:21:@4708.4]
  assign _T_130 = _T_116 | io_ins_7; // @[StickySelects.scala 22:54:@4717.4]
  assign _T_132 = io_ins_8 | _T_123; // @[StickySelects.scala 24:52:@4718.4]
  assign _T_133 = _T_130 ? 1'h0 : _T_132; // @[StickySelects.scala 24:21:@4719.4]
  assign io_outs_0 = _T_26 ? 1'h0 : _T_28; // @[StickySelects.scala 28:52:@4721.4]
  assign io_outs_1 = _T_39 ? 1'h0 : _T_41; // @[StickySelects.scala 28:52:@4722.4]
  assign io_outs_2 = _T_52 ? 1'h0 : _T_54; // @[StickySelects.scala 28:52:@4723.4]
  assign io_outs_3 = _T_65 ? 1'h0 : _T_67; // @[StickySelects.scala 28:52:@4724.4]
  assign io_outs_4 = _T_78 ? 1'h0 : _T_80; // @[StickySelects.scala 28:52:@4725.4]
  assign io_outs_5 = _T_91 ? 1'h0 : _T_93; // @[StickySelects.scala 28:52:@4726.4]
  assign io_outs_6 = _T_104 ? 1'h0 : _T_106; // @[StickySelects.scala 28:52:@4727.4]
  assign io_outs_7 = _T_117 ? 1'h0 : _T_119; // @[StickySelects.scala 28:52:@4728.4]
  assign io_outs_8 = _T_130 ? 1'h0 : _T_132; // @[StickySelects.scala 28:52:@4729.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_32 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_58 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_71 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_84 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_97 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_110 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_123 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_26) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_28;
      end
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      if (_T_39) begin
        _T_32 <= 1'h0;
      end else begin
        _T_32 <= _T_41;
      end
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      if (_T_52) begin
        _T_45 <= 1'h0;
      end else begin
        _T_45 <= _T_54;
      end
    end
    if (reset) begin
      _T_58 <= 1'h0;
    end else begin
      if (_T_65) begin
        _T_58 <= 1'h0;
      end else begin
        _T_58 <= _T_67;
      end
    end
    if (reset) begin
      _T_71 <= 1'h0;
    end else begin
      if (_T_78) begin
        _T_71 <= 1'h0;
      end else begin
        _T_71 <= _T_80;
      end
    end
    if (reset) begin
      _T_84 <= 1'h0;
    end else begin
      if (_T_91) begin
        _T_84 <= 1'h0;
      end else begin
        _T_84 <= _T_93;
      end
    end
    if (reset) begin
      _T_97 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_97 <= 1'h0;
      end else begin
        _T_97 <= _T_106;
      end
    end
    if (reset) begin
      _T_110 <= 1'h0;
    end else begin
      if (_T_117) begin
        _T_110 <= 1'h0;
      end else begin
        _T_110 <= _T_119;
      end
    end
    if (reset) begin
      _T_123 <= 1'h0;
    end else begin
      if (_T_130) begin
        _T_123 <= 1'h0;
      end else begin
        _T_123 <= _T_132;
      end
    end
  end
endmodule
module RetimeWrapper_32( // @[:@5997.2]
  input   clock, // @[:@5998.4]
  input   reset, // @[:@5999.4]
  input   io_flow, // @[:@6000.4]
  input   io_in, // @[:@6000.4]
  output  io_out // @[:@6000.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6002.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6002.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6002.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6002.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6002.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6002.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@6002.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6015.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6014.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6013.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6012.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6011.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6009.4]
endmodule
module x218_lb_0( // @[:@9441.2]
  input        clock, // @[:@9442.4]
  input        reset, // @[:@9443.4]
  input  [1:0] io_rPort_8_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_8_ofs_0, // @[:@9444.4]
  input        io_rPort_8_en_0, // @[:@9444.4]
  input        io_rPort_8_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_8_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_7_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_7_ofs_0, // @[:@9444.4]
  input        io_rPort_7_en_0, // @[:@9444.4]
  input        io_rPort_7_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_7_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_6_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_6_ofs_0, // @[:@9444.4]
  input        io_rPort_6_en_0, // @[:@9444.4]
  input        io_rPort_6_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_6_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_5_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_5_ofs_0, // @[:@9444.4]
  input        io_rPort_5_en_0, // @[:@9444.4]
  input        io_rPort_5_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_5_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_4_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_4_ofs_0, // @[:@9444.4]
  input        io_rPort_4_en_0, // @[:@9444.4]
  input        io_rPort_4_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_4_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_3_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_3_ofs_0, // @[:@9444.4]
  input        io_rPort_3_en_0, // @[:@9444.4]
  input        io_rPort_3_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_3_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_2_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_2_ofs_0, // @[:@9444.4]
  input        io_rPort_2_en_0, // @[:@9444.4]
  input        io_rPort_2_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_2_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_1_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_1_ofs_0, // @[:@9444.4]
  input        io_rPort_1_en_0, // @[:@9444.4]
  input        io_rPort_1_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_1_output_0, // @[:@9444.4]
  input  [1:0] io_rPort_0_banks_1, // @[:@9444.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@9444.4]
  input  [8:0] io_rPort_0_ofs_0, // @[:@9444.4]
  input        io_rPort_0_en_0, // @[:@9444.4]
  input        io_rPort_0_backpressure, // @[:@9444.4]
  output [7:0] io_rPort_0_output_0, // @[:@9444.4]
  input  [1:0] io_wPort_0_banks_1, // @[:@9444.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@9444.4]
  input  [8:0] io_wPort_0_ofs_0, // @[:@9444.4]
  input  [7:0] io_wPort_0_data_0, // @[:@9444.4]
  input        io_wPort_0_en_0 // @[:@9444.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@9509.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@9509.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9509.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9509.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9509.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@9509.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@9509.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@9509.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@9525.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@9525.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9525.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9525.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9525.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@9525.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@9525.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@9525.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@9541.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@9541.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9541.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9541.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9541.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@9541.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@9541.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@9541.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@9557.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@9557.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9557.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9557.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9557.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@9557.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@9557.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@9557.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@9573.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@9573.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9573.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9573.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9573.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@9573.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@9573.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@9573.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@9589.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@9589.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9589.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9589.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9589.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@9589.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@9589.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@9589.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@9605.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@9605.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9605.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9605.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9605.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@9605.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@9605.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@9605.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@9621.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@9621.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9621.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9621.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9621.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@9621.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@9621.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@9621.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@9637.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@9637.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9637.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9637.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9637.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@9637.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@9637.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@9637.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@9653.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@9653.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9653.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9653.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9653.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@9653.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@9653.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@9653.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@9669.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@9669.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9669.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9669.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9669.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@9669.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@9669.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@9669.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@9685.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@9685.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9685.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9685.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9685.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@9685.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@9685.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@9685.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 121:29:@9881.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 121:29:@9970.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 121:29:@10059.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 121:29:@10148.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 121:29:@10237.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 121:29:@10326.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 121:29:@10415.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 121:29:@10504.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 121:29:@10593.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 121:29:@10682.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 121:29:@10771.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 121:29:@10860.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10950.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10950.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10950.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10950.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10950.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10958.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10958.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10958.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10958.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10958.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10966.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10966.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10966.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10966.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10966.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10974.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10974.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10974.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10974.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10974.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10982.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10982.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10982.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10982.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10982.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10990.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10990.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10990.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10990.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10990.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10998.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10998.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10998.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10998.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10998.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@11006.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@11006.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@11006.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@11006.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@11006.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@11014.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@11014.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@11014.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@11014.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@11014.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@11022.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@11022.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@11022.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@11022.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@11022.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@11030.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@11030.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@11030.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@11030.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@11030.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@11038.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@11038.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@11038.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@11038.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@11038.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@11094.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@11094.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@11094.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@11094.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@11094.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@11102.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@11102.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@11102.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@11102.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@11102.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@11110.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@11110.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@11110.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@11110.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@11110.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@11118.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@11118.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@11118.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@11118.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@11118.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@11126.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@11126.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@11126.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@11126.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@11126.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@11134.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@11134.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@11134.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@11134.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@11134.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@11142.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@11142.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@11142.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@11142.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@11142.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@11150.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@11150.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@11150.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@11150.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@11150.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@11158.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@11158.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@11158.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@11158.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@11158.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@11166.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@11166.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@11166.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@11166.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@11166.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@11174.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@11174.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@11174.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@11174.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@11174.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@11182.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@11182.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@11182.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@11182.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@11182.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@11246.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@11246.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@11246.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@11246.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@11246.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@11254.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@11254.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@11254.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@11254.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@11254.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@11262.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@11262.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@11262.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@11262.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@11262.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@11270.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@11270.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@11270.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@11270.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@11270.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@11278.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@11278.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@11278.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@11278.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@11278.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@11286.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@11286.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@11286.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@11286.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@11286.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@11294.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@11294.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@11294.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@11294.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@11294.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@11302.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@11302.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@11302.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@11302.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@11302.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@11310.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@11310.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@11310.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@11310.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@11310.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@11318.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@11318.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@11318.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@11318.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@11318.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@11326.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@11326.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@11326.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@11326.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@11326.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@11382.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@11382.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@11382.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@11382.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@11382.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@11390.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@11390.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@11390.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@11390.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@11390.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@11398.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@11398.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@11398.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@11398.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@11398.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@11406.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@11406.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@11406.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@11406.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@11406.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@11414.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@11414.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@11414.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@11414.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@11414.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@11422.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@11422.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@11422.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@11422.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@11422.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@11430.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@11430.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@11430.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@11430.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@11430.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@11438.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@11438.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@11438.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@11438.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@11438.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@11446.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@11446.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@11446.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@11446.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@11446.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@11454.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@11454.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@11454.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@11454.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@11454.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@11462.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@11462.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@11462.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@11462.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@11462.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@11470.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@11470.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@11470.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@11470.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@11470.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@11526.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@11526.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@11526.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@11526.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@11526.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@11534.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@11534.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@11534.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@11534.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@11534.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@11542.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@11542.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@11542.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@11542.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@11542.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@11550.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@11550.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@11550.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@11550.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@11550.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@11558.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@11558.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@11558.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@11558.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@11558.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@11566.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@11566.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@11566.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@11566.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@11566.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@11574.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@11574.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@11574.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@11574.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@11574.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@11582.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@11582.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@11582.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@11582.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@11582.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@11590.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@11590.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@11590.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@11590.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@11590.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@11598.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@11598.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@11598.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@11598.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@11598.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@11606.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@11606.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@11606.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@11606.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@11606.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@11614.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@11614.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@11614.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@11614.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@11614.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@11670.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@11670.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@11670.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@11670.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@11670.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@11678.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@11678.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@11678.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@11678.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@11678.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@11686.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@11686.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@11686.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@11686.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@11686.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@11694.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@11694.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@11694.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@11694.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@11694.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@11702.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@11702.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@11702.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@11702.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@11702.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@11710.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@11710.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@11710.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@11710.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@11710.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@11718.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@11718.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@11718.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@11718.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@11718.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@11726.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@11726.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@11726.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@11726.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@11726.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@11734.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@11734.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@11734.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@11734.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@11734.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@11742.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@11742.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@11742.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@11742.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@11742.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@11750.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@11750.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@11750.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@11750.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@11750.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@11758.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@11758.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@11758.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@11758.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@11758.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@11814.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@11814.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@11814.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@11814.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@11814.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@11822.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@11822.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@11822.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@11822.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@11822.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@11830.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@11830.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@11830.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@11830.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@11830.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@11838.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@11838.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@11838.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@11838.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@11838.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@11846.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@11846.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@11846.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@11846.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@11846.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@11854.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@11854.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@11854.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@11854.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@11854.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@11862.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@11862.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@11862.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@11862.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@11862.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@11870.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@11870.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@11870.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@11870.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@11870.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@11878.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@11878.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@11878.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@11878.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@11878.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@11886.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@11886.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@11886.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@11886.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@11886.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@11894.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@11894.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@11894.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@11894.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@11894.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@11902.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@11902.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@11902.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@11902.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@11902.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@11958.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@11958.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@11958.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@11958.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@11958.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@11966.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@11966.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@11966.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@11966.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@11966.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@11974.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@11974.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@11974.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@11974.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@11974.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@11982.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@11982.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@11982.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@11982.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@11982.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@11990.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@11990.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@11990.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@11990.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@11990.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@11998.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@11998.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@11998.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@11998.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@11998.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@12006.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@12006.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@12006.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@12006.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@12006.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@12014.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@12014.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@12014.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@12014.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@12014.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@12022.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@12022.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@12022.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@12022.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@12022.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@12030.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@12030.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@12030.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@12030.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@12030.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@12038.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@12038.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@12038.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@12038.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@12038.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@12046.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@12046.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@12046.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@12046.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@12046.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@12118.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@12118.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@12118.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@12118.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@12118.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@12126.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@12126.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@12126.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@12126.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@12126.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@12134.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@12134.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@12134.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@12134.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@12134.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@12142.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@12142.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@12142.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@12142.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@12142.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@12150.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@12150.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@12150.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@12150.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@12150.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@12158.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@12158.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@12158.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@12158.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@12158.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@12166.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@12166.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@12166.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@12166.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@12166.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@12174.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@12174.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@12174.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@12174.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@12174.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@12182.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@12182.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@12182.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@12182.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@12182.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@12190.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@12190.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@12190.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@12190.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@12190.4]
  wire  _T_316; // @[MemPrimitives.scala 82:210:@9701.4]
  wire  _T_318; // @[MemPrimitives.scala 82:210:@9702.4]
  wire  _T_319; // @[MemPrimitives.scala 82:228:@9703.4]
  wire  _T_320; // @[MemPrimitives.scala 83:102:@9704.4]
  wire [17:0] _T_322; // @[Cat.scala 30:58:@9706.4]
  wire  _T_329; // @[MemPrimitives.scala 82:210:@9714.4]
  wire  _T_330; // @[MemPrimitives.scala 82:228:@9715.4]
  wire  _T_331; // @[MemPrimitives.scala 83:102:@9716.4]
  wire [17:0] _T_333; // @[Cat.scala 30:58:@9718.4]
  wire  _T_340; // @[MemPrimitives.scala 82:210:@9726.4]
  wire  _T_341; // @[MemPrimitives.scala 82:228:@9727.4]
  wire  _T_342; // @[MemPrimitives.scala 83:102:@9728.4]
  wire [17:0] _T_344; // @[Cat.scala 30:58:@9730.4]
  wire  _T_349; // @[MemPrimitives.scala 82:210:@9737.4]
  wire  _T_352; // @[MemPrimitives.scala 82:228:@9739.4]
  wire  _T_353; // @[MemPrimitives.scala 83:102:@9740.4]
  wire [17:0] _T_355; // @[Cat.scala 30:58:@9742.4]
  wire  _T_363; // @[MemPrimitives.scala 82:228:@9751.4]
  wire  _T_364; // @[MemPrimitives.scala 83:102:@9752.4]
  wire [17:0] _T_366; // @[Cat.scala 30:58:@9754.4]
  wire  _T_374; // @[MemPrimitives.scala 82:228:@9763.4]
  wire  _T_375; // @[MemPrimitives.scala 83:102:@9764.4]
  wire [17:0] _T_377; // @[Cat.scala 30:58:@9766.4]
  wire  _T_382; // @[MemPrimitives.scala 82:210:@9773.4]
  wire  _T_385; // @[MemPrimitives.scala 82:228:@9775.4]
  wire  _T_386; // @[MemPrimitives.scala 83:102:@9776.4]
  wire [17:0] _T_388; // @[Cat.scala 30:58:@9778.4]
  wire  _T_396; // @[MemPrimitives.scala 82:228:@9787.4]
  wire  _T_397; // @[MemPrimitives.scala 83:102:@9788.4]
  wire [17:0] _T_399; // @[Cat.scala 30:58:@9790.4]
  wire  _T_407; // @[MemPrimitives.scala 82:228:@9799.4]
  wire  _T_408; // @[MemPrimitives.scala 83:102:@9800.4]
  wire [17:0] _T_410; // @[Cat.scala 30:58:@9802.4]
  wire  _T_415; // @[MemPrimitives.scala 82:210:@9809.4]
  wire  _T_418; // @[MemPrimitives.scala 82:228:@9811.4]
  wire  _T_419; // @[MemPrimitives.scala 83:102:@9812.4]
  wire [17:0] _T_421; // @[Cat.scala 30:58:@9814.4]
  wire  _T_429; // @[MemPrimitives.scala 82:228:@9823.4]
  wire  _T_430; // @[MemPrimitives.scala 83:102:@9824.4]
  wire [17:0] _T_432; // @[Cat.scala 30:58:@9826.4]
  wire  _T_440; // @[MemPrimitives.scala 82:228:@9835.4]
  wire  _T_441; // @[MemPrimitives.scala 83:102:@9836.4]
  wire [17:0] _T_443; // @[Cat.scala 30:58:@9838.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@9845.4]
  wire  _T_450; // @[MemPrimitives.scala 110:210:@9846.4]
  wire  _T_451; // @[MemPrimitives.scala 110:228:@9847.4]
  wire  _T_454; // @[MemPrimitives.scala 110:210:@9849.4]
  wire  _T_456; // @[MemPrimitives.scala 110:210:@9850.4]
  wire  _T_457; // @[MemPrimitives.scala 110:228:@9851.4]
  wire  _T_460; // @[MemPrimitives.scala 110:210:@9853.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@9854.4]
  wire  _T_463; // @[MemPrimitives.scala 110:228:@9855.4]
  wire  _T_466; // @[MemPrimitives.scala 110:210:@9857.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@9858.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@9859.4]
  wire  _T_472; // @[MemPrimitives.scala 110:210:@9861.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@9862.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@9863.4]
  wire  _T_478; // @[MemPrimitives.scala 110:210:@9865.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@9866.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@9867.4]
  wire  _T_484; // @[MemPrimitives.scala 110:210:@9869.4]
  wire  _T_486; // @[MemPrimitives.scala 110:210:@9870.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@9871.4]
  wire  _T_490; // @[MemPrimitives.scala 110:210:@9873.4]
  wire  _T_492; // @[MemPrimitives.scala 110:210:@9874.4]
  wire  _T_493; // @[MemPrimitives.scala 110:228:@9875.4]
  wire  _T_496; // @[MemPrimitives.scala 110:210:@9877.4]
  wire  _T_498; // @[MemPrimitives.scala 110:210:@9878.4]
  wire  _T_499; // @[MemPrimitives.scala 110:228:@9879.4]
  wire  _T_501; // @[MemPrimitives.scala 123:41:@9893.4]
  wire  _T_502; // @[MemPrimitives.scala 123:41:@9894.4]
  wire  _T_503; // @[MemPrimitives.scala 123:41:@9895.4]
  wire  _T_504; // @[MemPrimitives.scala 123:41:@9896.4]
  wire  _T_505; // @[MemPrimitives.scala 123:41:@9897.4]
  wire  _T_506; // @[MemPrimitives.scala 123:41:@9898.4]
  wire  _T_507; // @[MemPrimitives.scala 123:41:@9899.4]
  wire  _T_508; // @[MemPrimitives.scala 123:41:@9900.4]
  wire  _T_509; // @[MemPrimitives.scala 123:41:@9901.4]
  wire [10:0] _T_511; // @[Cat.scala 30:58:@9903.4]
  wire [10:0] _T_513; // @[Cat.scala 30:58:@9905.4]
  wire [10:0] _T_515; // @[Cat.scala 30:58:@9907.4]
  wire [10:0] _T_517; // @[Cat.scala 30:58:@9909.4]
  wire [10:0] _T_519; // @[Cat.scala 30:58:@9911.4]
  wire [10:0] _T_521; // @[Cat.scala 30:58:@9913.4]
  wire [10:0] _T_523; // @[Cat.scala 30:58:@9915.4]
  wire [10:0] _T_525; // @[Cat.scala 30:58:@9917.4]
  wire [10:0] _T_527; // @[Cat.scala 30:58:@9919.4]
  wire [10:0] _T_528; // @[Mux.scala 31:69:@9920.4]
  wire [10:0] _T_529; // @[Mux.scala 31:69:@9921.4]
  wire [10:0] _T_530; // @[Mux.scala 31:69:@9922.4]
  wire [10:0] _T_531; // @[Mux.scala 31:69:@9923.4]
  wire [10:0] _T_532; // @[Mux.scala 31:69:@9924.4]
  wire [10:0] _T_533; // @[Mux.scala 31:69:@9925.4]
  wire [10:0] _T_534; // @[Mux.scala 31:69:@9926.4]
  wire [10:0] _T_535; // @[Mux.scala 31:69:@9927.4]
  wire  _T_542; // @[MemPrimitives.scala 110:210:@9935.4]
  wire  _T_543; // @[MemPrimitives.scala 110:228:@9936.4]
  wire  _T_548; // @[MemPrimitives.scala 110:210:@9939.4]
  wire  _T_549; // @[MemPrimitives.scala 110:228:@9940.4]
  wire  _T_554; // @[MemPrimitives.scala 110:210:@9943.4]
  wire  _T_555; // @[MemPrimitives.scala 110:228:@9944.4]
  wire  _T_560; // @[MemPrimitives.scala 110:210:@9947.4]
  wire  _T_561; // @[MemPrimitives.scala 110:228:@9948.4]
  wire  _T_566; // @[MemPrimitives.scala 110:210:@9951.4]
  wire  _T_567; // @[MemPrimitives.scala 110:228:@9952.4]
  wire  _T_572; // @[MemPrimitives.scala 110:210:@9955.4]
  wire  _T_573; // @[MemPrimitives.scala 110:228:@9956.4]
  wire  _T_578; // @[MemPrimitives.scala 110:210:@9959.4]
  wire  _T_579; // @[MemPrimitives.scala 110:228:@9960.4]
  wire  _T_584; // @[MemPrimitives.scala 110:210:@9963.4]
  wire  _T_585; // @[MemPrimitives.scala 110:228:@9964.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@9967.4]
  wire  _T_591; // @[MemPrimitives.scala 110:228:@9968.4]
  wire  _T_593; // @[MemPrimitives.scala 123:41:@9982.4]
  wire  _T_594; // @[MemPrimitives.scala 123:41:@9983.4]
  wire  _T_595; // @[MemPrimitives.scala 123:41:@9984.4]
  wire  _T_596; // @[MemPrimitives.scala 123:41:@9985.4]
  wire  _T_597; // @[MemPrimitives.scala 123:41:@9986.4]
  wire  _T_598; // @[MemPrimitives.scala 123:41:@9987.4]
  wire  _T_599; // @[MemPrimitives.scala 123:41:@9988.4]
  wire  _T_600; // @[MemPrimitives.scala 123:41:@9989.4]
  wire  _T_601; // @[MemPrimitives.scala 123:41:@9990.4]
  wire [10:0] _T_603; // @[Cat.scala 30:58:@9992.4]
  wire [10:0] _T_605; // @[Cat.scala 30:58:@9994.4]
  wire [10:0] _T_607; // @[Cat.scala 30:58:@9996.4]
  wire [10:0] _T_609; // @[Cat.scala 30:58:@9998.4]
  wire [10:0] _T_611; // @[Cat.scala 30:58:@10000.4]
  wire [10:0] _T_613; // @[Cat.scala 30:58:@10002.4]
  wire [10:0] _T_615; // @[Cat.scala 30:58:@10004.4]
  wire [10:0] _T_617; // @[Cat.scala 30:58:@10006.4]
  wire [10:0] _T_619; // @[Cat.scala 30:58:@10008.4]
  wire [10:0] _T_620; // @[Mux.scala 31:69:@10009.4]
  wire [10:0] _T_621; // @[Mux.scala 31:69:@10010.4]
  wire [10:0] _T_622; // @[Mux.scala 31:69:@10011.4]
  wire [10:0] _T_623; // @[Mux.scala 31:69:@10012.4]
  wire [10:0] _T_624; // @[Mux.scala 31:69:@10013.4]
  wire [10:0] _T_625; // @[Mux.scala 31:69:@10014.4]
  wire [10:0] _T_626; // @[Mux.scala 31:69:@10015.4]
  wire [10:0] _T_627; // @[Mux.scala 31:69:@10016.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@10024.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@10025.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@10028.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@10029.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@10032.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@10033.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@10036.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@10037.4]
  wire  _T_658; // @[MemPrimitives.scala 110:210:@10040.4]
  wire  _T_659; // @[MemPrimitives.scala 110:228:@10041.4]
  wire  _T_664; // @[MemPrimitives.scala 110:210:@10044.4]
  wire  _T_665; // @[MemPrimitives.scala 110:228:@10045.4]
  wire  _T_670; // @[MemPrimitives.scala 110:210:@10048.4]
  wire  _T_671; // @[MemPrimitives.scala 110:228:@10049.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@10052.4]
  wire  _T_677; // @[MemPrimitives.scala 110:228:@10053.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@10056.4]
  wire  _T_683; // @[MemPrimitives.scala 110:228:@10057.4]
  wire  _T_685; // @[MemPrimitives.scala 123:41:@10071.4]
  wire  _T_686; // @[MemPrimitives.scala 123:41:@10072.4]
  wire  _T_687; // @[MemPrimitives.scala 123:41:@10073.4]
  wire  _T_688; // @[MemPrimitives.scala 123:41:@10074.4]
  wire  _T_689; // @[MemPrimitives.scala 123:41:@10075.4]
  wire  _T_690; // @[MemPrimitives.scala 123:41:@10076.4]
  wire  _T_691; // @[MemPrimitives.scala 123:41:@10077.4]
  wire  _T_692; // @[MemPrimitives.scala 123:41:@10078.4]
  wire  _T_693; // @[MemPrimitives.scala 123:41:@10079.4]
  wire [10:0] _T_695; // @[Cat.scala 30:58:@10081.4]
  wire [10:0] _T_697; // @[Cat.scala 30:58:@10083.4]
  wire [10:0] _T_699; // @[Cat.scala 30:58:@10085.4]
  wire [10:0] _T_701; // @[Cat.scala 30:58:@10087.4]
  wire [10:0] _T_703; // @[Cat.scala 30:58:@10089.4]
  wire [10:0] _T_705; // @[Cat.scala 30:58:@10091.4]
  wire [10:0] _T_707; // @[Cat.scala 30:58:@10093.4]
  wire [10:0] _T_709; // @[Cat.scala 30:58:@10095.4]
  wire [10:0] _T_711; // @[Cat.scala 30:58:@10097.4]
  wire [10:0] _T_712; // @[Mux.scala 31:69:@10098.4]
  wire [10:0] _T_713; // @[Mux.scala 31:69:@10099.4]
  wire [10:0] _T_714; // @[Mux.scala 31:69:@10100.4]
  wire [10:0] _T_715; // @[Mux.scala 31:69:@10101.4]
  wire [10:0] _T_716; // @[Mux.scala 31:69:@10102.4]
  wire [10:0] _T_717; // @[Mux.scala 31:69:@10103.4]
  wire [10:0] _T_718; // @[Mux.scala 31:69:@10104.4]
  wire [10:0] _T_719; // @[Mux.scala 31:69:@10105.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@10112.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@10114.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@10116.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@10118.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@10120.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@10122.4]
  wire  _T_742; // @[MemPrimitives.scala 110:210:@10124.4]
  wire  _T_745; // @[MemPrimitives.scala 110:228:@10126.4]
  wire  _T_748; // @[MemPrimitives.scala 110:210:@10128.4]
  wire  _T_751; // @[MemPrimitives.scala 110:228:@10130.4]
  wire  _T_754; // @[MemPrimitives.scala 110:210:@10132.4]
  wire  _T_757; // @[MemPrimitives.scala 110:228:@10134.4]
  wire  _T_760; // @[MemPrimitives.scala 110:210:@10136.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@10138.4]
  wire  _T_766; // @[MemPrimitives.scala 110:210:@10140.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@10142.4]
  wire  _T_772; // @[MemPrimitives.scala 110:210:@10144.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@10146.4]
  wire  _T_777; // @[MemPrimitives.scala 123:41:@10160.4]
  wire  _T_778; // @[MemPrimitives.scala 123:41:@10161.4]
  wire  _T_779; // @[MemPrimitives.scala 123:41:@10162.4]
  wire  _T_780; // @[MemPrimitives.scala 123:41:@10163.4]
  wire  _T_781; // @[MemPrimitives.scala 123:41:@10164.4]
  wire  _T_782; // @[MemPrimitives.scala 123:41:@10165.4]
  wire  _T_783; // @[MemPrimitives.scala 123:41:@10166.4]
  wire  _T_784; // @[MemPrimitives.scala 123:41:@10167.4]
  wire  _T_785; // @[MemPrimitives.scala 123:41:@10168.4]
  wire [10:0] _T_787; // @[Cat.scala 30:58:@10170.4]
  wire [10:0] _T_789; // @[Cat.scala 30:58:@10172.4]
  wire [10:0] _T_791; // @[Cat.scala 30:58:@10174.4]
  wire [10:0] _T_793; // @[Cat.scala 30:58:@10176.4]
  wire [10:0] _T_795; // @[Cat.scala 30:58:@10178.4]
  wire [10:0] _T_797; // @[Cat.scala 30:58:@10180.4]
  wire [10:0] _T_799; // @[Cat.scala 30:58:@10182.4]
  wire [10:0] _T_801; // @[Cat.scala 30:58:@10184.4]
  wire [10:0] _T_803; // @[Cat.scala 30:58:@10186.4]
  wire [10:0] _T_804; // @[Mux.scala 31:69:@10187.4]
  wire [10:0] _T_805; // @[Mux.scala 31:69:@10188.4]
  wire [10:0] _T_806; // @[Mux.scala 31:69:@10189.4]
  wire [10:0] _T_807; // @[Mux.scala 31:69:@10190.4]
  wire [10:0] _T_808; // @[Mux.scala 31:69:@10191.4]
  wire [10:0] _T_809; // @[Mux.scala 31:69:@10192.4]
  wire [10:0] _T_810; // @[Mux.scala 31:69:@10193.4]
  wire [10:0] _T_811; // @[Mux.scala 31:69:@10194.4]
  wire  _T_819; // @[MemPrimitives.scala 110:228:@10203.4]
  wire  _T_825; // @[MemPrimitives.scala 110:228:@10207.4]
  wire  _T_831; // @[MemPrimitives.scala 110:228:@10211.4]
  wire  _T_837; // @[MemPrimitives.scala 110:228:@10215.4]
  wire  _T_843; // @[MemPrimitives.scala 110:228:@10219.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@10223.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@10227.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@10231.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@10235.4]
  wire  _T_869; // @[MemPrimitives.scala 123:41:@10249.4]
  wire  _T_870; // @[MemPrimitives.scala 123:41:@10250.4]
  wire  _T_871; // @[MemPrimitives.scala 123:41:@10251.4]
  wire  _T_872; // @[MemPrimitives.scala 123:41:@10252.4]
  wire  _T_873; // @[MemPrimitives.scala 123:41:@10253.4]
  wire  _T_874; // @[MemPrimitives.scala 123:41:@10254.4]
  wire  _T_875; // @[MemPrimitives.scala 123:41:@10255.4]
  wire  _T_876; // @[MemPrimitives.scala 123:41:@10256.4]
  wire  _T_877; // @[MemPrimitives.scala 123:41:@10257.4]
  wire [10:0] _T_879; // @[Cat.scala 30:58:@10259.4]
  wire [10:0] _T_881; // @[Cat.scala 30:58:@10261.4]
  wire [10:0] _T_883; // @[Cat.scala 30:58:@10263.4]
  wire [10:0] _T_885; // @[Cat.scala 30:58:@10265.4]
  wire [10:0] _T_887; // @[Cat.scala 30:58:@10267.4]
  wire [10:0] _T_889; // @[Cat.scala 30:58:@10269.4]
  wire [10:0] _T_891; // @[Cat.scala 30:58:@10271.4]
  wire [10:0] _T_893; // @[Cat.scala 30:58:@10273.4]
  wire [10:0] _T_895; // @[Cat.scala 30:58:@10275.4]
  wire [10:0] _T_896; // @[Mux.scala 31:69:@10276.4]
  wire [10:0] _T_897; // @[Mux.scala 31:69:@10277.4]
  wire [10:0] _T_898; // @[Mux.scala 31:69:@10278.4]
  wire [10:0] _T_899; // @[Mux.scala 31:69:@10279.4]
  wire [10:0] _T_900; // @[Mux.scala 31:69:@10280.4]
  wire [10:0] _T_901; // @[Mux.scala 31:69:@10281.4]
  wire [10:0] _T_902; // @[Mux.scala 31:69:@10282.4]
  wire [10:0] _T_903; // @[Mux.scala 31:69:@10283.4]
  wire  _T_911; // @[MemPrimitives.scala 110:228:@10292.4]
  wire  _T_917; // @[MemPrimitives.scala 110:228:@10296.4]
  wire  _T_923; // @[MemPrimitives.scala 110:228:@10300.4]
  wire  _T_929; // @[MemPrimitives.scala 110:228:@10304.4]
  wire  _T_935; // @[MemPrimitives.scala 110:228:@10308.4]
  wire  _T_941; // @[MemPrimitives.scala 110:228:@10312.4]
  wire  _T_947; // @[MemPrimitives.scala 110:228:@10316.4]
  wire  _T_953; // @[MemPrimitives.scala 110:228:@10320.4]
  wire  _T_959; // @[MemPrimitives.scala 110:228:@10324.4]
  wire  _T_961; // @[MemPrimitives.scala 123:41:@10338.4]
  wire  _T_962; // @[MemPrimitives.scala 123:41:@10339.4]
  wire  _T_963; // @[MemPrimitives.scala 123:41:@10340.4]
  wire  _T_964; // @[MemPrimitives.scala 123:41:@10341.4]
  wire  _T_965; // @[MemPrimitives.scala 123:41:@10342.4]
  wire  _T_966; // @[MemPrimitives.scala 123:41:@10343.4]
  wire  _T_967; // @[MemPrimitives.scala 123:41:@10344.4]
  wire  _T_968; // @[MemPrimitives.scala 123:41:@10345.4]
  wire  _T_969; // @[MemPrimitives.scala 123:41:@10346.4]
  wire [10:0] _T_971; // @[Cat.scala 30:58:@10348.4]
  wire [10:0] _T_973; // @[Cat.scala 30:58:@10350.4]
  wire [10:0] _T_975; // @[Cat.scala 30:58:@10352.4]
  wire [10:0] _T_977; // @[Cat.scala 30:58:@10354.4]
  wire [10:0] _T_979; // @[Cat.scala 30:58:@10356.4]
  wire [10:0] _T_981; // @[Cat.scala 30:58:@10358.4]
  wire [10:0] _T_983; // @[Cat.scala 30:58:@10360.4]
  wire [10:0] _T_985; // @[Cat.scala 30:58:@10362.4]
  wire [10:0] _T_987; // @[Cat.scala 30:58:@10364.4]
  wire [10:0] _T_988; // @[Mux.scala 31:69:@10365.4]
  wire [10:0] _T_989; // @[Mux.scala 31:69:@10366.4]
  wire [10:0] _T_990; // @[Mux.scala 31:69:@10367.4]
  wire [10:0] _T_991; // @[Mux.scala 31:69:@10368.4]
  wire [10:0] _T_992; // @[Mux.scala 31:69:@10369.4]
  wire [10:0] _T_993; // @[Mux.scala 31:69:@10370.4]
  wire [10:0] _T_994; // @[Mux.scala 31:69:@10371.4]
  wire [10:0] _T_995; // @[Mux.scala 31:69:@10372.4]
  wire  _T_1000; // @[MemPrimitives.scala 110:210:@10379.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@10381.4]
  wire  _T_1006; // @[MemPrimitives.scala 110:210:@10383.4]
  wire  _T_1009; // @[MemPrimitives.scala 110:228:@10385.4]
  wire  _T_1012; // @[MemPrimitives.scala 110:210:@10387.4]
  wire  _T_1015; // @[MemPrimitives.scala 110:228:@10389.4]
  wire  _T_1018; // @[MemPrimitives.scala 110:210:@10391.4]
  wire  _T_1021; // @[MemPrimitives.scala 110:228:@10393.4]
  wire  _T_1024; // @[MemPrimitives.scala 110:210:@10395.4]
  wire  _T_1027; // @[MemPrimitives.scala 110:228:@10397.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@10399.4]
  wire  _T_1033; // @[MemPrimitives.scala 110:228:@10401.4]
  wire  _T_1036; // @[MemPrimitives.scala 110:210:@10403.4]
  wire  _T_1039; // @[MemPrimitives.scala 110:228:@10405.4]
  wire  _T_1042; // @[MemPrimitives.scala 110:210:@10407.4]
  wire  _T_1045; // @[MemPrimitives.scala 110:228:@10409.4]
  wire  _T_1048; // @[MemPrimitives.scala 110:210:@10411.4]
  wire  _T_1051; // @[MemPrimitives.scala 110:228:@10413.4]
  wire  _T_1053; // @[MemPrimitives.scala 123:41:@10427.4]
  wire  _T_1054; // @[MemPrimitives.scala 123:41:@10428.4]
  wire  _T_1055; // @[MemPrimitives.scala 123:41:@10429.4]
  wire  _T_1056; // @[MemPrimitives.scala 123:41:@10430.4]
  wire  _T_1057; // @[MemPrimitives.scala 123:41:@10431.4]
  wire  _T_1058; // @[MemPrimitives.scala 123:41:@10432.4]
  wire  _T_1059; // @[MemPrimitives.scala 123:41:@10433.4]
  wire  _T_1060; // @[MemPrimitives.scala 123:41:@10434.4]
  wire  _T_1061; // @[MemPrimitives.scala 123:41:@10435.4]
  wire [10:0] _T_1063; // @[Cat.scala 30:58:@10437.4]
  wire [10:0] _T_1065; // @[Cat.scala 30:58:@10439.4]
  wire [10:0] _T_1067; // @[Cat.scala 30:58:@10441.4]
  wire [10:0] _T_1069; // @[Cat.scala 30:58:@10443.4]
  wire [10:0] _T_1071; // @[Cat.scala 30:58:@10445.4]
  wire [10:0] _T_1073; // @[Cat.scala 30:58:@10447.4]
  wire [10:0] _T_1075; // @[Cat.scala 30:58:@10449.4]
  wire [10:0] _T_1077; // @[Cat.scala 30:58:@10451.4]
  wire [10:0] _T_1079; // @[Cat.scala 30:58:@10453.4]
  wire [10:0] _T_1080; // @[Mux.scala 31:69:@10454.4]
  wire [10:0] _T_1081; // @[Mux.scala 31:69:@10455.4]
  wire [10:0] _T_1082; // @[Mux.scala 31:69:@10456.4]
  wire [10:0] _T_1083; // @[Mux.scala 31:69:@10457.4]
  wire [10:0] _T_1084; // @[Mux.scala 31:69:@10458.4]
  wire [10:0] _T_1085; // @[Mux.scala 31:69:@10459.4]
  wire [10:0] _T_1086; // @[Mux.scala 31:69:@10460.4]
  wire [10:0] _T_1087; // @[Mux.scala 31:69:@10461.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@10470.4]
  wire  _T_1101; // @[MemPrimitives.scala 110:228:@10474.4]
  wire  _T_1107; // @[MemPrimitives.scala 110:228:@10478.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:228:@10482.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@10486.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@10490.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@10494.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@10498.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@10502.4]
  wire  _T_1145; // @[MemPrimitives.scala 123:41:@10516.4]
  wire  _T_1146; // @[MemPrimitives.scala 123:41:@10517.4]
  wire  _T_1147; // @[MemPrimitives.scala 123:41:@10518.4]
  wire  _T_1148; // @[MemPrimitives.scala 123:41:@10519.4]
  wire  _T_1149; // @[MemPrimitives.scala 123:41:@10520.4]
  wire  _T_1150; // @[MemPrimitives.scala 123:41:@10521.4]
  wire  _T_1151; // @[MemPrimitives.scala 123:41:@10522.4]
  wire  _T_1152; // @[MemPrimitives.scala 123:41:@10523.4]
  wire  _T_1153; // @[MemPrimitives.scala 123:41:@10524.4]
  wire [10:0] _T_1155; // @[Cat.scala 30:58:@10526.4]
  wire [10:0] _T_1157; // @[Cat.scala 30:58:@10528.4]
  wire [10:0] _T_1159; // @[Cat.scala 30:58:@10530.4]
  wire [10:0] _T_1161; // @[Cat.scala 30:58:@10532.4]
  wire [10:0] _T_1163; // @[Cat.scala 30:58:@10534.4]
  wire [10:0] _T_1165; // @[Cat.scala 30:58:@10536.4]
  wire [10:0] _T_1167; // @[Cat.scala 30:58:@10538.4]
  wire [10:0] _T_1169; // @[Cat.scala 30:58:@10540.4]
  wire [10:0] _T_1171; // @[Cat.scala 30:58:@10542.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@10543.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@10544.4]
  wire [10:0] _T_1174; // @[Mux.scala 31:69:@10545.4]
  wire [10:0] _T_1175; // @[Mux.scala 31:69:@10546.4]
  wire [10:0] _T_1176; // @[Mux.scala 31:69:@10547.4]
  wire [10:0] _T_1177; // @[Mux.scala 31:69:@10548.4]
  wire [10:0] _T_1178; // @[Mux.scala 31:69:@10549.4]
  wire [10:0] _T_1179; // @[Mux.scala 31:69:@10550.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@10559.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@10563.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@10567.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@10571.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@10575.4]
  wire  _T_1217; // @[MemPrimitives.scala 110:228:@10579.4]
  wire  _T_1223; // @[MemPrimitives.scala 110:228:@10583.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:228:@10587.4]
  wire  _T_1235; // @[MemPrimitives.scala 110:228:@10591.4]
  wire  _T_1237; // @[MemPrimitives.scala 123:41:@10605.4]
  wire  _T_1238; // @[MemPrimitives.scala 123:41:@10606.4]
  wire  _T_1239; // @[MemPrimitives.scala 123:41:@10607.4]
  wire  _T_1240; // @[MemPrimitives.scala 123:41:@10608.4]
  wire  _T_1241; // @[MemPrimitives.scala 123:41:@10609.4]
  wire  _T_1242; // @[MemPrimitives.scala 123:41:@10610.4]
  wire  _T_1243; // @[MemPrimitives.scala 123:41:@10611.4]
  wire  _T_1244; // @[MemPrimitives.scala 123:41:@10612.4]
  wire  _T_1245; // @[MemPrimitives.scala 123:41:@10613.4]
  wire [10:0] _T_1247; // @[Cat.scala 30:58:@10615.4]
  wire [10:0] _T_1249; // @[Cat.scala 30:58:@10617.4]
  wire [10:0] _T_1251; // @[Cat.scala 30:58:@10619.4]
  wire [10:0] _T_1253; // @[Cat.scala 30:58:@10621.4]
  wire [10:0] _T_1255; // @[Cat.scala 30:58:@10623.4]
  wire [10:0] _T_1257; // @[Cat.scala 30:58:@10625.4]
  wire [10:0] _T_1259; // @[Cat.scala 30:58:@10627.4]
  wire [10:0] _T_1261; // @[Cat.scala 30:58:@10629.4]
  wire [10:0] _T_1263; // @[Cat.scala 30:58:@10631.4]
  wire [10:0] _T_1264; // @[Mux.scala 31:69:@10632.4]
  wire [10:0] _T_1265; // @[Mux.scala 31:69:@10633.4]
  wire [10:0] _T_1266; // @[Mux.scala 31:69:@10634.4]
  wire [10:0] _T_1267; // @[Mux.scala 31:69:@10635.4]
  wire [10:0] _T_1268; // @[Mux.scala 31:69:@10636.4]
  wire [10:0] _T_1269; // @[Mux.scala 31:69:@10637.4]
  wire [10:0] _T_1270; // @[Mux.scala 31:69:@10638.4]
  wire [10:0] _T_1271; // @[Mux.scala 31:69:@10639.4]
  wire  _T_1276; // @[MemPrimitives.scala 110:210:@10646.4]
  wire  _T_1279; // @[MemPrimitives.scala 110:228:@10648.4]
  wire  _T_1282; // @[MemPrimitives.scala 110:210:@10650.4]
  wire  _T_1285; // @[MemPrimitives.scala 110:228:@10652.4]
  wire  _T_1288; // @[MemPrimitives.scala 110:210:@10654.4]
  wire  _T_1291; // @[MemPrimitives.scala 110:228:@10656.4]
  wire  _T_1294; // @[MemPrimitives.scala 110:210:@10658.4]
  wire  _T_1297; // @[MemPrimitives.scala 110:228:@10660.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@10662.4]
  wire  _T_1303; // @[MemPrimitives.scala 110:228:@10664.4]
  wire  _T_1306; // @[MemPrimitives.scala 110:210:@10666.4]
  wire  _T_1309; // @[MemPrimitives.scala 110:228:@10668.4]
  wire  _T_1312; // @[MemPrimitives.scala 110:210:@10670.4]
  wire  _T_1315; // @[MemPrimitives.scala 110:228:@10672.4]
  wire  _T_1318; // @[MemPrimitives.scala 110:210:@10674.4]
  wire  _T_1321; // @[MemPrimitives.scala 110:228:@10676.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@10678.4]
  wire  _T_1327; // @[MemPrimitives.scala 110:228:@10680.4]
  wire  _T_1329; // @[MemPrimitives.scala 123:41:@10694.4]
  wire  _T_1330; // @[MemPrimitives.scala 123:41:@10695.4]
  wire  _T_1331; // @[MemPrimitives.scala 123:41:@10696.4]
  wire  _T_1332; // @[MemPrimitives.scala 123:41:@10697.4]
  wire  _T_1333; // @[MemPrimitives.scala 123:41:@10698.4]
  wire  _T_1334; // @[MemPrimitives.scala 123:41:@10699.4]
  wire  _T_1335; // @[MemPrimitives.scala 123:41:@10700.4]
  wire  _T_1336; // @[MemPrimitives.scala 123:41:@10701.4]
  wire  _T_1337; // @[MemPrimitives.scala 123:41:@10702.4]
  wire [10:0] _T_1339; // @[Cat.scala 30:58:@10704.4]
  wire [10:0] _T_1341; // @[Cat.scala 30:58:@10706.4]
  wire [10:0] _T_1343; // @[Cat.scala 30:58:@10708.4]
  wire [10:0] _T_1345; // @[Cat.scala 30:58:@10710.4]
  wire [10:0] _T_1347; // @[Cat.scala 30:58:@10712.4]
  wire [10:0] _T_1349; // @[Cat.scala 30:58:@10714.4]
  wire [10:0] _T_1351; // @[Cat.scala 30:58:@10716.4]
  wire [10:0] _T_1353; // @[Cat.scala 30:58:@10718.4]
  wire [10:0] _T_1355; // @[Cat.scala 30:58:@10720.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@10721.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@10722.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@10723.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@10724.4]
  wire [10:0] _T_1360; // @[Mux.scala 31:69:@10725.4]
  wire [10:0] _T_1361; // @[Mux.scala 31:69:@10726.4]
  wire [10:0] _T_1362; // @[Mux.scala 31:69:@10727.4]
  wire [10:0] _T_1363; // @[Mux.scala 31:69:@10728.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@10737.4]
  wire  _T_1377; // @[MemPrimitives.scala 110:228:@10741.4]
  wire  _T_1383; // @[MemPrimitives.scala 110:228:@10745.4]
  wire  _T_1389; // @[MemPrimitives.scala 110:228:@10749.4]
  wire  _T_1395; // @[MemPrimitives.scala 110:228:@10753.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:228:@10757.4]
  wire  _T_1407; // @[MemPrimitives.scala 110:228:@10761.4]
  wire  _T_1413; // @[MemPrimitives.scala 110:228:@10765.4]
  wire  _T_1419; // @[MemPrimitives.scala 110:228:@10769.4]
  wire  _T_1421; // @[MemPrimitives.scala 123:41:@10783.4]
  wire  _T_1422; // @[MemPrimitives.scala 123:41:@10784.4]
  wire  _T_1423; // @[MemPrimitives.scala 123:41:@10785.4]
  wire  _T_1424; // @[MemPrimitives.scala 123:41:@10786.4]
  wire  _T_1425; // @[MemPrimitives.scala 123:41:@10787.4]
  wire  _T_1426; // @[MemPrimitives.scala 123:41:@10788.4]
  wire  _T_1427; // @[MemPrimitives.scala 123:41:@10789.4]
  wire  _T_1428; // @[MemPrimitives.scala 123:41:@10790.4]
  wire  _T_1429; // @[MemPrimitives.scala 123:41:@10791.4]
  wire [10:0] _T_1431; // @[Cat.scala 30:58:@10793.4]
  wire [10:0] _T_1433; // @[Cat.scala 30:58:@10795.4]
  wire [10:0] _T_1435; // @[Cat.scala 30:58:@10797.4]
  wire [10:0] _T_1437; // @[Cat.scala 30:58:@10799.4]
  wire [10:0] _T_1439; // @[Cat.scala 30:58:@10801.4]
  wire [10:0] _T_1441; // @[Cat.scala 30:58:@10803.4]
  wire [10:0] _T_1443; // @[Cat.scala 30:58:@10805.4]
  wire [10:0] _T_1445; // @[Cat.scala 30:58:@10807.4]
  wire [10:0] _T_1447; // @[Cat.scala 30:58:@10809.4]
  wire [10:0] _T_1448; // @[Mux.scala 31:69:@10810.4]
  wire [10:0] _T_1449; // @[Mux.scala 31:69:@10811.4]
  wire [10:0] _T_1450; // @[Mux.scala 31:69:@10812.4]
  wire [10:0] _T_1451; // @[Mux.scala 31:69:@10813.4]
  wire [10:0] _T_1452; // @[Mux.scala 31:69:@10814.4]
  wire [10:0] _T_1453; // @[Mux.scala 31:69:@10815.4]
  wire [10:0] _T_1454; // @[Mux.scala 31:69:@10816.4]
  wire [10:0] _T_1455; // @[Mux.scala 31:69:@10817.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@10826.4]
  wire  _T_1469; // @[MemPrimitives.scala 110:228:@10830.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:228:@10834.4]
  wire  _T_1481; // @[MemPrimitives.scala 110:228:@10838.4]
  wire  _T_1487; // @[MemPrimitives.scala 110:228:@10842.4]
  wire  _T_1493; // @[MemPrimitives.scala 110:228:@10846.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:228:@10850.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:228:@10854.4]
  wire  _T_1511; // @[MemPrimitives.scala 110:228:@10858.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@10872.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@10873.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@10874.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@10875.4]
  wire  _T_1517; // @[MemPrimitives.scala 123:41:@10876.4]
  wire  _T_1518; // @[MemPrimitives.scala 123:41:@10877.4]
  wire  _T_1519; // @[MemPrimitives.scala 123:41:@10878.4]
  wire  _T_1520; // @[MemPrimitives.scala 123:41:@10879.4]
  wire  _T_1521; // @[MemPrimitives.scala 123:41:@10880.4]
  wire [10:0] _T_1523; // @[Cat.scala 30:58:@10882.4]
  wire [10:0] _T_1525; // @[Cat.scala 30:58:@10884.4]
  wire [10:0] _T_1527; // @[Cat.scala 30:58:@10886.4]
  wire [10:0] _T_1529; // @[Cat.scala 30:58:@10888.4]
  wire [10:0] _T_1531; // @[Cat.scala 30:58:@10890.4]
  wire [10:0] _T_1533; // @[Cat.scala 30:58:@10892.4]
  wire [10:0] _T_1535; // @[Cat.scala 30:58:@10894.4]
  wire [10:0] _T_1537; // @[Cat.scala 30:58:@10896.4]
  wire [10:0] _T_1539; // @[Cat.scala 30:58:@10898.4]
  wire [10:0] _T_1540; // @[Mux.scala 31:69:@10899.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@10900.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@10901.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@10902.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@10903.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@10904.4]
  wire [10:0] _T_1546; // @[Mux.scala 31:69:@10905.4]
  wire [10:0] _T_1547; // @[Mux.scala 31:69:@10906.4]
  wire  _T_1643; // @[package.scala 96:25:@11035.4 package.scala 96:25:@11036.4]
  wire [7:0] _T_1647; // @[Mux.scala 31:69:@11045.4]
  wire  _T_1640; // @[package.scala 96:25:@11027.4 package.scala 96:25:@11028.4]
  wire [7:0] _T_1648; // @[Mux.scala 31:69:@11046.4]
  wire  _T_1637; // @[package.scala 96:25:@11019.4 package.scala 96:25:@11020.4]
  wire [7:0] _T_1649; // @[Mux.scala 31:69:@11047.4]
  wire  _T_1634; // @[package.scala 96:25:@11011.4 package.scala 96:25:@11012.4]
  wire [7:0] _T_1650; // @[Mux.scala 31:69:@11048.4]
  wire  _T_1631; // @[package.scala 96:25:@11003.4 package.scala 96:25:@11004.4]
  wire [7:0] _T_1651; // @[Mux.scala 31:69:@11049.4]
  wire  _T_1628; // @[package.scala 96:25:@10995.4 package.scala 96:25:@10996.4]
  wire [7:0] _T_1652; // @[Mux.scala 31:69:@11050.4]
  wire  _T_1625; // @[package.scala 96:25:@10987.4 package.scala 96:25:@10988.4]
  wire [7:0] _T_1653; // @[Mux.scala 31:69:@11051.4]
  wire  _T_1622; // @[package.scala 96:25:@10979.4 package.scala 96:25:@10980.4]
  wire [7:0] _T_1654; // @[Mux.scala 31:69:@11052.4]
  wire  _T_1619; // @[package.scala 96:25:@10971.4 package.scala 96:25:@10972.4]
  wire [7:0] _T_1655; // @[Mux.scala 31:69:@11053.4]
  wire  _T_1616; // @[package.scala 96:25:@10963.4 package.scala 96:25:@10964.4]
  wire [7:0] _T_1656; // @[Mux.scala 31:69:@11054.4]
  wire  _T_1613; // @[package.scala 96:25:@10955.4 package.scala 96:25:@10956.4]
  wire  _T_1750; // @[package.scala 96:25:@11179.4 package.scala 96:25:@11180.4]
  wire [7:0] _T_1754; // @[Mux.scala 31:69:@11189.4]
  wire  _T_1747; // @[package.scala 96:25:@11171.4 package.scala 96:25:@11172.4]
  wire [7:0] _T_1755; // @[Mux.scala 31:69:@11190.4]
  wire  _T_1744; // @[package.scala 96:25:@11163.4 package.scala 96:25:@11164.4]
  wire [7:0] _T_1756; // @[Mux.scala 31:69:@11191.4]
  wire  _T_1741; // @[package.scala 96:25:@11155.4 package.scala 96:25:@11156.4]
  wire [7:0] _T_1757; // @[Mux.scala 31:69:@11192.4]
  wire  _T_1738; // @[package.scala 96:25:@11147.4 package.scala 96:25:@11148.4]
  wire [7:0] _T_1758; // @[Mux.scala 31:69:@11193.4]
  wire  _T_1735; // @[package.scala 96:25:@11139.4 package.scala 96:25:@11140.4]
  wire [7:0] _T_1759; // @[Mux.scala 31:69:@11194.4]
  wire  _T_1732; // @[package.scala 96:25:@11131.4 package.scala 96:25:@11132.4]
  wire [7:0] _T_1760; // @[Mux.scala 31:69:@11195.4]
  wire  _T_1729; // @[package.scala 96:25:@11123.4 package.scala 96:25:@11124.4]
  wire [7:0] _T_1761; // @[Mux.scala 31:69:@11196.4]
  wire  _T_1726; // @[package.scala 96:25:@11115.4 package.scala 96:25:@11116.4]
  wire [7:0] _T_1762; // @[Mux.scala 31:69:@11197.4]
  wire  _T_1723; // @[package.scala 96:25:@11107.4 package.scala 96:25:@11108.4]
  wire [7:0] _T_1763; // @[Mux.scala 31:69:@11198.4]
  wire  _T_1720; // @[package.scala 96:25:@11099.4 package.scala 96:25:@11100.4]
  wire  _T_1857; // @[package.scala 96:25:@11323.4 package.scala 96:25:@11324.4]
  wire [7:0] _T_1861; // @[Mux.scala 31:69:@11333.4]
  wire  _T_1854; // @[package.scala 96:25:@11315.4 package.scala 96:25:@11316.4]
  wire [7:0] _T_1862; // @[Mux.scala 31:69:@11334.4]
  wire  _T_1851; // @[package.scala 96:25:@11307.4 package.scala 96:25:@11308.4]
  wire [7:0] _T_1863; // @[Mux.scala 31:69:@11335.4]
  wire  _T_1848; // @[package.scala 96:25:@11299.4 package.scala 96:25:@11300.4]
  wire [7:0] _T_1864; // @[Mux.scala 31:69:@11336.4]
  wire  _T_1845; // @[package.scala 96:25:@11291.4 package.scala 96:25:@11292.4]
  wire [7:0] _T_1865; // @[Mux.scala 31:69:@11337.4]
  wire  _T_1842; // @[package.scala 96:25:@11283.4 package.scala 96:25:@11284.4]
  wire [7:0] _T_1866; // @[Mux.scala 31:69:@11338.4]
  wire  _T_1839; // @[package.scala 96:25:@11275.4 package.scala 96:25:@11276.4]
  wire [7:0] _T_1867; // @[Mux.scala 31:69:@11339.4]
  wire  _T_1836; // @[package.scala 96:25:@11267.4 package.scala 96:25:@11268.4]
  wire [7:0] _T_1868; // @[Mux.scala 31:69:@11340.4]
  wire  _T_1833; // @[package.scala 96:25:@11259.4 package.scala 96:25:@11260.4]
  wire [7:0] _T_1869; // @[Mux.scala 31:69:@11341.4]
  wire  _T_1830; // @[package.scala 96:25:@11251.4 package.scala 96:25:@11252.4]
  wire [7:0] _T_1870; // @[Mux.scala 31:69:@11342.4]
  wire  _T_1827; // @[package.scala 96:25:@11243.4 package.scala 96:25:@11244.4]
  wire  _T_1964; // @[package.scala 96:25:@11467.4 package.scala 96:25:@11468.4]
  wire [7:0] _T_1968; // @[Mux.scala 31:69:@11477.4]
  wire  _T_1961; // @[package.scala 96:25:@11459.4 package.scala 96:25:@11460.4]
  wire [7:0] _T_1969; // @[Mux.scala 31:69:@11478.4]
  wire  _T_1958; // @[package.scala 96:25:@11451.4 package.scala 96:25:@11452.4]
  wire [7:0] _T_1970; // @[Mux.scala 31:69:@11479.4]
  wire  _T_1955; // @[package.scala 96:25:@11443.4 package.scala 96:25:@11444.4]
  wire [7:0] _T_1971; // @[Mux.scala 31:69:@11480.4]
  wire  _T_1952; // @[package.scala 96:25:@11435.4 package.scala 96:25:@11436.4]
  wire [7:0] _T_1972; // @[Mux.scala 31:69:@11481.4]
  wire  _T_1949; // @[package.scala 96:25:@11427.4 package.scala 96:25:@11428.4]
  wire [7:0] _T_1973; // @[Mux.scala 31:69:@11482.4]
  wire  _T_1946; // @[package.scala 96:25:@11419.4 package.scala 96:25:@11420.4]
  wire [7:0] _T_1974; // @[Mux.scala 31:69:@11483.4]
  wire  _T_1943; // @[package.scala 96:25:@11411.4 package.scala 96:25:@11412.4]
  wire [7:0] _T_1975; // @[Mux.scala 31:69:@11484.4]
  wire  _T_1940; // @[package.scala 96:25:@11403.4 package.scala 96:25:@11404.4]
  wire [7:0] _T_1976; // @[Mux.scala 31:69:@11485.4]
  wire  _T_1937; // @[package.scala 96:25:@11395.4 package.scala 96:25:@11396.4]
  wire [7:0] _T_1977; // @[Mux.scala 31:69:@11486.4]
  wire  _T_1934; // @[package.scala 96:25:@11387.4 package.scala 96:25:@11388.4]
  wire  _T_2071; // @[package.scala 96:25:@11611.4 package.scala 96:25:@11612.4]
  wire [7:0] _T_2075; // @[Mux.scala 31:69:@11621.4]
  wire  _T_2068; // @[package.scala 96:25:@11603.4 package.scala 96:25:@11604.4]
  wire [7:0] _T_2076; // @[Mux.scala 31:69:@11622.4]
  wire  _T_2065; // @[package.scala 96:25:@11595.4 package.scala 96:25:@11596.4]
  wire [7:0] _T_2077; // @[Mux.scala 31:69:@11623.4]
  wire  _T_2062; // @[package.scala 96:25:@11587.4 package.scala 96:25:@11588.4]
  wire [7:0] _T_2078; // @[Mux.scala 31:69:@11624.4]
  wire  _T_2059; // @[package.scala 96:25:@11579.4 package.scala 96:25:@11580.4]
  wire [7:0] _T_2079; // @[Mux.scala 31:69:@11625.4]
  wire  _T_2056; // @[package.scala 96:25:@11571.4 package.scala 96:25:@11572.4]
  wire [7:0] _T_2080; // @[Mux.scala 31:69:@11626.4]
  wire  _T_2053; // @[package.scala 96:25:@11563.4 package.scala 96:25:@11564.4]
  wire [7:0] _T_2081; // @[Mux.scala 31:69:@11627.4]
  wire  _T_2050; // @[package.scala 96:25:@11555.4 package.scala 96:25:@11556.4]
  wire [7:0] _T_2082; // @[Mux.scala 31:69:@11628.4]
  wire  _T_2047; // @[package.scala 96:25:@11547.4 package.scala 96:25:@11548.4]
  wire [7:0] _T_2083; // @[Mux.scala 31:69:@11629.4]
  wire  _T_2044; // @[package.scala 96:25:@11539.4 package.scala 96:25:@11540.4]
  wire [7:0] _T_2084; // @[Mux.scala 31:69:@11630.4]
  wire  _T_2041; // @[package.scala 96:25:@11531.4 package.scala 96:25:@11532.4]
  wire  _T_2178; // @[package.scala 96:25:@11755.4 package.scala 96:25:@11756.4]
  wire [7:0] _T_2182; // @[Mux.scala 31:69:@11765.4]
  wire  _T_2175; // @[package.scala 96:25:@11747.4 package.scala 96:25:@11748.4]
  wire [7:0] _T_2183; // @[Mux.scala 31:69:@11766.4]
  wire  _T_2172; // @[package.scala 96:25:@11739.4 package.scala 96:25:@11740.4]
  wire [7:0] _T_2184; // @[Mux.scala 31:69:@11767.4]
  wire  _T_2169; // @[package.scala 96:25:@11731.4 package.scala 96:25:@11732.4]
  wire [7:0] _T_2185; // @[Mux.scala 31:69:@11768.4]
  wire  _T_2166; // @[package.scala 96:25:@11723.4 package.scala 96:25:@11724.4]
  wire [7:0] _T_2186; // @[Mux.scala 31:69:@11769.4]
  wire  _T_2163; // @[package.scala 96:25:@11715.4 package.scala 96:25:@11716.4]
  wire [7:0] _T_2187; // @[Mux.scala 31:69:@11770.4]
  wire  _T_2160; // @[package.scala 96:25:@11707.4 package.scala 96:25:@11708.4]
  wire [7:0] _T_2188; // @[Mux.scala 31:69:@11771.4]
  wire  _T_2157; // @[package.scala 96:25:@11699.4 package.scala 96:25:@11700.4]
  wire [7:0] _T_2189; // @[Mux.scala 31:69:@11772.4]
  wire  _T_2154; // @[package.scala 96:25:@11691.4 package.scala 96:25:@11692.4]
  wire [7:0] _T_2190; // @[Mux.scala 31:69:@11773.4]
  wire  _T_2151; // @[package.scala 96:25:@11683.4 package.scala 96:25:@11684.4]
  wire [7:0] _T_2191; // @[Mux.scala 31:69:@11774.4]
  wire  _T_2148; // @[package.scala 96:25:@11675.4 package.scala 96:25:@11676.4]
  wire  _T_2285; // @[package.scala 96:25:@11899.4 package.scala 96:25:@11900.4]
  wire [7:0] _T_2289; // @[Mux.scala 31:69:@11909.4]
  wire  _T_2282; // @[package.scala 96:25:@11891.4 package.scala 96:25:@11892.4]
  wire [7:0] _T_2290; // @[Mux.scala 31:69:@11910.4]
  wire  _T_2279; // @[package.scala 96:25:@11883.4 package.scala 96:25:@11884.4]
  wire [7:0] _T_2291; // @[Mux.scala 31:69:@11911.4]
  wire  _T_2276; // @[package.scala 96:25:@11875.4 package.scala 96:25:@11876.4]
  wire [7:0] _T_2292; // @[Mux.scala 31:69:@11912.4]
  wire  _T_2273; // @[package.scala 96:25:@11867.4 package.scala 96:25:@11868.4]
  wire [7:0] _T_2293; // @[Mux.scala 31:69:@11913.4]
  wire  _T_2270; // @[package.scala 96:25:@11859.4 package.scala 96:25:@11860.4]
  wire [7:0] _T_2294; // @[Mux.scala 31:69:@11914.4]
  wire  _T_2267; // @[package.scala 96:25:@11851.4 package.scala 96:25:@11852.4]
  wire [7:0] _T_2295; // @[Mux.scala 31:69:@11915.4]
  wire  _T_2264; // @[package.scala 96:25:@11843.4 package.scala 96:25:@11844.4]
  wire [7:0] _T_2296; // @[Mux.scala 31:69:@11916.4]
  wire  _T_2261; // @[package.scala 96:25:@11835.4 package.scala 96:25:@11836.4]
  wire [7:0] _T_2297; // @[Mux.scala 31:69:@11917.4]
  wire  _T_2258; // @[package.scala 96:25:@11827.4 package.scala 96:25:@11828.4]
  wire [7:0] _T_2298; // @[Mux.scala 31:69:@11918.4]
  wire  _T_2255; // @[package.scala 96:25:@11819.4 package.scala 96:25:@11820.4]
  wire  _T_2392; // @[package.scala 96:25:@12043.4 package.scala 96:25:@12044.4]
  wire [7:0] _T_2396; // @[Mux.scala 31:69:@12053.4]
  wire  _T_2389; // @[package.scala 96:25:@12035.4 package.scala 96:25:@12036.4]
  wire [7:0] _T_2397; // @[Mux.scala 31:69:@12054.4]
  wire  _T_2386; // @[package.scala 96:25:@12027.4 package.scala 96:25:@12028.4]
  wire [7:0] _T_2398; // @[Mux.scala 31:69:@12055.4]
  wire  _T_2383; // @[package.scala 96:25:@12019.4 package.scala 96:25:@12020.4]
  wire [7:0] _T_2399; // @[Mux.scala 31:69:@12056.4]
  wire  _T_2380; // @[package.scala 96:25:@12011.4 package.scala 96:25:@12012.4]
  wire [7:0] _T_2400; // @[Mux.scala 31:69:@12057.4]
  wire  _T_2377; // @[package.scala 96:25:@12003.4 package.scala 96:25:@12004.4]
  wire [7:0] _T_2401; // @[Mux.scala 31:69:@12058.4]
  wire  _T_2374; // @[package.scala 96:25:@11995.4 package.scala 96:25:@11996.4]
  wire [7:0] _T_2402; // @[Mux.scala 31:69:@12059.4]
  wire  _T_2371; // @[package.scala 96:25:@11987.4 package.scala 96:25:@11988.4]
  wire [7:0] _T_2403; // @[Mux.scala 31:69:@12060.4]
  wire  _T_2368; // @[package.scala 96:25:@11979.4 package.scala 96:25:@11980.4]
  wire [7:0] _T_2404; // @[Mux.scala 31:69:@12061.4]
  wire  _T_2365; // @[package.scala 96:25:@11971.4 package.scala 96:25:@11972.4]
  wire [7:0] _T_2405; // @[Mux.scala 31:69:@12062.4]
  wire  _T_2362; // @[package.scala 96:25:@11963.4 package.scala 96:25:@11964.4]
  wire  _T_2499; // @[package.scala 96:25:@12187.4 package.scala 96:25:@12188.4]
  wire [7:0] _T_2503; // @[Mux.scala 31:69:@12197.4]
  wire  _T_2496; // @[package.scala 96:25:@12179.4 package.scala 96:25:@12180.4]
  wire [7:0] _T_2504; // @[Mux.scala 31:69:@12198.4]
  wire  _T_2493; // @[package.scala 96:25:@12171.4 package.scala 96:25:@12172.4]
  wire [7:0] _T_2505; // @[Mux.scala 31:69:@12199.4]
  wire  _T_2490; // @[package.scala 96:25:@12163.4 package.scala 96:25:@12164.4]
  wire [7:0] _T_2506; // @[Mux.scala 31:69:@12200.4]
  wire  _T_2487; // @[package.scala 96:25:@12155.4 package.scala 96:25:@12156.4]
  wire [7:0] _T_2507; // @[Mux.scala 31:69:@12201.4]
  wire  _T_2484; // @[package.scala 96:25:@12147.4 package.scala 96:25:@12148.4]
  wire [7:0] _T_2508; // @[Mux.scala 31:69:@12202.4]
  wire  _T_2481; // @[package.scala 96:25:@12139.4 package.scala 96:25:@12140.4]
  wire [7:0] _T_2509; // @[Mux.scala 31:69:@12203.4]
  wire  _T_2478; // @[package.scala 96:25:@12131.4 package.scala 96:25:@12132.4]
  wire [7:0] _T_2510; // @[Mux.scala 31:69:@12204.4]
  wire  _T_2475; // @[package.scala 96:25:@12123.4 package.scala 96:25:@12124.4]
  wire [7:0] _T_2511; // @[Mux.scala 31:69:@12205.4]
  wire  _T_2472; // @[package.scala 96:25:@12115.4 package.scala 96:25:@12116.4]
  wire [7:0] _T_2512; // @[Mux.scala 31:69:@12206.4]
  wire  _T_2469; // @[package.scala 96:25:@12107.4 package.scala 96:25:@12108.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@9509.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@9525.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@9541.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@9557.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@9573.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@9589.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@9605.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@9621.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@9637.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@9653.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@9669.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@9685.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@9881.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@9970.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@10059.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@10148.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@10237.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@10326.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@10415.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@10504.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@10593.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@10682.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects StickySelects_10 ( // @[MemPrimitives.scala 121:29:@10771.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects StickySelects_11 ( // @[MemPrimitives.scala 121:29:@10860.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  RetimeWrapper_32 RetimeWrapper ( // @[package.scala 93:22:@10950.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_1 ( // @[package.scala 93:22:@10958.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_2 ( // @[package.scala 93:22:@10966.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_3 ( // @[package.scala 93:22:@10974.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_4 ( // @[package.scala 93:22:@10982.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_5 ( // @[package.scala 93:22:@10990.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_6 ( // @[package.scala 93:22:@10998.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_7 ( // @[package.scala 93:22:@11006.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_8 ( // @[package.scala 93:22:@11014.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_9 ( // @[package.scala 93:22:@11022.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_10 ( // @[package.scala 93:22:@11030.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_11 ( // @[package.scala 93:22:@11038.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_12 ( // @[package.scala 93:22:@11094.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_13 ( // @[package.scala 93:22:@11102.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_14 ( // @[package.scala 93:22:@11110.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_15 ( // @[package.scala 93:22:@11118.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_16 ( // @[package.scala 93:22:@11126.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_17 ( // @[package.scala 93:22:@11134.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_18 ( // @[package.scala 93:22:@11142.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_19 ( // @[package.scala 93:22:@11150.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_20 ( // @[package.scala 93:22:@11158.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_21 ( // @[package.scala 93:22:@11166.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_22 ( // @[package.scala 93:22:@11174.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_23 ( // @[package.scala 93:22:@11182.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_24 ( // @[package.scala 93:22:@11238.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_25 ( // @[package.scala 93:22:@11246.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_26 ( // @[package.scala 93:22:@11254.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_27 ( // @[package.scala 93:22:@11262.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_28 ( // @[package.scala 93:22:@11270.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_29 ( // @[package.scala 93:22:@11278.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_30 ( // @[package.scala 93:22:@11286.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_31 ( // @[package.scala 93:22:@11294.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_32 ( // @[package.scala 93:22:@11302.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_33 ( // @[package.scala 93:22:@11310.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_34 ( // @[package.scala 93:22:@11318.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_35 ( // @[package.scala 93:22:@11326.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_36 ( // @[package.scala 93:22:@11382.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_37 ( // @[package.scala 93:22:@11390.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_38 ( // @[package.scala 93:22:@11398.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_39 ( // @[package.scala 93:22:@11406.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_40 ( // @[package.scala 93:22:@11414.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_41 ( // @[package.scala 93:22:@11422.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_42 ( // @[package.scala 93:22:@11430.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_43 ( // @[package.scala 93:22:@11438.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_44 ( // @[package.scala 93:22:@11446.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_45 ( // @[package.scala 93:22:@11454.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_46 ( // @[package.scala 93:22:@11462.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_47 ( // @[package.scala 93:22:@11470.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_48 ( // @[package.scala 93:22:@11526.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_49 ( // @[package.scala 93:22:@11534.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_50 ( // @[package.scala 93:22:@11542.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_51 ( // @[package.scala 93:22:@11550.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_52 ( // @[package.scala 93:22:@11558.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_53 ( // @[package.scala 93:22:@11566.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_54 ( // @[package.scala 93:22:@11574.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_55 ( // @[package.scala 93:22:@11582.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_56 ( // @[package.scala 93:22:@11590.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_57 ( // @[package.scala 93:22:@11598.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_58 ( // @[package.scala 93:22:@11606.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_59 ( // @[package.scala 93:22:@11614.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_60 ( // @[package.scala 93:22:@11670.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_61 ( // @[package.scala 93:22:@11678.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_62 ( // @[package.scala 93:22:@11686.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_63 ( // @[package.scala 93:22:@11694.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_64 ( // @[package.scala 93:22:@11702.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_65 ( // @[package.scala 93:22:@11710.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_66 ( // @[package.scala 93:22:@11718.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_67 ( // @[package.scala 93:22:@11726.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_68 ( // @[package.scala 93:22:@11734.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_69 ( // @[package.scala 93:22:@11742.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_70 ( // @[package.scala 93:22:@11750.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_71 ( // @[package.scala 93:22:@11758.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_72 ( // @[package.scala 93:22:@11814.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_73 ( // @[package.scala 93:22:@11822.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_74 ( // @[package.scala 93:22:@11830.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_75 ( // @[package.scala 93:22:@11838.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_76 ( // @[package.scala 93:22:@11846.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_77 ( // @[package.scala 93:22:@11854.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_78 ( // @[package.scala 93:22:@11862.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_79 ( // @[package.scala 93:22:@11870.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_80 ( // @[package.scala 93:22:@11878.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_81 ( // @[package.scala 93:22:@11886.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_82 ( // @[package.scala 93:22:@11894.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_83 ( // @[package.scala 93:22:@11902.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_84 ( // @[package.scala 93:22:@11958.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_85 ( // @[package.scala 93:22:@11966.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_86 ( // @[package.scala 93:22:@11974.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_87 ( // @[package.scala 93:22:@11982.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_88 ( // @[package.scala 93:22:@11990.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_89 ( // @[package.scala 93:22:@11998.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_90 ( // @[package.scala 93:22:@12006.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_91 ( // @[package.scala 93:22:@12014.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_92 ( // @[package.scala 93:22:@12022.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_93 ( // @[package.scala 93:22:@12030.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_94 ( // @[package.scala 93:22:@12038.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_95 ( // @[package.scala 93:22:@12046.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_96 ( // @[package.scala 93:22:@12102.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_97 ( // @[package.scala 93:22:@12110.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_98 ( // @[package.scala 93:22:@12118.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_99 ( // @[package.scala 93:22:@12126.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_100 ( // @[package.scala 93:22:@12134.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_101 ( // @[package.scala 93:22:@12142.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_102 ( // @[package.scala 93:22:@12150.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_103 ( // @[package.scala 93:22:@12158.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_104 ( // @[package.scala 93:22:@12166.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_105 ( // @[package.scala 93:22:@12174.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_106 ( // @[package.scala 93:22:@12182.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_107 ( // @[package.scala 93:22:@12190.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  assign _T_316 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9701.4]
  assign _T_318 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@9702.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 82:228:@9703.4]
  assign _T_320 = io_wPort_0_en_0 & _T_319; // @[MemPrimitives.scala 83:102:@9704.4]
  assign _T_322 = {_T_320,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9706.4]
  assign _T_329 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@9714.4]
  assign _T_330 = _T_316 & _T_329; // @[MemPrimitives.scala 82:228:@9715.4]
  assign _T_331 = io_wPort_0_en_0 & _T_330; // @[MemPrimitives.scala 83:102:@9716.4]
  assign _T_333 = {_T_331,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9718.4]
  assign _T_340 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@9726.4]
  assign _T_341 = _T_316 & _T_340; // @[MemPrimitives.scala 82:228:@9727.4]
  assign _T_342 = io_wPort_0_en_0 & _T_341; // @[MemPrimitives.scala 83:102:@9728.4]
  assign _T_344 = {_T_342,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9730.4]
  assign _T_349 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9737.4]
  assign _T_352 = _T_349 & _T_318; // @[MemPrimitives.scala 82:228:@9739.4]
  assign _T_353 = io_wPort_0_en_0 & _T_352; // @[MemPrimitives.scala 83:102:@9740.4]
  assign _T_355 = {_T_353,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9742.4]
  assign _T_363 = _T_349 & _T_329; // @[MemPrimitives.scala 82:228:@9751.4]
  assign _T_364 = io_wPort_0_en_0 & _T_363; // @[MemPrimitives.scala 83:102:@9752.4]
  assign _T_366 = {_T_364,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9754.4]
  assign _T_374 = _T_349 & _T_340; // @[MemPrimitives.scala 82:228:@9763.4]
  assign _T_375 = io_wPort_0_en_0 & _T_374; // @[MemPrimitives.scala 83:102:@9764.4]
  assign _T_377 = {_T_375,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9766.4]
  assign _T_382 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9773.4]
  assign _T_385 = _T_382 & _T_318; // @[MemPrimitives.scala 82:228:@9775.4]
  assign _T_386 = io_wPort_0_en_0 & _T_385; // @[MemPrimitives.scala 83:102:@9776.4]
  assign _T_388 = {_T_386,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9778.4]
  assign _T_396 = _T_382 & _T_329; // @[MemPrimitives.scala 82:228:@9787.4]
  assign _T_397 = io_wPort_0_en_0 & _T_396; // @[MemPrimitives.scala 83:102:@9788.4]
  assign _T_399 = {_T_397,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9790.4]
  assign _T_407 = _T_382 & _T_340; // @[MemPrimitives.scala 82:228:@9799.4]
  assign _T_408 = io_wPort_0_en_0 & _T_407; // @[MemPrimitives.scala 83:102:@9800.4]
  assign _T_410 = {_T_408,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9802.4]
  assign _T_415 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9809.4]
  assign _T_418 = _T_415 & _T_318; // @[MemPrimitives.scala 82:228:@9811.4]
  assign _T_419 = io_wPort_0_en_0 & _T_418; // @[MemPrimitives.scala 83:102:@9812.4]
  assign _T_421 = {_T_419,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9814.4]
  assign _T_429 = _T_415 & _T_329; // @[MemPrimitives.scala 82:228:@9823.4]
  assign _T_430 = io_wPort_0_en_0 & _T_429; // @[MemPrimitives.scala 83:102:@9824.4]
  assign _T_432 = {_T_430,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9826.4]
  assign _T_440 = _T_415 & _T_340; // @[MemPrimitives.scala 82:228:@9835.4]
  assign _T_441 = io_wPort_0_en_0 & _T_440; // @[MemPrimitives.scala 83:102:@9836.4]
  assign _T_443 = {_T_441,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9838.4]
  assign _T_448 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9845.4]
  assign _T_450 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9846.4]
  assign _T_451 = _T_448 & _T_450; // @[MemPrimitives.scala 110:228:@9847.4]
  assign _T_454 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9849.4]
  assign _T_456 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9850.4]
  assign _T_457 = _T_454 & _T_456; // @[MemPrimitives.scala 110:228:@9851.4]
  assign _T_460 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9853.4]
  assign _T_462 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9854.4]
  assign _T_463 = _T_460 & _T_462; // @[MemPrimitives.scala 110:228:@9855.4]
  assign _T_466 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9857.4]
  assign _T_468 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9858.4]
  assign _T_469 = _T_466 & _T_468; // @[MemPrimitives.scala 110:228:@9859.4]
  assign _T_472 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9861.4]
  assign _T_474 = io_rPort_4_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9862.4]
  assign _T_475 = _T_472 & _T_474; // @[MemPrimitives.scala 110:228:@9863.4]
  assign _T_478 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9865.4]
  assign _T_480 = io_rPort_5_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9866.4]
  assign _T_481 = _T_478 & _T_480; // @[MemPrimitives.scala 110:228:@9867.4]
  assign _T_484 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9869.4]
  assign _T_486 = io_rPort_6_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9870.4]
  assign _T_487 = _T_484 & _T_486; // @[MemPrimitives.scala 110:228:@9871.4]
  assign _T_490 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9873.4]
  assign _T_492 = io_rPort_7_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9874.4]
  assign _T_493 = _T_490 & _T_492; // @[MemPrimitives.scala 110:228:@9875.4]
  assign _T_496 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9877.4]
  assign _T_498 = io_rPort_8_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@9878.4]
  assign _T_499 = _T_496 & _T_498; // @[MemPrimitives.scala 110:228:@9879.4]
  assign _T_501 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@9893.4]
  assign _T_502 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@9894.4]
  assign _T_503 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@9895.4]
  assign _T_504 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@9896.4]
  assign _T_505 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@9897.4]
  assign _T_506 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@9898.4]
  assign _T_507 = StickySelects_io_outs_6; // @[MemPrimitives.scala 123:41:@9899.4]
  assign _T_508 = StickySelects_io_outs_7; // @[MemPrimitives.scala 123:41:@9900.4]
  assign _T_509 = StickySelects_io_outs_8; // @[MemPrimitives.scala 123:41:@9901.4]
  assign _T_511 = {_T_501,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9903.4]
  assign _T_513 = {_T_502,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9905.4]
  assign _T_515 = {_T_503,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9907.4]
  assign _T_517 = {_T_504,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9909.4]
  assign _T_519 = {_T_505,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9911.4]
  assign _T_521 = {_T_506,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9913.4]
  assign _T_523 = {_T_507,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9915.4]
  assign _T_525 = {_T_508,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9917.4]
  assign _T_527 = {_T_509,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9919.4]
  assign _T_528 = _T_508 ? _T_525 : _T_527; // @[Mux.scala 31:69:@9920.4]
  assign _T_529 = _T_507 ? _T_523 : _T_528; // @[Mux.scala 31:69:@9921.4]
  assign _T_530 = _T_506 ? _T_521 : _T_529; // @[Mux.scala 31:69:@9922.4]
  assign _T_531 = _T_505 ? _T_519 : _T_530; // @[Mux.scala 31:69:@9923.4]
  assign _T_532 = _T_504 ? _T_517 : _T_531; // @[Mux.scala 31:69:@9924.4]
  assign _T_533 = _T_503 ? _T_515 : _T_532; // @[Mux.scala 31:69:@9925.4]
  assign _T_534 = _T_502 ? _T_513 : _T_533; // @[Mux.scala 31:69:@9926.4]
  assign _T_535 = _T_501 ? _T_511 : _T_534; // @[Mux.scala 31:69:@9927.4]
  assign _T_542 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9935.4]
  assign _T_543 = _T_448 & _T_542; // @[MemPrimitives.scala 110:228:@9936.4]
  assign _T_548 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9939.4]
  assign _T_549 = _T_454 & _T_548; // @[MemPrimitives.scala 110:228:@9940.4]
  assign _T_554 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9943.4]
  assign _T_555 = _T_460 & _T_554; // @[MemPrimitives.scala 110:228:@9944.4]
  assign _T_560 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9947.4]
  assign _T_561 = _T_466 & _T_560; // @[MemPrimitives.scala 110:228:@9948.4]
  assign _T_566 = io_rPort_4_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9951.4]
  assign _T_567 = _T_472 & _T_566; // @[MemPrimitives.scala 110:228:@9952.4]
  assign _T_572 = io_rPort_5_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9955.4]
  assign _T_573 = _T_478 & _T_572; // @[MemPrimitives.scala 110:228:@9956.4]
  assign _T_578 = io_rPort_6_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9959.4]
  assign _T_579 = _T_484 & _T_578; // @[MemPrimitives.scala 110:228:@9960.4]
  assign _T_584 = io_rPort_7_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9963.4]
  assign _T_585 = _T_490 & _T_584; // @[MemPrimitives.scala 110:228:@9964.4]
  assign _T_590 = io_rPort_8_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@9967.4]
  assign _T_591 = _T_496 & _T_590; // @[MemPrimitives.scala 110:228:@9968.4]
  assign _T_593 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@9982.4]
  assign _T_594 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@9983.4]
  assign _T_595 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@9984.4]
  assign _T_596 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@9985.4]
  assign _T_597 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@9986.4]
  assign _T_598 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@9987.4]
  assign _T_599 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 123:41:@9988.4]
  assign _T_600 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 123:41:@9989.4]
  assign _T_601 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 123:41:@9990.4]
  assign _T_603 = {_T_593,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9992.4]
  assign _T_605 = {_T_594,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9994.4]
  assign _T_607 = {_T_595,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9996.4]
  assign _T_609 = {_T_596,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9998.4]
  assign _T_611 = {_T_597,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10000.4]
  assign _T_613 = {_T_598,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10002.4]
  assign _T_615 = {_T_599,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10004.4]
  assign _T_617 = {_T_600,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10006.4]
  assign _T_619 = {_T_601,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10008.4]
  assign _T_620 = _T_600 ? _T_617 : _T_619; // @[Mux.scala 31:69:@10009.4]
  assign _T_621 = _T_599 ? _T_615 : _T_620; // @[Mux.scala 31:69:@10010.4]
  assign _T_622 = _T_598 ? _T_613 : _T_621; // @[Mux.scala 31:69:@10011.4]
  assign _T_623 = _T_597 ? _T_611 : _T_622; // @[Mux.scala 31:69:@10012.4]
  assign _T_624 = _T_596 ? _T_609 : _T_623; // @[Mux.scala 31:69:@10013.4]
  assign _T_625 = _T_595 ? _T_607 : _T_624; // @[Mux.scala 31:69:@10014.4]
  assign _T_626 = _T_594 ? _T_605 : _T_625; // @[Mux.scala 31:69:@10015.4]
  assign _T_627 = _T_593 ? _T_603 : _T_626; // @[Mux.scala 31:69:@10016.4]
  assign _T_634 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10024.4]
  assign _T_635 = _T_448 & _T_634; // @[MemPrimitives.scala 110:228:@10025.4]
  assign _T_640 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10028.4]
  assign _T_641 = _T_454 & _T_640; // @[MemPrimitives.scala 110:228:@10029.4]
  assign _T_646 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10032.4]
  assign _T_647 = _T_460 & _T_646; // @[MemPrimitives.scala 110:228:@10033.4]
  assign _T_652 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10036.4]
  assign _T_653 = _T_466 & _T_652; // @[MemPrimitives.scala 110:228:@10037.4]
  assign _T_658 = io_rPort_4_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10040.4]
  assign _T_659 = _T_472 & _T_658; // @[MemPrimitives.scala 110:228:@10041.4]
  assign _T_664 = io_rPort_5_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10044.4]
  assign _T_665 = _T_478 & _T_664; // @[MemPrimitives.scala 110:228:@10045.4]
  assign _T_670 = io_rPort_6_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10048.4]
  assign _T_671 = _T_484 & _T_670; // @[MemPrimitives.scala 110:228:@10049.4]
  assign _T_676 = io_rPort_7_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10052.4]
  assign _T_677 = _T_490 & _T_676; // @[MemPrimitives.scala 110:228:@10053.4]
  assign _T_682 = io_rPort_8_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@10056.4]
  assign _T_683 = _T_496 & _T_682; // @[MemPrimitives.scala 110:228:@10057.4]
  assign _T_685 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@10071.4]
  assign _T_686 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@10072.4]
  assign _T_687 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@10073.4]
  assign _T_688 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@10074.4]
  assign _T_689 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@10075.4]
  assign _T_690 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@10076.4]
  assign _T_691 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@10077.4]
  assign _T_692 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@10078.4]
  assign _T_693 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 123:41:@10079.4]
  assign _T_695 = {_T_685,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10081.4]
  assign _T_697 = {_T_686,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10083.4]
  assign _T_699 = {_T_687,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10085.4]
  assign _T_701 = {_T_688,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10087.4]
  assign _T_703 = {_T_689,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10089.4]
  assign _T_705 = {_T_690,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10091.4]
  assign _T_707 = {_T_691,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10093.4]
  assign _T_709 = {_T_692,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10095.4]
  assign _T_711 = {_T_693,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10097.4]
  assign _T_712 = _T_692 ? _T_709 : _T_711; // @[Mux.scala 31:69:@10098.4]
  assign _T_713 = _T_691 ? _T_707 : _T_712; // @[Mux.scala 31:69:@10099.4]
  assign _T_714 = _T_690 ? _T_705 : _T_713; // @[Mux.scala 31:69:@10100.4]
  assign _T_715 = _T_689 ? _T_703 : _T_714; // @[Mux.scala 31:69:@10101.4]
  assign _T_716 = _T_688 ? _T_701 : _T_715; // @[Mux.scala 31:69:@10102.4]
  assign _T_717 = _T_687 ? _T_699 : _T_716; // @[Mux.scala 31:69:@10103.4]
  assign _T_718 = _T_686 ? _T_697 : _T_717; // @[Mux.scala 31:69:@10104.4]
  assign _T_719 = _T_685 ? _T_695 : _T_718; // @[Mux.scala 31:69:@10105.4]
  assign _T_724 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10112.4]
  assign _T_727 = _T_724 & _T_450; // @[MemPrimitives.scala 110:228:@10114.4]
  assign _T_730 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10116.4]
  assign _T_733 = _T_730 & _T_456; // @[MemPrimitives.scala 110:228:@10118.4]
  assign _T_736 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10120.4]
  assign _T_739 = _T_736 & _T_462; // @[MemPrimitives.scala 110:228:@10122.4]
  assign _T_742 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10124.4]
  assign _T_745 = _T_742 & _T_468; // @[MemPrimitives.scala 110:228:@10126.4]
  assign _T_748 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10128.4]
  assign _T_751 = _T_748 & _T_474; // @[MemPrimitives.scala 110:228:@10130.4]
  assign _T_754 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10132.4]
  assign _T_757 = _T_754 & _T_480; // @[MemPrimitives.scala 110:228:@10134.4]
  assign _T_760 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10136.4]
  assign _T_763 = _T_760 & _T_486; // @[MemPrimitives.scala 110:228:@10138.4]
  assign _T_766 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10140.4]
  assign _T_769 = _T_766 & _T_492; // @[MemPrimitives.scala 110:228:@10142.4]
  assign _T_772 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10144.4]
  assign _T_775 = _T_772 & _T_498; // @[MemPrimitives.scala 110:228:@10146.4]
  assign _T_777 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@10160.4]
  assign _T_778 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@10161.4]
  assign _T_779 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@10162.4]
  assign _T_780 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@10163.4]
  assign _T_781 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@10164.4]
  assign _T_782 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@10165.4]
  assign _T_783 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@10166.4]
  assign _T_784 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@10167.4]
  assign _T_785 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 123:41:@10168.4]
  assign _T_787 = {_T_777,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10170.4]
  assign _T_789 = {_T_778,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10172.4]
  assign _T_791 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10174.4]
  assign _T_793 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10176.4]
  assign _T_795 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10178.4]
  assign _T_797 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10180.4]
  assign _T_799 = {_T_783,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10182.4]
  assign _T_801 = {_T_784,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10184.4]
  assign _T_803 = {_T_785,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10186.4]
  assign _T_804 = _T_784 ? _T_801 : _T_803; // @[Mux.scala 31:69:@10187.4]
  assign _T_805 = _T_783 ? _T_799 : _T_804; // @[Mux.scala 31:69:@10188.4]
  assign _T_806 = _T_782 ? _T_797 : _T_805; // @[Mux.scala 31:69:@10189.4]
  assign _T_807 = _T_781 ? _T_795 : _T_806; // @[Mux.scala 31:69:@10190.4]
  assign _T_808 = _T_780 ? _T_793 : _T_807; // @[Mux.scala 31:69:@10191.4]
  assign _T_809 = _T_779 ? _T_791 : _T_808; // @[Mux.scala 31:69:@10192.4]
  assign _T_810 = _T_778 ? _T_789 : _T_809; // @[Mux.scala 31:69:@10193.4]
  assign _T_811 = _T_777 ? _T_787 : _T_810; // @[Mux.scala 31:69:@10194.4]
  assign _T_819 = _T_724 & _T_542; // @[MemPrimitives.scala 110:228:@10203.4]
  assign _T_825 = _T_730 & _T_548; // @[MemPrimitives.scala 110:228:@10207.4]
  assign _T_831 = _T_736 & _T_554; // @[MemPrimitives.scala 110:228:@10211.4]
  assign _T_837 = _T_742 & _T_560; // @[MemPrimitives.scala 110:228:@10215.4]
  assign _T_843 = _T_748 & _T_566; // @[MemPrimitives.scala 110:228:@10219.4]
  assign _T_849 = _T_754 & _T_572; // @[MemPrimitives.scala 110:228:@10223.4]
  assign _T_855 = _T_760 & _T_578; // @[MemPrimitives.scala 110:228:@10227.4]
  assign _T_861 = _T_766 & _T_584; // @[MemPrimitives.scala 110:228:@10231.4]
  assign _T_867 = _T_772 & _T_590; // @[MemPrimitives.scala 110:228:@10235.4]
  assign _T_869 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@10249.4]
  assign _T_870 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@10250.4]
  assign _T_871 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@10251.4]
  assign _T_872 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@10252.4]
  assign _T_873 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@10253.4]
  assign _T_874 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@10254.4]
  assign _T_875 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 123:41:@10255.4]
  assign _T_876 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 123:41:@10256.4]
  assign _T_877 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 123:41:@10257.4]
  assign _T_879 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10259.4]
  assign _T_881 = {_T_870,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10261.4]
  assign _T_883 = {_T_871,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10263.4]
  assign _T_885 = {_T_872,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10265.4]
  assign _T_887 = {_T_873,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10267.4]
  assign _T_889 = {_T_874,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10269.4]
  assign _T_891 = {_T_875,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10271.4]
  assign _T_893 = {_T_876,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10273.4]
  assign _T_895 = {_T_877,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10275.4]
  assign _T_896 = _T_876 ? _T_893 : _T_895; // @[Mux.scala 31:69:@10276.4]
  assign _T_897 = _T_875 ? _T_891 : _T_896; // @[Mux.scala 31:69:@10277.4]
  assign _T_898 = _T_874 ? _T_889 : _T_897; // @[Mux.scala 31:69:@10278.4]
  assign _T_899 = _T_873 ? _T_887 : _T_898; // @[Mux.scala 31:69:@10279.4]
  assign _T_900 = _T_872 ? _T_885 : _T_899; // @[Mux.scala 31:69:@10280.4]
  assign _T_901 = _T_871 ? _T_883 : _T_900; // @[Mux.scala 31:69:@10281.4]
  assign _T_902 = _T_870 ? _T_881 : _T_901; // @[Mux.scala 31:69:@10282.4]
  assign _T_903 = _T_869 ? _T_879 : _T_902; // @[Mux.scala 31:69:@10283.4]
  assign _T_911 = _T_724 & _T_634; // @[MemPrimitives.scala 110:228:@10292.4]
  assign _T_917 = _T_730 & _T_640; // @[MemPrimitives.scala 110:228:@10296.4]
  assign _T_923 = _T_736 & _T_646; // @[MemPrimitives.scala 110:228:@10300.4]
  assign _T_929 = _T_742 & _T_652; // @[MemPrimitives.scala 110:228:@10304.4]
  assign _T_935 = _T_748 & _T_658; // @[MemPrimitives.scala 110:228:@10308.4]
  assign _T_941 = _T_754 & _T_664; // @[MemPrimitives.scala 110:228:@10312.4]
  assign _T_947 = _T_760 & _T_670; // @[MemPrimitives.scala 110:228:@10316.4]
  assign _T_953 = _T_766 & _T_676; // @[MemPrimitives.scala 110:228:@10320.4]
  assign _T_959 = _T_772 & _T_682; // @[MemPrimitives.scala 110:228:@10324.4]
  assign _T_961 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@10338.4]
  assign _T_962 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@10339.4]
  assign _T_963 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@10340.4]
  assign _T_964 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@10341.4]
  assign _T_965 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@10342.4]
  assign _T_966 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@10343.4]
  assign _T_967 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 123:41:@10344.4]
  assign _T_968 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 123:41:@10345.4]
  assign _T_969 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 123:41:@10346.4]
  assign _T_971 = {_T_961,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10348.4]
  assign _T_973 = {_T_962,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10350.4]
  assign _T_975 = {_T_963,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10352.4]
  assign _T_977 = {_T_964,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10354.4]
  assign _T_979 = {_T_965,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10356.4]
  assign _T_981 = {_T_966,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10358.4]
  assign _T_983 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10360.4]
  assign _T_985 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10362.4]
  assign _T_987 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10364.4]
  assign _T_988 = _T_968 ? _T_985 : _T_987; // @[Mux.scala 31:69:@10365.4]
  assign _T_989 = _T_967 ? _T_983 : _T_988; // @[Mux.scala 31:69:@10366.4]
  assign _T_990 = _T_966 ? _T_981 : _T_989; // @[Mux.scala 31:69:@10367.4]
  assign _T_991 = _T_965 ? _T_979 : _T_990; // @[Mux.scala 31:69:@10368.4]
  assign _T_992 = _T_964 ? _T_977 : _T_991; // @[Mux.scala 31:69:@10369.4]
  assign _T_993 = _T_963 ? _T_975 : _T_992; // @[Mux.scala 31:69:@10370.4]
  assign _T_994 = _T_962 ? _T_973 : _T_993; // @[Mux.scala 31:69:@10371.4]
  assign _T_995 = _T_961 ? _T_971 : _T_994; // @[Mux.scala 31:69:@10372.4]
  assign _T_1000 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10379.4]
  assign _T_1003 = _T_1000 & _T_450; // @[MemPrimitives.scala 110:228:@10381.4]
  assign _T_1006 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10383.4]
  assign _T_1009 = _T_1006 & _T_456; // @[MemPrimitives.scala 110:228:@10385.4]
  assign _T_1012 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10387.4]
  assign _T_1015 = _T_1012 & _T_462; // @[MemPrimitives.scala 110:228:@10389.4]
  assign _T_1018 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10391.4]
  assign _T_1021 = _T_1018 & _T_468; // @[MemPrimitives.scala 110:228:@10393.4]
  assign _T_1024 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10395.4]
  assign _T_1027 = _T_1024 & _T_474; // @[MemPrimitives.scala 110:228:@10397.4]
  assign _T_1030 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10399.4]
  assign _T_1033 = _T_1030 & _T_480; // @[MemPrimitives.scala 110:228:@10401.4]
  assign _T_1036 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10403.4]
  assign _T_1039 = _T_1036 & _T_486; // @[MemPrimitives.scala 110:228:@10405.4]
  assign _T_1042 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10407.4]
  assign _T_1045 = _T_1042 & _T_492; // @[MemPrimitives.scala 110:228:@10409.4]
  assign _T_1048 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10411.4]
  assign _T_1051 = _T_1048 & _T_498; // @[MemPrimitives.scala 110:228:@10413.4]
  assign _T_1053 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@10427.4]
  assign _T_1054 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@10428.4]
  assign _T_1055 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@10429.4]
  assign _T_1056 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@10430.4]
  assign _T_1057 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@10431.4]
  assign _T_1058 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@10432.4]
  assign _T_1059 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@10433.4]
  assign _T_1060 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@10434.4]
  assign _T_1061 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 123:41:@10435.4]
  assign _T_1063 = {_T_1053,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10437.4]
  assign _T_1065 = {_T_1054,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10439.4]
  assign _T_1067 = {_T_1055,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10441.4]
  assign _T_1069 = {_T_1056,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10443.4]
  assign _T_1071 = {_T_1057,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10445.4]
  assign _T_1073 = {_T_1058,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10447.4]
  assign _T_1075 = {_T_1059,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10449.4]
  assign _T_1077 = {_T_1060,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10451.4]
  assign _T_1079 = {_T_1061,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10453.4]
  assign _T_1080 = _T_1060 ? _T_1077 : _T_1079; // @[Mux.scala 31:69:@10454.4]
  assign _T_1081 = _T_1059 ? _T_1075 : _T_1080; // @[Mux.scala 31:69:@10455.4]
  assign _T_1082 = _T_1058 ? _T_1073 : _T_1081; // @[Mux.scala 31:69:@10456.4]
  assign _T_1083 = _T_1057 ? _T_1071 : _T_1082; // @[Mux.scala 31:69:@10457.4]
  assign _T_1084 = _T_1056 ? _T_1069 : _T_1083; // @[Mux.scala 31:69:@10458.4]
  assign _T_1085 = _T_1055 ? _T_1067 : _T_1084; // @[Mux.scala 31:69:@10459.4]
  assign _T_1086 = _T_1054 ? _T_1065 : _T_1085; // @[Mux.scala 31:69:@10460.4]
  assign _T_1087 = _T_1053 ? _T_1063 : _T_1086; // @[Mux.scala 31:69:@10461.4]
  assign _T_1095 = _T_1000 & _T_542; // @[MemPrimitives.scala 110:228:@10470.4]
  assign _T_1101 = _T_1006 & _T_548; // @[MemPrimitives.scala 110:228:@10474.4]
  assign _T_1107 = _T_1012 & _T_554; // @[MemPrimitives.scala 110:228:@10478.4]
  assign _T_1113 = _T_1018 & _T_560; // @[MemPrimitives.scala 110:228:@10482.4]
  assign _T_1119 = _T_1024 & _T_566; // @[MemPrimitives.scala 110:228:@10486.4]
  assign _T_1125 = _T_1030 & _T_572; // @[MemPrimitives.scala 110:228:@10490.4]
  assign _T_1131 = _T_1036 & _T_578; // @[MemPrimitives.scala 110:228:@10494.4]
  assign _T_1137 = _T_1042 & _T_584; // @[MemPrimitives.scala 110:228:@10498.4]
  assign _T_1143 = _T_1048 & _T_590; // @[MemPrimitives.scala 110:228:@10502.4]
  assign _T_1145 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@10516.4]
  assign _T_1146 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@10517.4]
  assign _T_1147 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@10518.4]
  assign _T_1148 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@10519.4]
  assign _T_1149 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@10520.4]
  assign _T_1150 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@10521.4]
  assign _T_1151 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@10522.4]
  assign _T_1152 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@10523.4]
  assign _T_1153 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 123:41:@10524.4]
  assign _T_1155 = {_T_1145,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10526.4]
  assign _T_1157 = {_T_1146,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10528.4]
  assign _T_1159 = {_T_1147,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10530.4]
  assign _T_1161 = {_T_1148,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10532.4]
  assign _T_1163 = {_T_1149,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10534.4]
  assign _T_1165 = {_T_1150,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10536.4]
  assign _T_1167 = {_T_1151,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10538.4]
  assign _T_1169 = {_T_1152,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10540.4]
  assign _T_1171 = {_T_1153,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10542.4]
  assign _T_1172 = _T_1152 ? _T_1169 : _T_1171; // @[Mux.scala 31:69:@10543.4]
  assign _T_1173 = _T_1151 ? _T_1167 : _T_1172; // @[Mux.scala 31:69:@10544.4]
  assign _T_1174 = _T_1150 ? _T_1165 : _T_1173; // @[Mux.scala 31:69:@10545.4]
  assign _T_1175 = _T_1149 ? _T_1163 : _T_1174; // @[Mux.scala 31:69:@10546.4]
  assign _T_1176 = _T_1148 ? _T_1161 : _T_1175; // @[Mux.scala 31:69:@10547.4]
  assign _T_1177 = _T_1147 ? _T_1159 : _T_1176; // @[Mux.scala 31:69:@10548.4]
  assign _T_1178 = _T_1146 ? _T_1157 : _T_1177; // @[Mux.scala 31:69:@10549.4]
  assign _T_1179 = _T_1145 ? _T_1155 : _T_1178; // @[Mux.scala 31:69:@10550.4]
  assign _T_1187 = _T_1000 & _T_634; // @[MemPrimitives.scala 110:228:@10559.4]
  assign _T_1193 = _T_1006 & _T_640; // @[MemPrimitives.scala 110:228:@10563.4]
  assign _T_1199 = _T_1012 & _T_646; // @[MemPrimitives.scala 110:228:@10567.4]
  assign _T_1205 = _T_1018 & _T_652; // @[MemPrimitives.scala 110:228:@10571.4]
  assign _T_1211 = _T_1024 & _T_658; // @[MemPrimitives.scala 110:228:@10575.4]
  assign _T_1217 = _T_1030 & _T_664; // @[MemPrimitives.scala 110:228:@10579.4]
  assign _T_1223 = _T_1036 & _T_670; // @[MemPrimitives.scala 110:228:@10583.4]
  assign _T_1229 = _T_1042 & _T_676; // @[MemPrimitives.scala 110:228:@10587.4]
  assign _T_1235 = _T_1048 & _T_682; // @[MemPrimitives.scala 110:228:@10591.4]
  assign _T_1237 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@10605.4]
  assign _T_1238 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@10606.4]
  assign _T_1239 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@10607.4]
  assign _T_1240 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@10608.4]
  assign _T_1241 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@10609.4]
  assign _T_1242 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@10610.4]
  assign _T_1243 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 123:41:@10611.4]
  assign _T_1244 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 123:41:@10612.4]
  assign _T_1245 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 123:41:@10613.4]
  assign _T_1247 = {_T_1237,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10615.4]
  assign _T_1249 = {_T_1238,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10617.4]
  assign _T_1251 = {_T_1239,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10619.4]
  assign _T_1253 = {_T_1240,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10621.4]
  assign _T_1255 = {_T_1241,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10623.4]
  assign _T_1257 = {_T_1242,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10625.4]
  assign _T_1259 = {_T_1243,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10627.4]
  assign _T_1261 = {_T_1244,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10629.4]
  assign _T_1263 = {_T_1245,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10631.4]
  assign _T_1264 = _T_1244 ? _T_1261 : _T_1263; // @[Mux.scala 31:69:@10632.4]
  assign _T_1265 = _T_1243 ? _T_1259 : _T_1264; // @[Mux.scala 31:69:@10633.4]
  assign _T_1266 = _T_1242 ? _T_1257 : _T_1265; // @[Mux.scala 31:69:@10634.4]
  assign _T_1267 = _T_1241 ? _T_1255 : _T_1266; // @[Mux.scala 31:69:@10635.4]
  assign _T_1268 = _T_1240 ? _T_1253 : _T_1267; // @[Mux.scala 31:69:@10636.4]
  assign _T_1269 = _T_1239 ? _T_1251 : _T_1268; // @[Mux.scala 31:69:@10637.4]
  assign _T_1270 = _T_1238 ? _T_1249 : _T_1269; // @[Mux.scala 31:69:@10638.4]
  assign _T_1271 = _T_1237 ? _T_1247 : _T_1270; // @[Mux.scala 31:69:@10639.4]
  assign _T_1276 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10646.4]
  assign _T_1279 = _T_1276 & _T_450; // @[MemPrimitives.scala 110:228:@10648.4]
  assign _T_1282 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10650.4]
  assign _T_1285 = _T_1282 & _T_456; // @[MemPrimitives.scala 110:228:@10652.4]
  assign _T_1288 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10654.4]
  assign _T_1291 = _T_1288 & _T_462; // @[MemPrimitives.scala 110:228:@10656.4]
  assign _T_1294 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10658.4]
  assign _T_1297 = _T_1294 & _T_468; // @[MemPrimitives.scala 110:228:@10660.4]
  assign _T_1300 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10662.4]
  assign _T_1303 = _T_1300 & _T_474; // @[MemPrimitives.scala 110:228:@10664.4]
  assign _T_1306 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10666.4]
  assign _T_1309 = _T_1306 & _T_480; // @[MemPrimitives.scala 110:228:@10668.4]
  assign _T_1312 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10670.4]
  assign _T_1315 = _T_1312 & _T_486; // @[MemPrimitives.scala 110:228:@10672.4]
  assign _T_1318 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10674.4]
  assign _T_1321 = _T_1318 & _T_492; // @[MemPrimitives.scala 110:228:@10676.4]
  assign _T_1324 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10678.4]
  assign _T_1327 = _T_1324 & _T_498; // @[MemPrimitives.scala 110:228:@10680.4]
  assign _T_1329 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@10694.4]
  assign _T_1330 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@10695.4]
  assign _T_1331 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@10696.4]
  assign _T_1332 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@10697.4]
  assign _T_1333 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@10698.4]
  assign _T_1334 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@10699.4]
  assign _T_1335 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 123:41:@10700.4]
  assign _T_1336 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 123:41:@10701.4]
  assign _T_1337 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 123:41:@10702.4]
  assign _T_1339 = {_T_1329,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10704.4]
  assign _T_1341 = {_T_1330,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10706.4]
  assign _T_1343 = {_T_1331,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10708.4]
  assign _T_1345 = {_T_1332,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10710.4]
  assign _T_1347 = {_T_1333,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10712.4]
  assign _T_1349 = {_T_1334,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10714.4]
  assign _T_1351 = {_T_1335,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10716.4]
  assign _T_1353 = {_T_1336,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10718.4]
  assign _T_1355 = {_T_1337,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10720.4]
  assign _T_1356 = _T_1336 ? _T_1353 : _T_1355; // @[Mux.scala 31:69:@10721.4]
  assign _T_1357 = _T_1335 ? _T_1351 : _T_1356; // @[Mux.scala 31:69:@10722.4]
  assign _T_1358 = _T_1334 ? _T_1349 : _T_1357; // @[Mux.scala 31:69:@10723.4]
  assign _T_1359 = _T_1333 ? _T_1347 : _T_1358; // @[Mux.scala 31:69:@10724.4]
  assign _T_1360 = _T_1332 ? _T_1345 : _T_1359; // @[Mux.scala 31:69:@10725.4]
  assign _T_1361 = _T_1331 ? _T_1343 : _T_1360; // @[Mux.scala 31:69:@10726.4]
  assign _T_1362 = _T_1330 ? _T_1341 : _T_1361; // @[Mux.scala 31:69:@10727.4]
  assign _T_1363 = _T_1329 ? _T_1339 : _T_1362; // @[Mux.scala 31:69:@10728.4]
  assign _T_1371 = _T_1276 & _T_542; // @[MemPrimitives.scala 110:228:@10737.4]
  assign _T_1377 = _T_1282 & _T_548; // @[MemPrimitives.scala 110:228:@10741.4]
  assign _T_1383 = _T_1288 & _T_554; // @[MemPrimitives.scala 110:228:@10745.4]
  assign _T_1389 = _T_1294 & _T_560; // @[MemPrimitives.scala 110:228:@10749.4]
  assign _T_1395 = _T_1300 & _T_566; // @[MemPrimitives.scala 110:228:@10753.4]
  assign _T_1401 = _T_1306 & _T_572; // @[MemPrimitives.scala 110:228:@10757.4]
  assign _T_1407 = _T_1312 & _T_578; // @[MemPrimitives.scala 110:228:@10761.4]
  assign _T_1413 = _T_1318 & _T_584; // @[MemPrimitives.scala 110:228:@10765.4]
  assign _T_1419 = _T_1324 & _T_590; // @[MemPrimitives.scala 110:228:@10769.4]
  assign _T_1421 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@10783.4]
  assign _T_1422 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@10784.4]
  assign _T_1423 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@10785.4]
  assign _T_1424 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@10786.4]
  assign _T_1425 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@10787.4]
  assign _T_1426 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@10788.4]
  assign _T_1427 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@10789.4]
  assign _T_1428 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@10790.4]
  assign _T_1429 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 123:41:@10791.4]
  assign _T_1431 = {_T_1421,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10793.4]
  assign _T_1433 = {_T_1422,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10795.4]
  assign _T_1435 = {_T_1423,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10797.4]
  assign _T_1437 = {_T_1424,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10799.4]
  assign _T_1439 = {_T_1425,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10801.4]
  assign _T_1441 = {_T_1426,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10803.4]
  assign _T_1443 = {_T_1427,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10805.4]
  assign _T_1445 = {_T_1428,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10807.4]
  assign _T_1447 = {_T_1429,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10809.4]
  assign _T_1448 = _T_1428 ? _T_1445 : _T_1447; // @[Mux.scala 31:69:@10810.4]
  assign _T_1449 = _T_1427 ? _T_1443 : _T_1448; // @[Mux.scala 31:69:@10811.4]
  assign _T_1450 = _T_1426 ? _T_1441 : _T_1449; // @[Mux.scala 31:69:@10812.4]
  assign _T_1451 = _T_1425 ? _T_1439 : _T_1450; // @[Mux.scala 31:69:@10813.4]
  assign _T_1452 = _T_1424 ? _T_1437 : _T_1451; // @[Mux.scala 31:69:@10814.4]
  assign _T_1453 = _T_1423 ? _T_1435 : _T_1452; // @[Mux.scala 31:69:@10815.4]
  assign _T_1454 = _T_1422 ? _T_1433 : _T_1453; // @[Mux.scala 31:69:@10816.4]
  assign _T_1455 = _T_1421 ? _T_1431 : _T_1454; // @[Mux.scala 31:69:@10817.4]
  assign _T_1463 = _T_1276 & _T_634; // @[MemPrimitives.scala 110:228:@10826.4]
  assign _T_1469 = _T_1282 & _T_640; // @[MemPrimitives.scala 110:228:@10830.4]
  assign _T_1475 = _T_1288 & _T_646; // @[MemPrimitives.scala 110:228:@10834.4]
  assign _T_1481 = _T_1294 & _T_652; // @[MemPrimitives.scala 110:228:@10838.4]
  assign _T_1487 = _T_1300 & _T_658; // @[MemPrimitives.scala 110:228:@10842.4]
  assign _T_1493 = _T_1306 & _T_664; // @[MemPrimitives.scala 110:228:@10846.4]
  assign _T_1499 = _T_1312 & _T_670; // @[MemPrimitives.scala 110:228:@10850.4]
  assign _T_1505 = _T_1318 & _T_676; // @[MemPrimitives.scala 110:228:@10854.4]
  assign _T_1511 = _T_1324 & _T_682; // @[MemPrimitives.scala 110:228:@10858.4]
  assign _T_1513 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@10872.4]
  assign _T_1514 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@10873.4]
  assign _T_1515 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@10874.4]
  assign _T_1516 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@10875.4]
  assign _T_1517 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@10876.4]
  assign _T_1518 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@10877.4]
  assign _T_1519 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@10878.4]
  assign _T_1520 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@10879.4]
  assign _T_1521 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 123:41:@10880.4]
  assign _T_1523 = {_T_1513,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10882.4]
  assign _T_1525 = {_T_1514,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10884.4]
  assign _T_1527 = {_T_1515,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10886.4]
  assign _T_1529 = {_T_1516,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10888.4]
  assign _T_1531 = {_T_1517,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10890.4]
  assign _T_1533 = {_T_1518,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10892.4]
  assign _T_1535 = {_T_1519,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10894.4]
  assign _T_1537 = {_T_1520,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10896.4]
  assign _T_1539 = {_T_1521,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10898.4]
  assign _T_1540 = _T_1520 ? _T_1537 : _T_1539; // @[Mux.scala 31:69:@10899.4]
  assign _T_1541 = _T_1519 ? _T_1535 : _T_1540; // @[Mux.scala 31:69:@10900.4]
  assign _T_1542 = _T_1518 ? _T_1533 : _T_1541; // @[Mux.scala 31:69:@10901.4]
  assign _T_1543 = _T_1517 ? _T_1531 : _T_1542; // @[Mux.scala 31:69:@10902.4]
  assign _T_1544 = _T_1516 ? _T_1529 : _T_1543; // @[Mux.scala 31:69:@10903.4]
  assign _T_1545 = _T_1515 ? _T_1527 : _T_1544; // @[Mux.scala 31:69:@10904.4]
  assign _T_1546 = _T_1514 ? _T_1525 : _T_1545; // @[Mux.scala 31:69:@10905.4]
  assign _T_1547 = _T_1513 ? _T_1523 : _T_1546; // @[Mux.scala 31:69:@10906.4]
  assign _T_1643 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@11035.4 package.scala 96:25:@11036.4]
  assign _T_1647 = _T_1643 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@11045.4]
  assign _T_1640 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@11027.4 package.scala 96:25:@11028.4]
  assign _T_1648 = _T_1640 ? Mem1D_9_io_output : _T_1647; // @[Mux.scala 31:69:@11046.4]
  assign _T_1637 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@11019.4 package.scala 96:25:@11020.4]
  assign _T_1649 = _T_1637 ? Mem1D_8_io_output : _T_1648; // @[Mux.scala 31:69:@11047.4]
  assign _T_1634 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@11011.4 package.scala 96:25:@11012.4]
  assign _T_1650 = _T_1634 ? Mem1D_7_io_output : _T_1649; // @[Mux.scala 31:69:@11048.4]
  assign _T_1631 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@11003.4 package.scala 96:25:@11004.4]
  assign _T_1651 = _T_1631 ? Mem1D_6_io_output : _T_1650; // @[Mux.scala 31:69:@11049.4]
  assign _T_1628 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10995.4 package.scala 96:25:@10996.4]
  assign _T_1652 = _T_1628 ? Mem1D_5_io_output : _T_1651; // @[Mux.scala 31:69:@11050.4]
  assign _T_1625 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10987.4 package.scala 96:25:@10988.4]
  assign _T_1653 = _T_1625 ? Mem1D_4_io_output : _T_1652; // @[Mux.scala 31:69:@11051.4]
  assign _T_1622 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@10979.4 package.scala 96:25:@10980.4]
  assign _T_1654 = _T_1622 ? Mem1D_3_io_output : _T_1653; // @[Mux.scala 31:69:@11052.4]
  assign _T_1619 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@10971.4 package.scala 96:25:@10972.4]
  assign _T_1655 = _T_1619 ? Mem1D_2_io_output : _T_1654; // @[Mux.scala 31:69:@11053.4]
  assign _T_1616 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@10963.4 package.scala 96:25:@10964.4]
  assign _T_1656 = _T_1616 ? Mem1D_1_io_output : _T_1655; // @[Mux.scala 31:69:@11054.4]
  assign _T_1613 = RetimeWrapper_io_out; // @[package.scala 96:25:@10955.4 package.scala 96:25:@10956.4]
  assign _T_1750 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@11179.4 package.scala 96:25:@11180.4]
  assign _T_1754 = _T_1750 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@11189.4]
  assign _T_1747 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@11171.4 package.scala 96:25:@11172.4]
  assign _T_1755 = _T_1747 ? Mem1D_9_io_output : _T_1754; // @[Mux.scala 31:69:@11190.4]
  assign _T_1744 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@11163.4 package.scala 96:25:@11164.4]
  assign _T_1756 = _T_1744 ? Mem1D_8_io_output : _T_1755; // @[Mux.scala 31:69:@11191.4]
  assign _T_1741 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@11155.4 package.scala 96:25:@11156.4]
  assign _T_1757 = _T_1741 ? Mem1D_7_io_output : _T_1756; // @[Mux.scala 31:69:@11192.4]
  assign _T_1738 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@11147.4 package.scala 96:25:@11148.4]
  assign _T_1758 = _T_1738 ? Mem1D_6_io_output : _T_1757; // @[Mux.scala 31:69:@11193.4]
  assign _T_1735 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@11139.4 package.scala 96:25:@11140.4]
  assign _T_1759 = _T_1735 ? Mem1D_5_io_output : _T_1758; // @[Mux.scala 31:69:@11194.4]
  assign _T_1732 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@11131.4 package.scala 96:25:@11132.4]
  assign _T_1760 = _T_1732 ? Mem1D_4_io_output : _T_1759; // @[Mux.scala 31:69:@11195.4]
  assign _T_1729 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@11123.4 package.scala 96:25:@11124.4]
  assign _T_1761 = _T_1729 ? Mem1D_3_io_output : _T_1760; // @[Mux.scala 31:69:@11196.4]
  assign _T_1726 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@11115.4 package.scala 96:25:@11116.4]
  assign _T_1762 = _T_1726 ? Mem1D_2_io_output : _T_1761; // @[Mux.scala 31:69:@11197.4]
  assign _T_1723 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@11107.4 package.scala 96:25:@11108.4]
  assign _T_1763 = _T_1723 ? Mem1D_1_io_output : _T_1762; // @[Mux.scala 31:69:@11198.4]
  assign _T_1720 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@11099.4 package.scala 96:25:@11100.4]
  assign _T_1857 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@11323.4 package.scala 96:25:@11324.4]
  assign _T_1861 = _T_1857 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@11333.4]
  assign _T_1854 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@11315.4 package.scala 96:25:@11316.4]
  assign _T_1862 = _T_1854 ? Mem1D_9_io_output : _T_1861; // @[Mux.scala 31:69:@11334.4]
  assign _T_1851 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@11307.4 package.scala 96:25:@11308.4]
  assign _T_1863 = _T_1851 ? Mem1D_8_io_output : _T_1862; // @[Mux.scala 31:69:@11335.4]
  assign _T_1848 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@11299.4 package.scala 96:25:@11300.4]
  assign _T_1864 = _T_1848 ? Mem1D_7_io_output : _T_1863; // @[Mux.scala 31:69:@11336.4]
  assign _T_1845 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@11291.4 package.scala 96:25:@11292.4]
  assign _T_1865 = _T_1845 ? Mem1D_6_io_output : _T_1864; // @[Mux.scala 31:69:@11337.4]
  assign _T_1842 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@11283.4 package.scala 96:25:@11284.4]
  assign _T_1866 = _T_1842 ? Mem1D_5_io_output : _T_1865; // @[Mux.scala 31:69:@11338.4]
  assign _T_1839 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@11275.4 package.scala 96:25:@11276.4]
  assign _T_1867 = _T_1839 ? Mem1D_4_io_output : _T_1866; // @[Mux.scala 31:69:@11339.4]
  assign _T_1836 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@11267.4 package.scala 96:25:@11268.4]
  assign _T_1868 = _T_1836 ? Mem1D_3_io_output : _T_1867; // @[Mux.scala 31:69:@11340.4]
  assign _T_1833 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@11259.4 package.scala 96:25:@11260.4]
  assign _T_1869 = _T_1833 ? Mem1D_2_io_output : _T_1868; // @[Mux.scala 31:69:@11341.4]
  assign _T_1830 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@11251.4 package.scala 96:25:@11252.4]
  assign _T_1870 = _T_1830 ? Mem1D_1_io_output : _T_1869; // @[Mux.scala 31:69:@11342.4]
  assign _T_1827 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@11243.4 package.scala 96:25:@11244.4]
  assign _T_1964 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@11467.4 package.scala 96:25:@11468.4]
  assign _T_1968 = _T_1964 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@11477.4]
  assign _T_1961 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@11459.4 package.scala 96:25:@11460.4]
  assign _T_1969 = _T_1961 ? Mem1D_9_io_output : _T_1968; // @[Mux.scala 31:69:@11478.4]
  assign _T_1958 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@11451.4 package.scala 96:25:@11452.4]
  assign _T_1970 = _T_1958 ? Mem1D_8_io_output : _T_1969; // @[Mux.scala 31:69:@11479.4]
  assign _T_1955 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@11443.4 package.scala 96:25:@11444.4]
  assign _T_1971 = _T_1955 ? Mem1D_7_io_output : _T_1970; // @[Mux.scala 31:69:@11480.4]
  assign _T_1952 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@11435.4 package.scala 96:25:@11436.4]
  assign _T_1972 = _T_1952 ? Mem1D_6_io_output : _T_1971; // @[Mux.scala 31:69:@11481.4]
  assign _T_1949 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@11427.4 package.scala 96:25:@11428.4]
  assign _T_1973 = _T_1949 ? Mem1D_5_io_output : _T_1972; // @[Mux.scala 31:69:@11482.4]
  assign _T_1946 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@11419.4 package.scala 96:25:@11420.4]
  assign _T_1974 = _T_1946 ? Mem1D_4_io_output : _T_1973; // @[Mux.scala 31:69:@11483.4]
  assign _T_1943 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@11411.4 package.scala 96:25:@11412.4]
  assign _T_1975 = _T_1943 ? Mem1D_3_io_output : _T_1974; // @[Mux.scala 31:69:@11484.4]
  assign _T_1940 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@11403.4 package.scala 96:25:@11404.4]
  assign _T_1976 = _T_1940 ? Mem1D_2_io_output : _T_1975; // @[Mux.scala 31:69:@11485.4]
  assign _T_1937 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@11395.4 package.scala 96:25:@11396.4]
  assign _T_1977 = _T_1937 ? Mem1D_1_io_output : _T_1976; // @[Mux.scala 31:69:@11486.4]
  assign _T_1934 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@11387.4 package.scala 96:25:@11388.4]
  assign _T_2071 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@11611.4 package.scala 96:25:@11612.4]
  assign _T_2075 = _T_2071 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@11621.4]
  assign _T_2068 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@11603.4 package.scala 96:25:@11604.4]
  assign _T_2076 = _T_2068 ? Mem1D_9_io_output : _T_2075; // @[Mux.scala 31:69:@11622.4]
  assign _T_2065 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@11595.4 package.scala 96:25:@11596.4]
  assign _T_2077 = _T_2065 ? Mem1D_8_io_output : _T_2076; // @[Mux.scala 31:69:@11623.4]
  assign _T_2062 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@11587.4 package.scala 96:25:@11588.4]
  assign _T_2078 = _T_2062 ? Mem1D_7_io_output : _T_2077; // @[Mux.scala 31:69:@11624.4]
  assign _T_2059 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@11579.4 package.scala 96:25:@11580.4]
  assign _T_2079 = _T_2059 ? Mem1D_6_io_output : _T_2078; // @[Mux.scala 31:69:@11625.4]
  assign _T_2056 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@11571.4 package.scala 96:25:@11572.4]
  assign _T_2080 = _T_2056 ? Mem1D_5_io_output : _T_2079; // @[Mux.scala 31:69:@11626.4]
  assign _T_2053 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@11563.4 package.scala 96:25:@11564.4]
  assign _T_2081 = _T_2053 ? Mem1D_4_io_output : _T_2080; // @[Mux.scala 31:69:@11627.4]
  assign _T_2050 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@11555.4 package.scala 96:25:@11556.4]
  assign _T_2082 = _T_2050 ? Mem1D_3_io_output : _T_2081; // @[Mux.scala 31:69:@11628.4]
  assign _T_2047 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@11547.4 package.scala 96:25:@11548.4]
  assign _T_2083 = _T_2047 ? Mem1D_2_io_output : _T_2082; // @[Mux.scala 31:69:@11629.4]
  assign _T_2044 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@11539.4 package.scala 96:25:@11540.4]
  assign _T_2084 = _T_2044 ? Mem1D_1_io_output : _T_2083; // @[Mux.scala 31:69:@11630.4]
  assign _T_2041 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@11531.4 package.scala 96:25:@11532.4]
  assign _T_2178 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@11755.4 package.scala 96:25:@11756.4]
  assign _T_2182 = _T_2178 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@11765.4]
  assign _T_2175 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@11747.4 package.scala 96:25:@11748.4]
  assign _T_2183 = _T_2175 ? Mem1D_9_io_output : _T_2182; // @[Mux.scala 31:69:@11766.4]
  assign _T_2172 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@11739.4 package.scala 96:25:@11740.4]
  assign _T_2184 = _T_2172 ? Mem1D_8_io_output : _T_2183; // @[Mux.scala 31:69:@11767.4]
  assign _T_2169 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@11731.4 package.scala 96:25:@11732.4]
  assign _T_2185 = _T_2169 ? Mem1D_7_io_output : _T_2184; // @[Mux.scala 31:69:@11768.4]
  assign _T_2166 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@11723.4 package.scala 96:25:@11724.4]
  assign _T_2186 = _T_2166 ? Mem1D_6_io_output : _T_2185; // @[Mux.scala 31:69:@11769.4]
  assign _T_2163 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@11715.4 package.scala 96:25:@11716.4]
  assign _T_2187 = _T_2163 ? Mem1D_5_io_output : _T_2186; // @[Mux.scala 31:69:@11770.4]
  assign _T_2160 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@11707.4 package.scala 96:25:@11708.4]
  assign _T_2188 = _T_2160 ? Mem1D_4_io_output : _T_2187; // @[Mux.scala 31:69:@11771.4]
  assign _T_2157 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@11699.4 package.scala 96:25:@11700.4]
  assign _T_2189 = _T_2157 ? Mem1D_3_io_output : _T_2188; // @[Mux.scala 31:69:@11772.4]
  assign _T_2154 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@11691.4 package.scala 96:25:@11692.4]
  assign _T_2190 = _T_2154 ? Mem1D_2_io_output : _T_2189; // @[Mux.scala 31:69:@11773.4]
  assign _T_2151 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@11683.4 package.scala 96:25:@11684.4]
  assign _T_2191 = _T_2151 ? Mem1D_1_io_output : _T_2190; // @[Mux.scala 31:69:@11774.4]
  assign _T_2148 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@11675.4 package.scala 96:25:@11676.4]
  assign _T_2285 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@11899.4 package.scala 96:25:@11900.4]
  assign _T_2289 = _T_2285 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@11909.4]
  assign _T_2282 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@11891.4 package.scala 96:25:@11892.4]
  assign _T_2290 = _T_2282 ? Mem1D_9_io_output : _T_2289; // @[Mux.scala 31:69:@11910.4]
  assign _T_2279 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@11883.4 package.scala 96:25:@11884.4]
  assign _T_2291 = _T_2279 ? Mem1D_8_io_output : _T_2290; // @[Mux.scala 31:69:@11911.4]
  assign _T_2276 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@11875.4 package.scala 96:25:@11876.4]
  assign _T_2292 = _T_2276 ? Mem1D_7_io_output : _T_2291; // @[Mux.scala 31:69:@11912.4]
  assign _T_2273 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@11867.4 package.scala 96:25:@11868.4]
  assign _T_2293 = _T_2273 ? Mem1D_6_io_output : _T_2292; // @[Mux.scala 31:69:@11913.4]
  assign _T_2270 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@11859.4 package.scala 96:25:@11860.4]
  assign _T_2294 = _T_2270 ? Mem1D_5_io_output : _T_2293; // @[Mux.scala 31:69:@11914.4]
  assign _T_2267 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@11851.4 package.scala 96:25:@11852.4]
  assign _T_2295 = _T_2267 ? Mem1D_4_io_output : _T_2294; // @[Mux.scala 31:69:@11915.4]
  assign _T_2264 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@11843.4 package.scala 96:25:@11844.4]
  assign _T_2296 = _T_2264 ? Mem1D_3_io_output : _T_2295; // @[Mux.scala 31:69:@11916.4]
  assign _T_2261 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@11835.4 package.scala 96:25:@11836.4]
  assign _T_2297 = _T_2261 ? Mem1D_2_io_output : _T_2296; // @[Mux.scala 31:69:@11917.4]
  assign _T_2258 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@11827.4 package.scala 96:25:@11828.4]
  assign _T_2298 = _T_2258 ? Mem1D_1_io_output : _T_2297; // @[Mux.scala 31:69:@11918.4]
  assign _T_2255 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@11819.4 package.scala 96:25:@11820.4]
  assign _T_2392 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@12043.4 package.scala 96:25:@12044.4]
  assign _T_2396 = _T_2392 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@12053.4]
  assign _T_2389 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@12035.4 package.scala 96:25:@12036.4]
  assign _T_2397 = _T_2389 ? Mem1D_9_io_output : _T_2396; // @[Mux.scala 31:69:@12054.4]
  assign _T_2386 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@12027.4 package.scala 96:25:@12028.4]
  assign _T_2398 = _T_2386 ? Mem1D_8_io_output : _T_2397; // @[Mux.scala 31:69:@12055.4]
  assign _T_2383 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@12019.4 package.scala 96:25:@12020.4]
  assign _T_2399 = _T_2383 ? Mem1D_7_io_output : _T_2398; // @[Mux.scala 31:69:@12056.4]
  assign _T_2380 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@12011.4 package.scala 96:25:@12012.4]
  assign _T_2400 = _T_2380 ? Mem1D_6_io_output : _T_2399; // @[Mux.scala 31:69:@12057.4]
  assign _T_2377 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@12003.4 package.scala 96:25:@12004.4]
  assign _T_2401 = _T_2377 ? Mem1D_5_io_output : _T_2400; // @[Mux.scala 31:69:@12058.4]
  assign _T_2374 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@11995.4 package.scala 96:25:@11996.4]
  assign _T_2402 = _T_2374 ? Mem1D_4_io_output : _T_2401; // @[Mux.scala 31:69:@12059.4]
  assign _T_2371 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@11987.4 package.scala 96:25:@11988.4]
  assign _T_2403 = _T_2371 ? Mem1D_3_io_output : _T_2402; // @[Mux.scala 31:69:@12060.4]
  assign _T_2368 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@11979.4 package.scala 96:25:@11980.4]
  assign _T_2404 = _T_2368 ? Mem1D_2_io_output : _T_2403; // @[Mux.scala 31:69:@12061.4]
  assign _T_2365 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@11971.4 package.scala 96:25:@11972.4]
  assign _T_2405 = _T_2365 ? Mem1D_1_io_output : _T_2404; // @[Mux.scala 31:69:@12062.4]
  assign _T_2362 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@11963.4 package.scala 96:25:@11964.4]
  assign _T_2499 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@12187.4 package.scala 96:25:@12188.4]
  assign _T_2503 = _T_2499 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@12197.4]
  assign _T_2496 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@12179.4 package.scala 96:25:@12180.4]
  assign _T_2504 = _T_2496 ? Mem1D_9_io_output : _T_2503; // @[Mux.scala 31:69:@12198.4]
  assign _T_2493 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@12171.4 package.scala 96:25:@12172.4]
  assign _T_2505 = _T_2493 ? Mem1D_8_io_output : _T_2504; // @[Mux.scala 31:69:@12199.4]
  assign _T_2490 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@12163.4 package.scala 96:25:@12164.4]
  assign _T_2506 = _T_2490 ? Mem1D_7_io_output : _T_2505; // @[Mux.scala 31:69:@12200.4]
  assign _T_2487 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@12155.4 package.scala 96:25:@12156.4]
  assign _T_2507 = _T_2487 ? Mem1D_6_io_output : _T_2506; // @[Mux.scala 31:69:@12201.4]
  assign _T_2484 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@12147.4 package.scala 96:25:@12148.4]
  assign _T_2508 = _T_2484 ? Mem1D_5_io_output : _T_2507; // @[Mux.scala 31:69:@12202.4]
  assign _T_2481 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@12139.4 package.scala 96:25:@12140.4]
  assign _T_2509 = _T_2481 ? Mem1D_4_io_output : _T_2508; // @[Mux.scala 31:69:@12203.4]
  assign _T_2478 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@12131.4 package.scala 96:25:@12132.4]
  assign _T_2510 = _T_2478 ? Mem1D_3_io_output : _T_2509; // @[Mux.scala 31:69:@12204.4]
  assign _T_2475 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@12123.4 package.scala 96:25:@12124.4]
  assign _T_2511 = _T_2475 ? Mem1D_2_io_output : _T_2510; // @[Mux.scala 31:69:@12205.4]
  assign _T_2472 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@12115.4 package.scala 96:25:@12116.4]
  assign _T_2512 = _T_2472 ? Mem1D_1_io_output : _T_2511; // @[Mux.scala 31:69:@12206.4]
  assign _T_2469 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@12107.4 package.scala 96:25:@12108.4]
  assign io_rPort_8_output_0 = _T_2469 ? Mem1D_io_output : _T_2512; // @[MemPrimitives.scala 148:13:@12208.4]
  assign io_rPort_7_output_0 = _T_2362 ? Mem1D_io_output : _T_2405; // @[MemPrimitives.scala 148:13:@12064.4]
  assign io_rPort_6_output_0 = _T_2255 ? Mem1D_io_output : _T_2298; // @[MemPrimitives.scala 148:13:@11920.4]
  assign io_rPort_5_output_0 = _T_2148 ? Mem1D_io_output : _T_2191; // @[MemPrimitives.scala 148:13:@11776.4]
  assign io_rPort_4_output_0 = _T_2041 ? Mem1D_io_output : _T_2084; // @[MemPrimitives.scala 148:13:@11632.4]
  assign io_rPort_3_output_0 = _T_1934 ? Mem1D_io_output : _T_1977; // @[MemPrimitives.scala 148:13:@11488.4]
  assign io_rPort_2_output_0 = _T_1827 ? Mem1D_io_output : _T_1870; // @[MemPrimitives.scala 148:13:@11344.4]
  assign io_rPort_1_output_0 = _T_1720 ? Mem1D_io_output : _T_1763; // @[MemPrimitives.scala 148:13:@11200.4]
  assign io_rPort_0_output_0 = _T_1613 ? Mem1D_io_output : _T_1656; // @[MemPrimitives.scala 148:13:@11056.4]
  assign Mem1D_clock = clock; // @[:@9510.4]
  assign Mem1D_reset = reset; // @[:@9511.4]
  assign Mem1D_io_r_ofs_0 = _T_535[8:0]; // @[MemPrimitives.scala 127:28:@9931.4]
  assign Mem1D_io_r_backpressure = _T_535[9]; // @[MemPrimitives.scala 128:32:@9932.4]
  assign Mem1D_io_w_ofs_0 = _T_322[8:0]; // @[MemPrimitives.scala 94:28:@9710.4]
  assign Mem1D_io_w_data_0 = _T_322[16:9]; // @[MemPrimitives.scala 95:29:@9711.4]
  assign Mem1D_io_w_en_0 = _T_322[17]; // @[MemPrimitives.scala 96:27:@9712.4]
  assign Mem1D_1_clock = clock; // @[:@9526.4]
  assign Mem1D_1_reset = reset; // @[:@9527.4]
  assign Mem1D_1_io_r_ofs_0 = _T_627[8:0]; // @[MemPrimitives.scala 127:28:@10020.4]
  assign Mem1D_1_io_r_backpressure = _T_627[9]; // @[MemPrimitives.scala 128:32:@10021.4]
  assign Mem1D_1_io_w_ofs_0 = _T_333[8:0]; // @[MemPrimitives.scala 94:28:@9722.4]
  assign Mem1D_1_io_w_data_0 = _T_333[16:9]; // @[MemPrimitives.scala 95:29:@9723.4]
  assign Mem1D_1_io_w_en_0 = _T_333[17]; // @[MemPrimitives.scala 96:27:@9724.4]
  assign Mem1D_2_clock = clock; // @[:@9542.4]
  assign Mem1D_2_reset = reset; // @[:@9543.4]
  assign Mem1D_2_io_r_ofs_0 = _T_719[8:0]; // @[MemPrimitives.scala 127:28:@10109.4]
  assign Mem1D_2_io_r_backpressure = _T_719[9]; // @[MemPrimitives.scala 128:32:@10110.4]
  assign Mem1D_2_io_w_ofs_0 = _T_344[8:0]; // @[MemPrimitives.scala 94:28:@9734.4]
  assign Mem1D_2_io_w_data_0 = _T_344[16:9]; // @[MemPrimitives.scala 95:29:@9735.4]
  assign Mem1D_2_io_w_en_0 = _T_344[17]; // @[MemPrimitives.scala 96:27:@9736.4]
  assign Mem1D_3_clock = clock; // @[:@9558.4]
  assign Mem1D_3_reset = reset; // @[:@9559.4]
  assign Mem1D_3_io_r_ofs_0 = _T_811[8:0]; // @[MemPrimitives.scala 127:28:@10198.4]
  assign Mem1D_3_io_r_backpressure = _T_811[9]; // @[MemPrimitives.scala 128:32:@10199.4]
  assign Mem1D_3_io_w_ofs_0 = _T_355[8:0]; // @[MemPrimitives.scala 94:28:@9746.4]
  assign Mem1D_3_io_w_data_0 = _T_355[16:9]; // @[MemPrimitives.scala 95:29:@9747.4]
  assign Mem1D_3_io_w_en_0 = _T_355[17]; // @[MemPrimitives.scala 96:27:@9748.4]
  assign Mem1D_4_clock = clock; // @[:@9574.4]
  assign Mem1D_4_reset = reset; // @[:@9575.4]
  assign Mem1D_4_io_r_ofs_0 = _T_903[8:0]; // @[MemPrimitives.scala 127:28:@10287.4]
  assign Mem1D_4_io_r_backpressure = _T_903[9]; // @[MemPrimitives.scala 128:32:@10288.4]
  assign Mem1D_4_io_w_ofs_0 = _T_366[8:0]; // @[MemPrimitives.scala 94:28:@9758.4]
  assign Mem1D_4_io_w_data_0 = _T_366[16:9]; // @[MemPrimitives.scala 95:29:@9759.4]
  assign Mem1D_4_io_w_en_0 = _T_366[17]; // @[MemPrimitives.scala 96:27:@9760.4]
  assign Mem1D_5_clock = clock; // @[:@9590.4]
  assign Mem1D_5_reset = reset; // @[:@9591.4]
  assign Mem1D_5_io_r_ofs_0 = _T_995[8:0]; // @[MemPrimitives.scala 127:28:@10376.4]
  assign Mem1D_5_io_r_backpressure = _T_995[9]; // @[MemPrimitives.scala 128:32:@10377.4]
  assign Mem1D_5_io_w_ofs_0 = _T_377[8:0]; // @[MemPrimitives.scala 94:28:@9770.4]
  assign Mem1D_5_io_w_data_0 = _T_377[16:9]; // @[MemPrimitives.scala 95:29:@9771.4]
  assign Mem1D_5_io_w_en_0 = _T_377[17]; // @[MemPrimitives.scala 96:27:@9772.4]
  assign Mem1D_6_clock = clock; // @[:@9606.4]
  assign Mem1D_6_reset = reset; // @[:@9607.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1087[8:0]; // @[MemPrimitives.scala 127:28:@10465.4]
  assign Mem1D_6_io_r_backpressure = _T_1087[9]; // @[MemPrimitives.scala 128:32:@10466.4]
  assign Mem1D_6_io_w_ofs_0 = _T_388[8:0]; // @[MemPrimitives.scala 94:28:@9782.4]
  assign Mem1D_6_io_w_data_0 = _T_388[16:9]; // @[MemPrimitives.scala 95:29:@9783.4]
  assign Mem1D_6_io_w_en_0 = _T_388[17]; // @[MemPrimitives.scala 96:27:@9784.4]
  assign Mem1D_7_clock = clock; // @[:@9622.4]
  assign Mem1D_7_reset = reset; // @[:@9623.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1179[8:0]; // @[MemPrimitives.scala 127:28:@10554.4]
  assign Mem1D_7_io_r_backpressure = _T_1179[9]; // @[MemPrimitives.scala 128:32:@10555.4]
  assign Mem1D_7_io_w_ofs_0 = _T_399[8:0]; // @[MemPrimitives.scala 94:28:@9794.4]
  assign Mem1D_7_io_w_data_0 = _T_399[16:9]; // @[MemPrimitives.scala 95:29:@9795.4]
  assign Mem1D_7_io_w_en_0 = _T_399[17]; // @[MemPrimitives.scala 96:27:@9796.4]
  assign Mem1D_8_clock = clock; // @[:@9638.4]
  assign Mem1D_8_reset = reset; // @[:@9639.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1271[8:0]; // @[MemPrimitives.scala 127:28:@10643.4]
  assign Mem1D_8_io_r_backpressure = _T_1271[9]; // @[MemPrimitives.scala 128:32:@10644.4]
  assign Mem1D_8_io_w_ofs_0 = _T_410[8:0]; // @[MemPrimitives.scala 94:28:@9806.4]
  assign Mem1D_8_io_w_data_0 = _T_410[16:9]; // @[MemPrimitives.scala 95:29:@9807.4]
  assign Mem1D_8_io_w_en_0 = _T_410[17]; // @[MemPrimitives.scala 96:27:@9808.4]
  assign Mem1D_9_clock = clock; // @[:@9654.4]
  assign Mem1D_9_reset = reset; // @[:@9655.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1363[8:0]; // @[MemPrimitives.scala 127:28:@10732.4]
  assign Mem1D_9_io_r_backpressure = _T_1363[9]; // @[MemPrimitives.scala 128:32:@10733.4]
  assign Mem1D_9_io_w_ofs_0 = _T_421[8:0]; // @[MemPrimitives.scala 94:28:@9818.4]
  assign Mem1D_9_io_w_data_0 = _T_421[16:9]; // @[MemPrimitives.scala 95:29:@9819.4]
  assign Mem1D_9_io_w_en_0 = _T_421[17]; // @[MemPrimitives.scala 96:27:@9820.4]
  assign Mem1D_10_clock = clock; // @[:@9670.4]
  assign Mem1D_10_reset = reset; // @[:@9671.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1455[8:0]; // @[MemPrimitives.scala 127:28:@10821.4]
  assign Mem1D_10_io_r_backpressure = _T_1455[9]; // @[MemPrimitives.scala 128:32:@10822.4]
  assign Mem1D_10_io_w_ofs_0 = _T_432[8:0]; // @[MemPrimitives.scala 94:28:@9830.4]
  assign Mem1D_10_io_w_data_0 = _T_432[16:9]; // @[MemPrimitives.scala 95:29:@9831.4]
  assign Mem1D_10_io_w_en_0 = _T_432[17]; // @[MemPrimitives.scala 96:27:@9832.4]
  assign Mem1D_11_clock = clock; // @[:@9686.4]
  assign Mem1D_11_reset = reset; // @[:@9687.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1547[8:0]; // @[MemPrimitives.scala 127:28:@10910.4]
  assign Mem1D_11_io_r_backpressure = _T_1547[9]; // @[MemPrimitives.scala 128:32:@10911.4]
  assign Mem1D_11_io_w_ofs_0 = _T_443[8:0]; // @[MemPrimitives.scala 94:28:@9842.4]
  assign Mem1D_11_io_w_data_0 = _T_443[16:9]; // @[MemPrimitives.scala 95:29:@9843.4]
  assign Mem1D_11_io_w_en_0 = _T_443[17]; // @[MemPrimitives.scala 96:27:@9844.4]
  assign StickySelects_clock = clock; // @[:@9882.4]
  assign StickySelects_reset = reset; // @[:@9883.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_451; // @[MemPrimitives.scala 122:60:@9884.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_457; // @[MemPrimitives.scala 122:60:@9885.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_463; // @[MemPrimitives.scala 122:60:@9886.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_469; // @[MemPrimitives.scala 122:60:@9887.4]
  assign StickySelects_io_ins_4 = io_rPort_4_en_0 & _T_475; // @[MemPrimitives.scala 122:60:@9888.4]
  assign StickySelects_io_ins_5 = io_rPort_5_en_0 & _T_481; // @[MemPrimitives.scala 122:60:@9889.4]
  assign StickySelects_io_ins_6 = io_rPort_6_en_0 & _T_487; // @[MemPrimitives.scala 122:60:@9890.4]
  assign StickySelects_io_ins_7 = io_rPort_7_en_0 & _T_493; // @[MemPrimitives.scala 122:60:@9891.4]
  assign StickySelects_io_ins_8 = io_rPort_8_en_0 & _T_499; // @[MemPrimitives.scala 122:60:@9892.4]
  assign StickySelects_1_clock = clock; // @[:@9971.4]
  assign StickySelects_1_reset = reset; // @[:@9972.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_543; // @[MemPrimitives.scala 122:60:@9973.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_549; // @[MemPrimitives.scala 122:60:@9974.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_555; // @[MemPrimitives.scala 122:60:@9975.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_561; // @[MemPrimitives.scala 122:60:@9976.4]
  assign StickySelects_1_io_ins_4 = io_rPort_4_en_0 & _T_567; // @[MemPrimitives.scala 122:60:@9977.4]
  assign StickySelects_1_io_ins_5 = io_rPort_5_en_0 & _T_573; // @[MemPrimitives.scala 122:60:@9978.4]
  assign StickySelects_1_io_ins_6 = io_rPort_6_en_0 & _T_579; // @[MemPrimitives.scala 122:60:@9979.4]
  assign StickySelects_1_io_ins_7 = io_rPort_7_en_0 & _T_585; // @[MemPrimitives.scala 122:60:@9980.4]
  assign StickySelects_1_io_ins_8 = io_rPort_8_en_0 & _T_591; // @[MemPrimitives.scala 122:60:@9981.4]
  assign StickySelects_2_clock = clock; // @[:@10060.4]
  assign StickySelects_2_reset = reset; // @[:@10061.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@10062.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_641; // @[MemPrimitives.scala 122:60:@10063.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_647; // @[MemPrimitives.scala 122:60:@10064.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_653; // @[MemPrimitives.scala 122:60:@10065.4]
  assign StickySelects_2_io_ins_4 = io_rPort_4_en_0 & _T_659; // @[MemPrimitives.scala 122:60:@10066.4]
  assign StickySelects_2_io_ins_5 = io_rPort_5_en_0 & _T_665; // @[MemPrimitives.scala 122:60:@10067.4]
  assign StickySelects_2_io_ins_6 = io_rPort_6_en_0 & _T_671; // @[MemPrimitives.scala 122:60:@10068.4]
  assign StickySelects_2_io_ins_7 = io_rPort_7_en_0 & _T_677; // @[MemPrimitives.scala 122:60:@10069.4]
  assign StickySelects_2_io_ins_8 = io_rPort_8_en_0 & _T_683; // @[MemPrimitives.scala 122:60:@10070.4]
  assign StickySelects_3_clock = clock; // @[:@10149.4]
  assign StickySelects_3_reset = reset; // @[:@10150.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_727; // @[MemPrimitives.scala 122:60:@10151.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_733; // @[MemPrimitives.scala 122:60:@10152.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_739; // @[MemPrimitives.scala 122:60:@10153.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_745; // @[MemPrimitives.scala 122:60:@10154.4]
  assign StickySelects_3_io_ins_4 = io_rPort_4_en_0 & _T_751; // @[MemPrimitives.scala 122:60:@10155.4]
  assign StickySelects_3_io_ins_5 = io_rPort_5_en_0 & _T_757; // @[MemPrimitives.scala 122:60:@10156.4]
  assign StickySelects_3_io_ins_6 = io_rPort_6_en_0 & _T_763; // @[MemPrimitives.scala 122:60:@10157.4]
  assign StickySelects_3_io_ins_7 = io_rPort_7_en_0 & _T_769; // @[MemPrimitives.scala 122:60:@10158.4]
  assign StickySelects_3_io_ins_8 = io_rPort_8_en_0 & _T_775; // @[MemPrimitives.scala 122:60:@10159.4]
  assign StickySelects_4_clock = clock; // @[:@10238.4]
  assign StickySelects_4_reset = reset; // @[:@10239.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_819; // @[MemPrimitives.scala 122:60:@10240.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_825; // @[MemPrimitives.scala 122:60:@10241.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_831; // @[MemPrimitives.scala 122:60:@10242.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_837; // @[MemPrimitives.scala 122:60:@10243.4]
  assign StickySelects_4_io_ins_4 = io_rPort_4_en_0 & _T_843; // @[MemPrimitives.scala 122:60:@10244.4]
  assign StickySelects_4_io_ins_5 = io_rPort_5_en_0 & _T_849; // @[MemPrimitives.scala 122:60:@10245.4]
  assign StickySelects_4_io_ins_6 = io_rPort_6_en_0 & _T_855; // @[MemPrimitives.scala 122:60:@10246.4]
  assign StickySelects_4_io_ins_7 = io_rPort_7_en_0 & _T_861; // @[MemPrimitives.scala 122:60:@10247.4]
  assign StickySelects_4_io_ins_8 = io_rPort_8_en_0 & _T_867; // @[MemPrimitives.scala 122:60:@10248.4]
  assign StickySelects_5_clock = clock; // @[:@10327.4]
  assign StickySelects_5_reset = reset; // @[:@10328.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_911; // @[MemPrimitives.scala 122:60:@10329.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_917; // @[MemPrimitives.scala 122:60:@10330.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_923; // @[MemPrimitives.scala 122:60:@10331.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_929; // @[MemPrimitives.scala 122:60:@10332.4]
  assign StickySelects_5_io_ins_4 = io_rPort_4_en_0 & _T_935; // @[MemPrimitives.scala 122:60:@10333.4]
  assign StickySelects_5_io_ins_5 = io_rPort_5_en_0 & _T_941; // @[MemPrimitives.scala 122:60:@10334.4]
  assign StickySelects_5_io_ins_6 = io_rPort_6_en_0 & _T_947; // @[MemPrimitives.scala 122:60:@10335.4]
  assign StickySelects_5_io_ins_7 = io_rPort_7_en_0 & _T_953; // @[MemPrimitives.scala 122:60:@10336.4]
  assign StickySelects_5_io_ins_8 = io_rPort_8_en_0 & _T_959; // @[MemPrimitives.scala 122:60:@10337.4]
  assign StickySelects_6_clock = clock; // @[:@10416.4]
  assign StickySelects_6_reset = reset; // @[:@10417.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1003; // @[MemPrimitives.scala 122:60:@10418.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1009; // @[MemPrimitives.scala 122:60:@10419.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_1015; // @[MemPrimitives.scala 122:60:@10420.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_1021; // @[MemPrimitives.scala 122:60:@10421.4]
  assign StickySelects_6_io_ins_4 = io_rPort_4_en_0 & _T_1027; // @[MemPrimitives.scala 122:60:@10422.4]
  assign StickySelects_6_io_ins_5 = io_rPort_5_en_0 & _T_1033; // @[MemPrimitives.scala 122:60:@10423.4]
  assign StickySelects_6_io_ins_6 = io_rPort_6_en_0 & _T_1039; // @[MemPrimitives.scala 122:60:@10424.4]
  assign StickySelects_6_io_ins_7 = io_rPort_7_en_0 & _T_1045; // @[MemPrimitives.scala 122:60:@10425.4]
  assign StickySelects_6_io_ins_8 = io_rPort_8_en_0 & _T_1051; // @[MemPrimitives.scala 122:60:@10426.4]
  assign StickySelects_7_clock = clock; // @[:@10505.4]
  assign StickySelects_7_reset = reset; // @[:@10506.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1095; // @[MemPrimitives.scala 122:60:@10507.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1101; // @[MemPrimitives.scala 122:60:@10508.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1107; // @[MemPrimitives.scala 122:60:@10509.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1113; // @[MemPrimitives.scala 122:60:@10510.4]
  assign StickySelects_7_io_ins_4 = io_rPort_4_en_0 & _T_1119; // @[MemPrimitives.scala 122:60:@10511.4]
  assign StickySelects_7_io_ins_5 = io_rPort_5_en_0 & _T_1125; // @[MemPrimitives.scala 122:60:@10512.4]
  assign StickySelects_7_io_ins_6 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 122:60:@10513.4]
  assign StickySelects_7_io_ins_7 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 122:60:@10514.4]
  assign StickySelects_7_io_ins_8 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 122:60:@10515.4]
  assign StickySelects_8_clock = clock; // @[:@10594.4]
  assign StickySelects_8_reset = reset; // @[:@10595.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1187; // @[MemPrimitives.scala 122:60:@10596.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1193; // @[MemPrimitives.scala 122:60:@10597.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_1199; // @[MemPrimitives.scala 122:60:@10598.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@10599.4]
  assign StickySelects_8_io_ins_4 = io_rPort_4_en_0 & _T_1211; // @[MemPrimitives.scala 122:60:@10600.4]
  assign StickySelects_8_io_ins_5 = io_rPort_5_en_0 & _T_1217; // @[MemPrimitives.scala 122:60:@10601.4]
  assign StickySelects_8_io_ins_6 = io_rPort_6_en_0 & _T_1223; // @[MemPrimitives.scala 122:60:@10602.4]
  assign StickySelects_8_io_ins_7 = io_rPort_7_en_0 & _T_1229; // @[MemPrimitives.scala 122:60:@10603.4]
  assign StickySelects_8_io_ins_8 = io_rPort_8_en_0 & _T_1235; // @[MemPrimitives.scala 122:60:@10604.4]
  assign StickySelects_9_clock = clock; // @[:@10683.4]
  assign StickySelects_9_reset = reset; // @[:@10684.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1279; // @[MemPrimitives.scala 122:60:@10685.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1285; // @[MemPrimitives.scala 122:60:@10686.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1291; // @[MemPrimitives.scala 122:60:@10687.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1297; // @[MemPrimitives.scala 122:60:@10688.4]
  assign StickySelects_9_io_ins_4 = io_rPort_4_en_0 & _T_1303; // @[MemPrimitives.scala 122:60:@10689.4]
  assign StickySelects_9_io_ins_5 = io_rPort_5_en_0 & _T_1309; // @[MemPrimitives.scala 122:60:@10690.4]
  assign StickySelects_9_io_ins_6 = io_rPort_6_en_0 & _T_1315; // @[MemPrimitives.scala 122:60:@10691.4]
  assign StickySelects_9_io_ins_7 = io_rPort_7_en_0 & _T_1321; // @[MemPrimitives.scala 122:60:@10692.4]
  assign StickySelects_9_io_ins_8 = io_rPort_8_en_0 & _T_1327; // @[MemPrimitives.scala 122:60:@10693.4]
  assign StickySelects_10_clock = clock; // @[:@10772.4]
  assign StickySelects_10_reset = reset; // @[:@10773.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1371; // @[MemPrimitives.scala 122:60:@10774.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_1377; // @[MemPrimitives.scala 122:60:@10775.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_1383; // @[MemPrimitives.scala 122:60:@10776.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_1389; // @[MemPrimitives.scala 122:60:@10777.4]
  assign StickySelects_10_io_ins_4 = io_rPort_4_en_0 & _T_1395; // @[MemPrimitives.scala 122:60:@10778.4]
  assign StickySelects_10_io_ins_5 = io_rPort_5_en_0 & _T_1401; // @[MemPrimitives.scala 122:60:@10779.4]
  assign StickySelects_10_io_ins_6 = io_rPort_6_en_0 & _T_1407; // @[MemPrimitives.scala 122:60:@10780.4]
  assign StickySelects_10_io_ins_7 = io_rPort_7_en_0 & _T_1413; // @[MemPrimitives.scala 122:60:@10781.4]
  assign StickySelects_10_io_ins_8 = io_rPort_8_en_0 & _T_1419; // @[MemPrimitives.scala 122:60:@10782.4]
  assign StickySelects_11_clock = clock; // @[:@10861.4]
  assign StickySelects_11_reset = reset; // @[:@10862.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1463; // @[MemPrimitives.scala 122:60:@10863.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1469; // @[MemPrimitives.scala 122:60:@10864.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1475; // @[MemPrimitives.scala 122:60:@10865.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1481; // @[MemPrimitives.scala 122:60:@10866.4]
  assign StickySelects_11_io_ins_4 = io_rPort_4_en_0 & _T_1487; // @[MemPrimitives.scala 122:60:@10867.4]
  assign StickySelects_11_io_ins_5 = io_rPort_5_en_0 & _T_1493; // @[MemPrimitives.scala 122:60:@10868.4]
  assign StickySelects_11_io_ins_6 = io_rPort_6_en_0 & _T_1499; // @[MemPrimitives.scala 122:60:@10869.4]
  assign StickySelects_11_io_ins_7 = io_rPort_7_en_0 & _T_1505; // @[MemPrimitives.scala 122:60:@10870.4]
  assign StickySelects_11_io_ins_8 = io_rPort_8_en_0 & _T_1511; // @[MemPrimitives.scala 122:60:@10871.4]
  assign RetimeWrapper_clock = clock; // @[:@10951.4]
  assign RetimeWrapper_reset = reset; // @[:@10952.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10954.4]
  assign RetimeWrapper_io_in = _T_451 & io_rPort_0_en_0; // @[package.scala 94:16:@10953.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10959.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10960.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10962.4]
  assign RetimeWrapper_1_io_in = _T_543 & io_rPort_0_en_0; // @[package.scala 94:16:@10961.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10967.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10968.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10970.4]
  assign RetimeWrapper_2_io_in = _T_635 & io_rPort_0_en_0; // @[package.scala 94:16:@10969.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10975.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10976.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10978.4]
  assign RetimeWrapper_3_io_in = _T_727 & io_rPort_0_en_0; // @[package.scala 94:16:@10977.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10983.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10984.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10986.4]
  assign RetimeWrapper_4_io_in = _T_819 & io_rPort_0_en_0; // @[package.scala 94:16:@10985.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10991.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10992.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10994.4]
  assign RetimeWrapper_5_io_in = _T_911 & io_rPort_0_en_0; // @[package.scala 94:16:@10993.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10999.4]
  assign RetimeWrapper_6_reset = reset; // @[:@11000.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@11002.4]
  assign RetimeWrapper_6_io_in = _T_1003 & io_rPort_0_en_0; // @[package.scala 94:16:@11001.4]
  assign RetimeWrapper_7_clock = clock; // @[:@11007.4]
  assign RetimeWrapper_7_reset = reset; // @[:@11008.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@11010.4]
  assign RetimeWrapper_7_io_in = _T_1095 & io_rPort_0_en_0; // @[package.scala 94:16:@11009.4]
  assign RetimeWrapper_8_clock = clock; // @[:@11015.4]
  assign RetimeWrapper_8_reset = reset; // @[:@11016.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@11018.4]
  assign RetimeWrapper_8_io_in = _T_1187 & io_rPort_0_en_0; // @[package.scala 94:16:@11017.4]
  assign RetimeWrapper_9_clock = clock; // @[:@11023.4]
  assign RetimeWrapper_9_reset = reset; // @[:@11024.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@11026.4]
  assign RetimeWrapper_9_io_in = _T_1279 & io_rPort_0_en_0; // @[package.scala 94:16:@11025.4]
  assign RetimeWrapper_10_clock = clock; // @[:@11031.4]
  assign RetimeWrapper_10_reset = reset; // @[:@11032.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@11034.4]
  assign RetimeWrapper_10_io_in = _T_1371 & io_rPort_0_en_0; // @[package.scala 94:16:@11033.4]
  assign RetimeWrapper_11_clock = clock; // @[:@11039.4]
  assign RetimeWrapper_11_reset = reset; // @[:@11040.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@11042.4]
  assign RetimeWrapper_11_io_in = _T_1463 & io_rPort_0_en_0; // @[package.scala 94:16:@11041.4]
  assign RetimeWrapper_12_clock = clock; // @[:@11095.4]
  assign RetimeWrapper_12_reset = reset; // @[:@11096.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11098.4]
  assign RetimeWrapper_12_io_in = _T_457 & io_rPort_1_en_0; // @[package.scala 94:16:@11097.4]
  assign RetimeWrapper_13_clock = clock; // @[:@11103.4]
  assign RetimeWrapper_13_reset = reset; // @[:@11104.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11106.4]
  assign RetimeWrapper_13_io_in = _T_549 & io_rPort_1_en_0; // @[package.scala 94:16:@11105.4]
  assign RetimeWrapper_14_clock = clock; // @[:@11111.4]
  assign RetimeWrapper_14_reset = reset; // @[:@11112.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11114.4]
  assign RetimeWrapper_14_io_in = _T_641 & io_rPort_1_en_0; // @[package.scala 94:16:@11113.4]
  assign RetimeWrapper_15_clock = clock; // @[:@11119.4]
  assign RetimeWrapper_15_reset = reset; // @[:@11120.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11122.4]
  assign RetimeWrapper_15_io_in = _T_733 & io_rPort_1_en_0; // @[package.scala 94:16:@11121.4]
  assign RetimeWrapper_16_clock = clock; // @[:@11127.4]
  assign RetimeWrapper_16_reset = reset; // @[:@11128.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11130.4]
  assign RetimeWrapper_16_io_in = _T_825 & io_rPort_1_en_0; // @[package.scala 94:16:@11129.4]
  assign RetimeWrapper_17_clock = clock; // @[:@11135.4]
  assign RetimeWrapper_17_reset = reset; // @[:@11136.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11138.4]
  assign RetimeWrapper_17_io_in = _T_917 & io_rPort_1_en_0; // @[package.scala 94:16:@11137.4]
  assign RetimeWrapper_18_clock = clock; // @[:@11143.4]
  assign RetimeWrapper_18_reset = reset; // @[:@11144.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11146.4]
  assign RetimeWrapper_18_io_in = _T_1009 & io_rPort_1_en_0; // @[package.scala 94:16:@11145.4]
  assign RetimeWrapper_19_clock = clock; // @[:@11151.4]
  assign RetimeWrapper_19_reset = reset; // @[:@11152.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11154.4]
  assign RetimeWrapper_19_io_in = _T_1101 & io_rPort_1_en_0; // @[package.scala 94:16:@11153.4]
  assign RetimeWrapper_20_clock = clock; // @[:@11159.4]
  assign RetimeWrapper_20_reset = reset; // @[:@11160.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11162.4]
  assign RetimeWrapper_20_io_in = _T_1193 & io_rPort_1_en_0; // @[package.scala 94:16:@11161.4]
  assign RetimeWrapper_21_clock = clock; // @[:@11167.4]
  assign RetimeWrapper_21_reset = reset; // @[:@11168.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11170.4]
  assign RetimeWrapper_21_io_in = _T_1285 & io_rPort_1_en_0; // @[package.scala 94:16:@11169.4]
  assign RetimeWrapper_22_clock = clock; // @[:@11175.4]
  assign RetimeWrapper_22_reset = reset; // @[:@11176.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11178.4]
  assign RetimeWrapper_22_io_in = _T_1377 & io_rPort_1_en_0; // @[package.scala 94:16:@11177.4]
  assign RetimeWrapper_23_clock = clock; // @[:@11183.4]
  assign RetimeWrapper_23_reset = reset; // @[:@11184.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@11186.4]
  assign RetimeWrapper_23_io_in = _T_1469 & io_rPort_1_en_0; // @[package.scala 94:16:@11185.4]
  assign RetimeWrapper_24_clock = clock; // @[:@11239.4]
  assign RetimeWrapper_24_reset = reset; // @[:@11240.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11242.4]
  assign RetimeWrapper_24_io_in = _T_463 & io_rPort_2_en_0; // @[package.scala 94:16:@11241.4]
  assign RetimeWrapper_25_clock = clock; // @[:@11247.4]
  assign RetimeWrapper_25_reset = reset; // @[:@11248.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11250.4]
  assign RetimeWrapper_25_io_in = _T_555 & io_rPort_2_en_0; // @[package.scala 94:16:@11249.4]
  assign RetimeWrapper_26_clock = clock; // @[:@11255.4]
  assign RetimeWrapper_26_reset = reset; // @[:@11256.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11258.4]
  assign RetimeWrapper_26_io_in = _T_647 & io_rPort_2_en_0; // @[package.scala 94:16:@11257.4]
  assign RetimeWrapper_27_clock = clock; // @[:@11263.4]
  assign RetimeWrapper_27_reset = reset; // @[:@11264.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11266.4]
  assign RetimeWrapper_27_io_in = _T_739 & io_rPort_2_en_0; // @[package.scala 94:16:@11265.4]
  assign RetimeWrapper_28_clock = clock; // @[:@11271.4]
  assign RetimeWrapper_28_reset = reset; // @[:@11272.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11274.4]
  assign RetimeWrapper_28_io_in = _T_831 & io_rPort_2_en_0; // @[package.scala 94:16:@11273.4]
  assign RetimeWrapper_29_clock = clock; // @[:@11279.4]
  assign RetimeWrapper_29_reset = reset; // @[:@11280.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11282.4]
  assign RetimeWrapper_29_io_in = _T_923 & io_rPort_2_en_0; // @[package.scala 94:16:@11281.4]
  assign RetimeWrapper_30_clock = clock; // @[:@11287.4]
  assign RetimeWrapper_30_reset = reset; // @[:@11288.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11290.4]
  assign RetimeWrapper_30_io_in = _T_1015 & io_rPort_2_en_0; // @[package.scala 94:16:@11289.4]
  assign RetimeWrapper_31_clock = clock; // @[:@11295.4]
  assign RetimeWrapper_31_reset = reset; // @[:@11296.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11298.4]
  assign RetimeWrapper_31_io_in = _T_1107 & io_rPort_2_en_0; // @[package.scala 94:16:@11297.4]
  assign RetimeWrapper_32_clock = clock; // @[:@11303.4]
  assign RetimeWrapper_32_reset = reset; // @[:@11304.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11306.4]
  assign RetimeWrapper_32_io_in = _T_1199 & io_rPort_2_en_0; // @[package.scala 94:16:@11305.4]
  assign RetimeWrapper_33_clock = clock; // @[:@11311.4]
  assign RetimeWrapper_33_reset = reset; // @[:@11312.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11314.4]
  assign RetimeWrapper_33_io_in = _T_1291 & io_rPort_2_en_0; // @[package.scala 94:16:@11313.4]
  assign RetimeWrapper_34_clock = clock; // @[:@11319.4]
  assign RetimeWrapper_34_reset = reset; // @[:@11320.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11322.4]
  assign RetimeWrapper_34_io_in = _T_1383 & io_rPort_2_en_0; // @[package.scala 94:16:@11321.4]
  assign RetimeWrapper_35_clock = clock; // @[:@11327.4]
  assign RetimeWrapper_35_reset = reset; // @[:@11328.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@11330.4]
  assign RetimeWrapper_35_io_in = _T_1475 & io_rPort_2_en_0; // @[package.scala 94:16:@11329.4]
  assign RetimeWrapper_36_clock = clock; // @[:@11383.4]
  assign RetimeWrapper_36_reset = reset; // @[:@11384.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11386.4]
  assign RetimeWrapper_36_io_in = _T_469 & io_rPort_3_en_0; // @[package.scala 94:16:@11385.4]
  assign RetimeWrapper_37_clock = clock; // @[:@11391.4]
  assign RetimeWrapper_37_reset = reset; // @[:@11392.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11394.4]
  assign RetimeWrapper_37_io_in = _T_561 & io_rPort_3_en_0; // @[package.scala 94:16:@11393.4]
  assign RetimeWrapper_38_clock = clock; // @[:@11399.4]
  assign RetimeWrapper_38_reset = reset; // @[:@11400.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11402.4]
  assign RetimeWrapper_38_io_in = _T_653 & io_rPort_3_en_0; // @[package.scala 94:16:@11401.4]
  assign RetimeWrapper_39_clock = clock; // @[:@11407.4]
  assign RetimeWrapper_39_reset = reset; // @[:@11408.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11410.4]
  assign RetimeWrapper_39_io_in = _T_745 & io_rPort_3_en_0; // @[package.scala 94:16:@11409.4]
  assign RetimeWrapper_40_clock = clock; // @[:@11415.4]
  assign RetimeWrapper_40_reset = reset; // @[:@11416.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11418.4]
  assign RetimeWrapper_40_io_in = _T_837 & io_rPort_3_en_0; // @[package.scala 94:16:@11417.4]
  assign RetimeWrapper_41_clock = clock; // @[:@11423.4]
  assign RetimeWrapper_41_reset = reset; // @[:@11424.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11426.4]
  assign RetimeWrapper_41_io_in = _T_929 & io_rPort_3_en_0; // @[package.scala 94:16:@11425.4]
  assign RetimeWrapper_42_clock = clock; // @[:@11431.4]
  assign RetimeWrapper_42_reset = reset; // @[:@11432.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11434.4]
  assign RetimeWrapper_42_io_in = _T_1021 & io_rPort_3_en_0; // @[package.scala 94:16:@11433.4]
  assign RetimeWrapper_43_clock = clock; // @[:@11439.4]
  assign RetimeWrapper_43_reset = reset; // @[:@11440.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11442.4]
  assign RetimeWrapper_43_io_in = _T_1113 & io_rPort_3_en_0; // @[package.scala 94:16:@11441.4]
  assign RetimeWrapper_44_clock = clock; // @[:@11447.4]
  assign RetimeWrapper_44_reset = reset; // @[:@11448.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11450.4]
  assign RetimeWrapper_44_io_in = _T_1205 & io_rPort_3_en_0; // @[package.scala 94:16:@11449.4]
  assign RetimeWrapper_45_clock = clock; // @[:@11455.4]
  assign RetimeWrapper_45_reset = reset; // @[:@11456.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11458.4]
  assign RetimeWrapper_45_io_in = _T_1297 & io_rPort_3_en_0; // @[package.scala 94:16:@11457.4]
  assign RetimeWrapper_46_clock = clock; // @[:@11463.4]
  assign RetimeWrapper_46_reset = reset; // @[:@11464.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11466.4]
  assign RetimeWrapper_46_io_in = _T_1389 & io_rPort_3_en_0; // @[package.scala 94:16:@11465.4]
  assign RetimeWrapper_47_clock = clock; // @[:@11471.4]
  assign RetimeWrapper_47_reset = reset; // @[:@11472.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@11474.4]
  assign RetimeWrapper_47_io_in = _T_1481 & io_rPort_3_en_0; // @[package.scala 94:16:@11473.4]
  assign RetimeWrapper_48_clock = clock; // @[:@11527.4]
  assign RetimeWrapper_48_reset = reset; // @[:@11528.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11530.4]
  assign RetimeWrapper_48_io_in = _T_475 & io_rPort_4_en_0; // @[package.scala 94:16:@11529.4]
  assign RetimeWrapper_49_clock = clock; // @[:@11535.4]
  assign RetimeWrapper_49_reset = reset; // @[:@11536.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11538.4]
  assign RetimeWrapper_49_io_in = _T_567 & io_rPort_4_en_0; // @[package.scala 94:16:@11537.4]
  assign RetimeWrapper_50_clock = clock; // @[:@11543.4]
  assign RetimeWrapper_50_reset = reset; // @[:@11544.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11546.4]
  assign RetimeWrapper_50_io_in = _T_659 & io_rPort_4_en_0; // @[package.scala 94:16:@11545.4]
  assign RetimeWrapper_51_clock = clock; // @[:@11551.4]
  assign RetimeWrapper_51_reset = reset; // @[:@11552.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11554.4]
  assign RetimeWrapper_51_io_in = _T_751 & io_rPort_4_en_0; // @[package.scala 94:16:@11553.4]
  assign RetimeWrapper_52_clock = clock; // @[:@11559.4]
  assign RetimeWrapper_52_reset = reset; // @[:@11560.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11562.4]
  assign RetimeWrapper_52_io_in = _T_843 & io_rPort_4_en_0; // @[package.scala 94:16:@11561.4]
  assign RetimeWrapper_53_clock = clock; // @[:@11567.4]
  assign RetimeWrapper_53_reset = reset; // @[:@11568.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11570.4]
  assign RetimeWrapper_53_io_in = _T_935 & io_rPort_4_en_0; // @[package.scala 94:16:@11569.4]
  assign RetimeWrapper_54_clock = clock; // @[:@11575.4]
  assign RetimeWrapper_54_reset = reset; // @[:@11576.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11578.4]
  assign RetimeWrapper_54_io_in = _T_1027 & io_rPort_4_en_0; // @[package.scala 94:16:@11577.4]
  assign RetimeWrapper_55_clock = clock; // @[:@11583.4]
  assign RetimeWrapper_55_reset = reset; // @[:@11584.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11586.4]
  assign RetimeWrapper_55_io_in = _T_1119 & io_rPort_4_en_0; // @[package.scala 94:16:@11585.4]
  assign RetimeWrapper_56_clock = clock; // @[:@11591.4]
  assign RetimeWrapper_56_reset = reset; // @[:@11592.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11594.4]
  assign RetimeWrapper_56_io_in = _T_1211 & io_rPort_4_en_0; // @[package.scala 94:16:@11593.4]
  assign RetimeWrapper_57_clock = clock; // @[:@11599.4]
  assign RetimeWrapper_57_reset = reset; // @[:@11600.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11602.4]
  assign RetimeWrapper_57_io_in = _T_1303 & io_rPort_4_en_0; // @[package.scala 94:16:@11601.4]
  assign RetimeWrapper_58_clock = clock; // @[:@11607.4]
  assign RetimeWrapper_58_reset = reset; // @[:@11608.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11610.4]
  assign RetimeWrapper_58_io_in = _T_1395 & io_rPort_4_en_0; // @[package.scala 94:16:@11609.4]
  assign RetimeWrapper_59_clock = clock; // @[:@11615.4]
  assign RetimeWrapper_59_reset = reset; // @[:@11616.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11618.4]
  assign RetimeWrapper_59_io_in = _T_1487 & io_rPort_4_en_0; // @[package.scala 94:16:@11617.4]
  assign RetimeWrapper_60_clock = clock; // @[:@11671.4]
  assign RetimeWrapper_60_reset = reset; // @[:@11672.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11674.4]
  assign RetimeWrapper_60_io_in = _T_481 & io_rPort_5_en_0; // @[package.scala 94:16:@11673.4]
  assign RetimeWrapper_61_clock = clock; // @[:@11679.4]
  assign RetimeWrapper_61_reset = reset; // @[:@11680.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11682.4]
  assign RetimeWrapper_61_io_in = _T_573 & io_rPort_5_en_0; // @[package.scala 94:16:@11681.4]
  assign RetimeWrapper_62_clock = clock; // @[:@11687.4]
  assign RetimeWrapper_62_reset = reset; // @[:@11688.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11690.4]
  assign RetimeWrapper_62_io_in = _T_665 & io_rPort_5_en_0; // @[package.scala 94:16:@11689.4]
  assign RetimeWrapper_63_clock = clock; // @[:@11695.4]
  assign RetimeWrapper_63_reset = reset; // @[:@11696.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11698.4]
  assign RetimeWrapper_63_io_in = _T_757 & io_rPort_5_en_0; // @[package.scala 94:16:@11697.4]
  assign RetimeWrapper_64_clock = clock; // @[:@11703.4]
  assign RetimeWrapper_64_reset = reset; // @[:@11704.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11706.4]
  assign RetimeWrapper_64_io_in = _T_849 & io_rPort_5_en_0; // @[package.scala 94:16:@11705.4]
  assign RetimeWrapper_65_clock = clock; // @[:@11711.4]
  assign RetimeWrapper_65_reset = reset; // @[:@11712.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11714.4]
  assign RetimeWrapper_65_io_in = _T_941 & io_rPort_5_en_0; // @[package.scala 94:16:@11713.4]
  assign RetimeWrapper_66_clock = clock; // @[:@11719.4]
  assign RetimeWrapper_66_reset = reset; // @[:@11720.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11722.4]
  assign RetimeWrapper_66_io_in = _T_1033 & io_rPort_5_en_0; // @[package.scala 94:16:@11721.4]
  assign RetimeWrapper_67_clock = clock; // @[:@11727.4]
  assign RetimeWrapper_67_reset = reset; // @[:@11728.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11730.4]
  assign RetimeWrapper_67_io_in = _T_1125 & io_rPort_5_en_0; // @[package.scala 94:16:@11729.4]
  assign RetimeWrapper_68_clock = clock; // @[:@11735.4]
  assign RetimeWrapper_68_reset = reset; // @[:@11736.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11738.4]
  assign RetimeWrapper_68_io_in = _T_1217 & io_rPort_5_en_0; // @[package.scala 94:16:@11737.4]
  assign RetimeWrapper_69_clock = clock; // @[:@11743.4]
  assign RetimeWrapper_69_reset = reset; // @[:@11744.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11746.4]
  assign RetimeWrapper_69_io_in = _T_1309 & io_rPort_5_en_0; // @[package.scala 94:16:@11745.4]
  assign RetimeWrapper_70_clock = clock; // @[:@11751.4]
  assign RetimeWrapper_70_reset = reset; // @[:@11752.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11754.4]
  assign RetimeWrapper_70_io_in = _T_1401 & io_rPort_5_en_0; // @[package.scala 94:16:@11753.4]
  assign RetimeWrapper_71_clock = clock; // @[:@11759.4]
  assign RetimeWrapper_71_reset = reset; // @[:@11760.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11762.4]
  assign RetimeWrapper_71_io_in = _T_1493 & io_rPort_5_en_0; // @[package.scala 94:16:@11761.4]
  assign RetimeWrapper_72_clock = clock; // @[:@11815.4]
  assign RetimeWrapper_72_reset = reset; // @[:@11816.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11818.4]
  assign RetimeWrapper_72_io_in = _T_487 & io_rPort_6_en_0; // @[package.scala 94:16:@11817.4]
  assign RetimeWrapper_73_clock = clock; // @[:@11823.4]
  assign RetimeWrapper_73_reset = reset; // @[:@11824.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11826.4]
  assign RetimeWrapper_73_io_in = _T_579 & io_rPort_6_en_0; // @[package.scala 94:16:@11825.4]
  assign RetimeWrapper_74_clock = clock; // @[:@11831.4]
  assign RetimeWrapper_74_reset = reset; // @[:@11832.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11834.4]
  assign RetimeWrapper_74_io_in = _T_671 & io_rPort_6_en_0; // @[package.scala 94:16:@11833.4]
  assign RetimeWrapper_75_clock = clock; // @[:@11839.4]
  assign RetimeWrapper_75_reset = reset; // @[:@11840.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11842.4]
  assign RetimeWrapper_75_io_in = _T_763 & io_rPort_6_en_0; // @[package.scala 94:16:@11841.4]
  assign RetimeWrapper_76_clock = clock; // @[:@11847.4]
  assign RetimeWrapper_76_reset = reset; // @[:@11848.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11850.4]
  assign RetimeWrapper_76_io_in = _T_855 & io_rPort_6_en_0; // @[package.scala 94:16:@11849.4]
  assign RetimeWrapper_77_clock = clock; // @[:@11855.4]
  assign RetimeWrapper_77_reset = reset; // @[:@11856.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11858.4]
  assign RetimeWrapper_77_io_in = _T_947 & io_rPort_6_en_0; // @[package.scala 94:16:@11857.4]
  assign RetimeWrapper_78_clock = clock; // @[:@11863.4]
  assign RetimeWrapper_78_reset = reset; // @[:@11864.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11866.4]
  assign RetimeWrapper_78_io_in = _T_1039 & io_rPort_6_en_0; // @[package.scala 94:16:@11865.4]
  assign RetimeWrapper_79_clock = clock; // @[:@11871.4]
  assign RetimeWrapper_79_reset = reset; // @[:@11872.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11874.4]
  assign RetimeWrapper_79_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@11873.4]
  assign RetimeWrapper_80_clock = clock; // @[:@11879.4]
  assign RetimeWrapper_80_reset = reset; // @[:@11880.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11882.4]
  assign RetimeWrapper_80_io_in = _T_1223 & io_rPort_6_en_0; // @[package.scala 94:16:@11881.4]
  assign RetimeWrapper_81_clock = clock; // @[:@11887.4]
  assign RetimeWrapper_81_reset = reset; // @[:@11888.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11890.4]
  assign RetimeWrapper_81_io_in = _T_1315 & io_rPort_6_en_0; // @[package.scala 94:16:@11889.4]
  assign RetimeWrapper_82_clock = clock; // @[:@11895.4]
  assign RetimeWrapper_82_reset = reset; // @[:@11896.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11898.4]
  assign RetimeWrapper_82_io_in = _T_1407 & io_rPort_6_en_0; // @[package.scala 94:16:@11897.4]
  assign RetimeWrapper_83_clock = clock; // @[:@11903.4]
  assign RetimeWrapper_83_reset = reset; // @[:@11904.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11906.4]
  assign RetimeWrapper_83_io_in = _T_1499 & io_rPort_6_en_0; // @[package.scala 94:16:@11905.4]
  assign RetimeWrapper_84_clock = clock; // @[:@11959.4]
  assign RetimeWrapper_84_reset = reset; // @[:@11960.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11962.4]
  assign RetimeWrapper_84_io_in = _T_493 & io_rPort_7_en_0; // @[package.scala 94:16:@11961.4]
  assign RetimeWrapper_85_clock = clock; // @[:@11967.4]
  assign RetimeWrapper_85_reset = reset; // @[:@11968.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11970.4]
  assign RetimeWrapper_85_io_in = _T_585 & io_rPort_7_en_0; // @[package.scala 94:16:@11969.4]
  assign RetimeWrapper_86_clock = clock; // @[:@11975.4]
  assign RetimeWrapper_86_reset = reset; // @[:@11976.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11978.4]
  assign RetimeWrapper_86_io_in = _T_677 & io_rPort_7_en_0; // @[package.scala 94:16:@11977.4]
  assign RetimeWrapper_87_clock = clock; // @[:@11983.4]
  assign RetimeWrapper_87_reset = reset; // @[:@11984.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11986.4]
  assign RetimeWrapper_87_io_in = _T_769 & io_rPort_7_en_0; // @[package.scala 94:16:@11985.4]
  assign RetimeWrapper_88_clock = clock; // @[:@11991.4]
  assign RetimeWrapper_88_reset = reset; // @[:@11992.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11994.4]
  assign RetimeWrapper_88_io_in = _T_861 & io_rPort_7_en_0; // @[package.scala 94:16:@11993.4]
  assign RetimeWrapper_89_clock = clock; // @[:@11999.4]
  assign RetimeWrapper_89_reset = reset; // @[:@12000.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@12002.4]
  assign RetimeWrapper_89_io_in = _T_953 & io_rPort_7_en_0; // @[package.scala 94:16:@12001.4]
  assign RetimeWrapper_90_clock = clock; // @[:@12007.4]
  assign RetimeWrapper_90_reset = reset; // @[:@12008.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@12010.4]
  assign RetimeWrapper_90_io_in = _T_1045 & io_rPort_7_en_0; // @[package.scala 94:16:@12009.4]
  assign RetimeWrapper_91_clock = clock; // @[:@12015.4]
  assign RetimeWrapper_91_reset = reset; // @[:@12016.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@12018.4]
  assign RetimeWrapper_91_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@12017.4]
  assign RetimeWrapper_92_clock = clock; // @[:@12023.4]
  assign RetimeWrapper_92_reset = reset; // @[:@12024.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@12026.4]
  assign RetimeWrapper_92_io_in = _T_1229 & io_rPort_7_en_0; // @[package.scala 94:16:@12025.4]
  assign RetimeWrapper_93_clock = clock; // @[:@12031.4]
  assign RetimeWrapper_93_reset = reset; // @[:@12032.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@12034.4]
  assign RetimeWrapper_93_io_in = _T_1321 & io_rPort_7_en_0; // @[package.scala 94:16:@12033.4]
  assign RetimeWrapper_94_clock = clock; // @[:@12039.4]
  assign RetimeWrapper_94_reset = reset; // @[:@12040.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@12042.4]
  assign RetimeWrapper_94_io_in = _T_1413 & io_rPort_7_en_0; // @[package.scala 94:16:@12041.4]
  assign RetimeWrapper_95_clock = clock; // @[:@12047.4]
  assign RetimeWrapper_95_reset = reset; // @[:@12048.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@12050.4]
  assign RetimeWrapper_95_io_in = _T_1505 & io_rPort_7_en_0; // @[package.scala 94:16:@12049.4]
  assign RetimeWrapper_96_clock = clock; // @[:@12103.4]
  assign RetimeWrapper_96_reset = reset; // @[:@12104.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12106.4]
  assign RetimeWrapper_96_io_in = _T_499 & io_rPort_8_en_0; // @[package.scala 94:16:@12105.4]
  assign RetimeWrapper_97_clock = clock; // @[:@12111.4]
  assign RetimeWrapper_97_reset = reset; // @[:@12112.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12114.4]
  assign RetimeWrapper_97_io_in = _T_591 & io_rPort_8_en_0; // @[package.scala 94:16:@12113.4]
  assign RetimeWrapper_98_clock = clock; // @[:@12119.4]
  assign RetimeWrapper_98_reset = reset; // @[:@12120.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12122.4]
  assign RetimeWrapper_98_io_in = _T_683 & io_rPort_8_en_0; // @[package.scala 94:16:@12121.4]
  assign RetimeWrapper_99_clock = clock; // @[:@12127.4]
  assign RetimeWrapper_99_reset = reset; // @[:@12128.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12130.4]
  assign RetimeWrapper_99_io_in = _T_775 & io_rPort_8_en_0; // @[package.scala 94:16:@12129.4]
  assign RetimeWrapper_100_clock = clock; // @[:@12135.4]
  assign RetimeWrapper_100_reset = reset; // @[:@12136.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12138.4]
  assign RetimeWrapper_100_io_in = _T_867 & io_rPort_8_en_0; // @[package.scala 94:16:@12137.4]
  assign RetimeWrapper_101_clock = clock; // @[:@12143.4]
  assign RetimeWrapper_101_reset = reset; // @[:@12144.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12146.4]
  assign RetimeWrapper_101_io_in = _T_959 & io_rPort_8_en_0; // @[package.scala 94:16:@12145.4]
  assign RetimeWrapper_102_clock = clock; // @[:@12151.4]
  assign RetimeWrapper_102_reset = reset; // @[:@12152.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12154.4]
  assign RetimeWrapper_102_io_in = _T_1051 & io_rPort_8_en_0; // @[package.scala 94:16:@12153.4]
  assign RetimeWrapper_103_clock = clock; // @[:@12159.4]
  assign RetimeWrapper_103_reset = reset; // @[:@12160.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12162.4]
  assign RetimeWrapper_103_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@12161.4]
  assign RetimeWrapper_104_clock = clock; // @[:@12167.4]
  assign RetimeWrapper_104_reset = reset; // @[:@12168.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12170.4]
  assign RetimeWrapper_104_io_in = _T_1235 & io_rPort_8_en_0; // @[package.scala 94:16:@12169.4]
  assign RetimeWrapper_105_clock = clock; // @[:@12175.4]
  assign RetimeWrapper_105_reset = reset; // @[:@12176.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12178.4]
  assign RetimeWrapper_105_io_in = _T_1327 & io_rPort_8_en_0; // @[package.scala 94:16:@12177.4]
  assign RetimeWrapper_106_clock = clock; // @[:@12183.4]
  assign RetimeWrapper_106_reset = reset; // @[:@12184.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12186.4]
  assign RetimeWrapper_106_io_in = _T_1419 & io_rPort_8_en_0; // @[package.scala 94:16:@12185.4]
  assign RetimeWrapper_107_clock = clock; // @[:@12191.4]
  assign RetimeWrapper_107_reset = reset; // @[:@12192.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@12194.4]
  assign RetimeWrapper_107_io_in = _T_1511 & io_rPort_8_en_0; // @[package.scala 94:16:@12193.4]
endmodule
module RetimeWrapper_140( // @[:@12222.2]
  input        clock, // @[:@12223.4]
  input        reset, // @[:@12224.4]
  input        io_flow, // @[:@12225.4]
  input  [7:0] io_in, // @[:@12225.4]
  output [7:0] io_out // @[:@12225.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12227.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12227.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12227.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12227.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12227.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12227.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@12227.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12240.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12239.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@12238.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12237.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12236.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12234.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@12242.2]
  input  [31:0] io_a, // @[:@12245.4]
  output [32:0] io_b // @[:@12245.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@12255.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@12255.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@12260.4]
endmodule
module __2( // @[:@12262.2]
  input  [31:0] io_b, // @[:@12265.4]
  output [32:0] io_result // @[:@12265.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@12270.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@12270.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@12270.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@12283.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@12278.4]
endmodule
module RetimeWrapper_141( // @[:@12340.2]
  input         clock, // @[:@12341.4]
  input         reset, // @[:@12342.4]
  input         io_flow, // @[:@12343.4]
  input  [31:0] io_in, // @[:@12343.4]
  output [31:0] io_out // @[:@12343.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12345.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12345.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12345.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12345.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12345.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12345.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@12345.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12358.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12357.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12356.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12355.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12354.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12352.4]
endmodule
module fix2fixBox( // @[:@12360.2]
  input         clock, // @[:@12361.4]
  input         reset, // @[:@12362.4]
  input  [32:0] io_a, // @[:@12363.4]
  input         io_flow, // @[:@12363.4]
  output [31:0] io_b // @[:@12363.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@12376.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@12376.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@12376.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@12376.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@12376.4]
  RetimeWrapper_141 RetimeWrapper ( // @[package.scala 93:22:@12376.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@12383.4]
  assign RetimeWrapper_clock = clock; // @[:@12377.4]
  assign RetimeWrapper_reset = reset; // @[:@12378.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@12380.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@12379.4]
endmodule
module x396_sum( // @[:@12385.2]
  input         clock, // @[:@12386.4]
  input         reset, // @[:@12387.4]
  input  [31:0] io_a, // @[:@12388.4]
  input  [31:0] io_b, // @[:@12388.4]
  input         io_flow, // @[:@12388.4]
  output [31:0] io_result // @[:@12388.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@12396.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@12396.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@12403.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@12403.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@12421.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@12421.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@12421.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@12421.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@12421.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@12401.4 Math.scala 713:14:@12402.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@12408.4 Math.scala 713:14:@12409.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@12410.4]
  __2 _ ( // @[Math.scala 709:24:@12396.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@12403.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@12421.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@12401.4 Math.scala 713:14:@12402.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@12408.4 Math.scala 713:14:@12409.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@12410.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@12429.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@12399.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@12406.4]
  assign fix2fixBox_clock = clock; // @[:@12422.4]
  assign fix2fixBox_reset = reset; // @[:@12423.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@12424.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@12427.4]
endmodule
module x414_sub( // @[:@13583.2]
  input         clock, // @[:@13584.4]
  input         reset, // @[:@13585.4]
  input  [31:0] io_a, // @[:@13586.4]
  input  [31:0] io_b, // @[:@13586.4]
  input         io_flow, // @[:@13586.4]
  output [31:0] io_result // @[:@13586.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@13594.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@13594.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@13601.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@13601.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@13620.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@13620.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@13620.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@13620.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@13620.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@13599.4 Math.scala 713:14:@13600.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@13606.4 Math.scala 713:14:@13607.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@13608.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@13609.4]
  __2 _ ( // @[Math.scala 709:24:@13594.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@13601.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@13620.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@13599.4 Math.scala 713:14:@13600.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@13606.4 Math.scala 713:14:@13607.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@13608.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@13609.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@13628.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@13597.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@13604.4]
  assign fix2fixBox_clock = clock; // @[:@13621.4]
  assign fix2fixBox_reset = reset; // @[:@13622.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@13623.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@13626.4]
endmodule
module RetimeWrapper_153( // @[:@13738.2]
  input         clock, // @[:@13739.4]
  input         reset, // @[:@13740.4]
  input         io_flow, // @[:@13741.4]
  input  [31:0] io_in, // @[:@13741.4]
  output [31:0] io_out // @[:@13741.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13743.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13743.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13743.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13743.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13743.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13743.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@13743.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13756.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13755.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@13754.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13753.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13752.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13750.4]
endmodule
module x232_div( // @[:@13799.2]
  input         clock, // @[:@13800.4]
  input         reset, // @[:@13801.4]
  input  [31:0] io_a, // @[:@13802.4]
  input         io_flow, // @[:@13802.4]
  output [31:0] io_result // @[:@13802.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13811.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13811.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13811.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@13811.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@13811.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@13824.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@13824.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@13808.4]
  wire [32:0] _T_17; // @[BigIPSim.scala 23:39:@13810.4]
  wire [32:0] _T_18; // @[package.scala 94:23:@13814.4]
  wire [31:0] _T_21; // @[package.scala 96:25:@13818.4]
  RetimeWrapper_153 RetimeWrapper ( // @[package.scala 93:22:@13811.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ _ ( // @[Math.scala 709:24:@13824.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@13808.4]
  assign _T_17 = $signed(_T_15) / $signed(32'sh3); // @[BigIPSim.scala 23:39:@13810.4]
  assign _T_18 = $unsigned(_T_17); // @[package.scala 94:23:@13814.4]
  assign _T_21 = $signed(RetimeWrapper_io_out); // @[package.scala 96:25:@13818.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@13832.4]
  assign RetimeWrapper_clock = clock; // @[:@13812.4]
  assign RetimeWrapper_reset = reset; // @[:@13813.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@13816.4]
  assign RetimeWrapper_io_in = _T_18[31:0]; // @[package.scala 94:16:@13815.4]
  assign __io_b = $unsigned(_T_21); // @[Math.scala 710:17:@13827.4]
endmodule
module RetimeWrapper_155( // @[:@13878.2]
  input         clock, // @[:@13879.4]
  input         reset, // @[:@13880.4]
  input         io_flow, // @[:@13881.4]
  input  [63:0] io_in, // @[:@13881.4]
  output [63:0] io_out // @[:@13881.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13883.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13883.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13883.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13883.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13883.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13883.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@13883.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13896.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13895.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@13894.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13893.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13892.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13890.4]
endmodule
module RetimeWrapper_156( // @[:@13910.2]
  input   clock, // @[:@13911.4]
  input   reset, // @[:@13912.4]
  input   io_flow, // @[:@13913.4]
  input   io_in // @[:@13913.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@13915.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@13915.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@13915.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13915.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13915.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13915.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@13915.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13927.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@13926.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13925.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13924.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13922.4]
endmodule
module fmamul_x416( // @[:@13980.2]
  input         clock, // @[:@13981.4]
  input         reset, // @[:@13982.4]
  input  [31:0] io_a, // @[:@13983.4]
  input         io_flow, // @[:@13983.4]
  output [31:0] io_result // @[:@13983.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13991.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13991.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13991.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@13991.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@13991.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14004.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14004.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14004.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14004.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14015.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14015.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14015.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14015.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@14022.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@14022.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@13996.4 package.scala 96:25:@13997.4]
  wire  _T_21; // @[FixedPoint.scala 50:25:@14001.4]
  RetimeWrapper_155 RetimeWrapper ( // @[package.scala 93:22:@13991.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_1 ( // @[package.scala 93:22:@14004.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in)
  );
  RetimeWrapper_156 RetimeWrapper_2 ( // @[package.scala 93:22:@14015.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in)
  );
  SimBlackBoxesfix2fixBox fix2fixBox ( // @[Math.scala 253:30:@14022.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@13996.4 package.scala 96:25:@13997.4]
  assign _T_21 = io_a[31]; // @[FixedPoint.scala 50:25:@14001.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@14030.4]
  assign RetimeWrapper_clock = clock; // @[:@13992.4]
  assign RetimeWrapper_reset = reset; // @[:@13993.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@13995.4]
  assign RetimeWrapper_io_in = io_a * 32'h156; // @[package.scala 94:16:@13994.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14005.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14006.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@14008.4]
  assign RetimeWrapper_1_io_in = io_a[31]; // @[package.scala 94:16:@14007.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14016.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14017.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@14019.4]
  assign RetimeWrapper_2_io_in = _T_21 == 1'h0; // @[package.scala 94:16:@14018.4]
  assign fix2fixBox_io_a = _T_18[31:0]; // @[Math.scala 254:23:@14025.4]
endmodule
module RetimeWrapper_158( // @[:@14044.2]
  input         clock, // @[:@14045.4]
  input         reset, // @[:@14046.4]
  input         io_flow, // @[:@14047.4]
  input  [31:0] io_in, // @[:@14047.4]
  output [31:0] io_out // @[:@14047.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14049.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14049.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14049.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14049.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14049.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14049.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@14049.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14062.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14061.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14060.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14059.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14058.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14056.4]
endmodule
module fix2fixBox_8( // @[:@14150.2]
  input  [32:0] io_a, // @[:@14153.4]
  output [31:0] io_b // @[:@14153.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@14166.4]
endmodule
module add( // @[:@14168.2]
  input  [31:0] io_a, // @[:@14171.4]
  input  [31:0] io_b, // @[:@14171.4]
  output [31:0] io_result // @[:@14171.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@14179.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@14179.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@14186.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@14186.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@14204.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@14204.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@14184.4 Math.scala 713:14:@14185.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@14191.4 Math.scala 713:14:@14192.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@14193.4]
  __2 _ ( // @[Math.scala 709:24:@14179.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@14186.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_8 fix2fixBox ( // @[Math.scala 141:30:@14204.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@14184.4 Math.scala 713:14:@14185.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@14191.4 Math.scala 713:14:@14192.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@14193.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@14212.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@14182.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@14189.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@14207.4]
endmodule
module x416( // @[:@14214.2]
  input         clock, // @[:@14215.4]
  input         reset, // @[:@14216.4]
  input  [31:0] io_m0, // @[:@14217.4]
  input  [31:0] io_add, // @[:@14217.4]
  input         io_flow, // @[:@14217.4]
  output [31:0] io_result // @[:@14217.4]
);
  wire  fmamul_x416_clock; // @[Math.scala 262:24:@14225.4]
  wire  fmamul_x416_reset; // @[Math.scala 262:24:@14225.4]
  wire [31:0] fmamul_x416_io_a; // @[Math.scala 262:24:@14225.4]
  wire  fmamul_x416_io_flow; // @[Math.scala 262:24:@14225.4]
  wire [31:0] fmamul_x416_io_result; // @[Math.scala 262:24:@14225.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14233.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14233.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14233.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@14233.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@14233.4]
  wire [31:0] add_1_io_a; // @[Math.scala 150:24:@14243.4]
  wire [31:0] add_1_io_b; // @[Math.scala 150:24:@14243.4]
  wire [31:0] add_1_io_result; // @[Math.scala 150:24:@14243.4]
  fmamul_x416 fmamul_x416 ( // @[Math.scala 262:24:@14225.4]
    .clock(fmamul_x416_clock),
    .reset(fmamul_x416_reset),
    .io_a(fmamul_x416_io_a),
    .io_flow(fmamul_x416_io_flow),
    .io_result(fmamul_x416_io_result)
  );
  RetimeWrapper_158 RetimeWrapper ( // @[package.scala 93:22:@14233.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  add add_1 ( // @[Math.scala 150:24:@14243.4]
    .io_a(add_1_io_a),
    .io_b(add_1_io_b),
    .io_result(add_1_io_result)
  );
  assign io_result = add_1_io_result; // @[Math.scala 846:17:@14251.4]
  assign fmamul_x416_clock = clock; // @[:@14226.4]
  assign fmamul_x416_reset = reset; // @[:@14227.4]
  assign fmamul_x416_io_a = io_m0; // @[Math.scala 263:17:@14228.4]
  assign fmamul_x416_io_flow = io_flow; // @[Math.scala 265:20:@14230.4]
  assign RetimeWrapper_clock = clock; // @[:@14234.4]
  assign RetimeWrapper_reset = reset; // @[:@14235.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@14237.4]
  assign RetimeWrapper_io_in = io_add; // @[package.scala 94:16:@14236.4]
  assign add_1_io_a = fmamul_x416_io_result; // @[Math.scala 151:17:@14246.4]
  assign add_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@14247.4]
endmodule
module RetimeWrapper_159( // @[:@14306.2]
  input   clock, // @[:@14307.4]
  input   reset, // @[:@14308.4]
  input   io_flow, // @[:@14309.4]
  input   io_in, // @[:@14309.4]
  output  io_out // @[:@14309.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@14311.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@14311.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@14311.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14311.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14311.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14311.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@14311.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14324.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14323.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@14322.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14321.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14320.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14318.4]
endmodule
module RetimeWrapper_161( // @[:@14370.2]
  input         clock, // @[:@14371.4]
  input         reset, // @[:@14372.4]
  input         io_flow, // @[:@14373.4]
  input  [31:0] io_in, // @[:@14373.4]
  output [31:0] io_out // @[:@14373.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14375.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14375.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14375.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14375.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14375.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14375.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@14375.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14388.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14387.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14386.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14385.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14384.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14382.4]
endmodule
module RetimeWrapper_162( // @[:@14402.2]
  input         clock, // @[:@14403.4]
  input         reset, // @[:@14404.4]
  input         io_flow, // @[:@14405.4]
  input  [31:0] io_in, // @[:@14405.4]
  output [31:0] io_out // @[:@14405.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14407.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14407.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14407.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14407.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14407.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14407.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@14407.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14420.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14419.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14418.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14417.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14416.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14414.4]
endmodule
module RetimeWrapper_163( // @[:@14434.2]
  input        clock, // @[:@14435.4]
  input        reset, // @[:@14436.4]
  input        io_flow, // @[:@14437.4]
  input  [7:0] io_in, // @[:@14437.4]
  output [7:0] io_out // @[:@14437.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14439.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14439.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14439.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14439.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14439.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14439.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(25)) sr ( // @[RetimeShiftRegister.scala 15:20:@14439.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14452.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14451.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@14450.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14449.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14448.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14446.4]
endmodule
module RetimeWrapper_165( // @[:@14498.2]
  input         clock, // @[:@14499.4]
  input         reset, // @[:@14500.4]
  input         io_flow, // @[:@14501.4]
  input  [31:0] io_in, // @[:@14501.4]
  output [31:0] io_out // @[:@14501.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14503.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14503.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14503.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14503.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14503.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14503.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(28)) sr ( // @[RetimeShiftRegister.scala 15:20:@14503.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14516.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14515.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14514.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14513.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14512.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14510.4]
endmodule
module RetimeWrapper_166( // @[:@14530.2]
  input         clock, // @[:@14531.4]
  input         reset, // @[:@14532.4]
  input         io_flow, // @[:@14533.4]
  input  [31:0] io_in, // @[:@14533.4]
  output [31:0] io_out // @[:@14533.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14535.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14535.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14535.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14535.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14535.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14535.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@14535.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14548.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14547.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14546.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14545.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14544.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14542.4]
endmodule
module fix2fixBox_9( // @[:@14550.2]
  input  [63:0] io_a, // @[:@14553.4]
  output [31:0] io_b // @[:@14553.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@14566.4]
endmodule
module x236( // @[:@14568.2]
  input         clock, // @[:@14569.4]
  input         reset, // @[:@14570.4]
  input  [31:0] io_a, // @[:@14571.4]
  input         io_flow, // @[:@14571.4]
  output [31:0] io_result // @[:@14571.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14580.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14580.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14580.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@14580.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@14580.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@14588.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@14588.4]
  wire [31:0] _T_19; // @[package.scala 96:25:@14585.4 package.scala 96:25:@14586.4]
  wire [31:0] _GEN_0; // @[package.scala 94:16:@14583.4]
  RetimeWrapper_166 RetimeWrapper ( // @[package.scala 93:22:@14580.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  fix2fixBox_9 fix2fixBox ( // @[Math.scala 357:30:@14588.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_19 = RetimeWrapper_io_out; // @[package.scala 96:25:@14585.4 package.scala 96:25:@14586.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@14596.4]
  assign RetimeWrapper_clock = clock; // @[:@14581.4]
  assign RetimeWrapper_reset = reset; // @[:@14582.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@14584.4]
  assign _GEN_0 = io_a % 32'h780; // @[package.scala 94:16:@14583.4]
  assign RetimeWrapper_io_in = _GEN_0[31:0]; // @[package.scala 94:16:@14583.4]
  assign fix2fixBox_io_a = {{32'd0}, _T_19}; // @[Math.scala 358:23:@14591.4]
endmodule
module RetimeWrapper_173( // @[:@14872.2]
  input         clock, // @[:@14873.4]
  input         reset, // @[:@14874.4]
  input         io_flow, // @[:@14875.4]
  input  [31:0] io_in, // @[:@14875.4]
  output [31:0] io_out // @[:@14875.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14877.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14877.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14877.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14877.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14877.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14877.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(30)) sr ( // @[RetimeShiftRegister.scala 15:20:@14877.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14890.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14889.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14888.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14887.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14886.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14884.4]
endmodule
module RetimeWrapper_175( // @[:@15093.2]
  input   clock, // @[:@15094.4]
  input   reset, // @[:@15095.4]
  input   io_flow, // @[:@15096.4]
  input   io_in, // @[:@15096.4]
  output  io_out // @[:@15096.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15098.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15098.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15098.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15098.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15098.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15098.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(55)) sr ( // @[RetimeShiftRegister.scala 15:20:@15098.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15111.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15110.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15109.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15108.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15107.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15105.4]
endmodule
module RetimeWrapper_176( // @[:@15125.2]
  input         clock, // @[:@15126.4]
  input         reset, // @[:@15127.4]
  input         io_flow, // @[:@15128.4]
  input  [31:0] io_in, // @[:@15128.4]
  output [31:0] io_out // @[:@15128.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15130.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15130.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15130.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15130.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15130.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15130.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@15130.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15143.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15142.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15141.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15140.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15139.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15137.4]
endmodule
module RetimeWrapper_178( // @[:@15189.2]
  input         clock, // @[:@15190.4]
  input         reset, // @[:@15191.4]
  input         io_flow, // @[:@15192.4]
  input  [31:0] io_in, // @[:@15192.4]
  output [31:0] io_out // @[:@15192.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15194.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15194.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15194.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15194.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15194.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15194.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@15194.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15207.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15206.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15205.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15204.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15203.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15201.4]
endmodule
module RetimeWrapper_180( // @[:@15253.2]
  input         clock, // @[:@15254.4]
  input         reset, // @[:@15255.4]
  input         io_flow, // @[:@15256.4]
  input  [31:0] io_in, // @[:@15256.4]
  output [31:0] io_out // @[:@15256.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15258.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15258.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15258.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15258.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15258.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15258.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(47)) sr ( // @[RetimeShiftRegister.scala 15:20:@15258.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15271.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15270.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15269.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15268.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15267.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15265.4]
endmodule
module RetimeWrapper_202( // @[:@17448.2]
  input   clock, // @[:@17449.4]
  input   reset, // @[:@17450.4]
  input   io_flow, // @[:@17451.4]
  input   io_in, // @[:@17451.4]
  output  io_out // @[:@17451.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(25)) sr ( // @[RetimeShiftRegister.scala 15:20:@17453.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17466.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17465.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@17464.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17463.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17462.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17460.4]
endmodule
module RetimeWrapper_232( // @[:@20175.2]
  input         clock, // @[:@20176.4]
  input         reset, // @[:@20177.4]
  input         io_flow, // @[:@20178.4]
  input  [31:0] io_in, // @[:@20178.4]
  output [31:0] io_out // @[:@20178.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20180.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20180.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20180.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20180.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20180.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20180.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(31)) sr ( // @[RetimeShiftRegister.scala 15:20:@20180.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20193.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20192.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20191.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20190.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20189.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20187.4]
endmodule
module RetimeWrapper_235( // @[:@20428.2]
  input         clock, // @[:@20429.4]
  input         reset, // @[:@20430.4]
  input         io_flow, // @[:@20431.4]
  input  [31:0] io_in, // @[:@20431.4]
  output [31:0] io_out // @[:@20431.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20433.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20433.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20433.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20433.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20433.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20433.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(10)) sr ( // @[RetimeShiftRegister.scala 15:20:@20433.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20446.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20445.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20444.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20443.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20442.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20440.4]
endmodule
module RetimeWrapper_236( // @[:@20460.2]
  input         clock, // @[:@20461.4]
  input         reset, // @[:@20462.4]
  input         io_flow, // @[:@20463.4]
  input  [31:0] io_in, // @[:@20463.4]
  output [31:0] io_out // @[:@20463.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20465.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20465.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20465.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20465.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20465.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20465.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@20465.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20478.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20477.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20476.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20475.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20474.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20472.4]
endmodule
module RetimeWrapper_238( // @[:@20524.2]
  input         clock, // @[:@20525.4]
  input         reset, // @[:@20526.4]
  input         io_flow, // @[:@20527.4]
  input  [31:0] io_in, // @[:@20527.4]
  output [31:0] io_out // @[:@20527.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20529.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20529.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20529.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20529.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20529.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20529.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@20529.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20542.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20541.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20540.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20539.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20538.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20536.4]
endmodule
module SimBlackBoxesfix2fixBox_76( // @[:@22501.2]
  input  [7:0] io_a, // @[:@22504.4]
  output [8:0] io_b // @[:@22504.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@22518.4]
endmodule
module __75( // @[:@22520.2]
  input  [7:0] io_b, // @[:@22523.4]
  output [8:0] io_result // @[:@22523.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@22528.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@22528.4]
  SimBlackBoxesfix2fixBox_76 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@22528.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@22541.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@22536.4]
endmodule
module fix2fixBox_42( // @[:@22617.2]
  input        clock, // @[:@22618.4]
  input        reset, // @[:@22619.4]
  input  [8:0] io_a, // @[:@22620.4]
  input        io_flow, // @[:@22620.4]
  output [7:0] io_b // @[:@22620.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22633.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22633.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22633.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@22633.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@22633.4]
  RetimeWrapper_140 RetimeWrapper ( // @[package.scala 93:22:@22633.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@22640.4]
  assign RetimeWrapper_clock = clock; // @[:@22634.4]
  assign RetimeWrapper_reset = reset; // @[:@22635.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@22637.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@22636.4]
endmodule
module x312_x11( // @[:@22642.2]
  input        clock, // @[:@22643.4]
  input        reset, // @[:@22644.4]
  input  [7:0] io_a, // @[:@22645.4]
  input  [7:0] io_b, // @[:@22645.4]
  input        io_flow, // @[:@22645.4]
  output [7:0] io_result // @[:@22645.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22653.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22653.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22660.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22660.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@22670.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@22670.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22670.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@22670.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22670.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22658.4 Math.scala 713:14:@22659.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22665.4 Math.scala 713:14:@22666.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22667.4]
  __75 _ ( // @[Math.scala 709:24:@22653.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __75 __1 ( // @[Math.scala 709:24:@22660.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_42 fix2fixBox ( // @[Math.scala 141:30:@22670.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22658.4 Math.scala 713:14:@22659.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22665.4 Math.scala 713:14:@22666.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22667.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22678.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22656.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22663.4]
  assign fix2fixBox_clock = clock; // @[:@22671.4]
  assign fix2fixBox_reset = reset; // @[:@22672.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22673.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@22676.4]
endmodule
module fix2fixBox_46( // @[:@23301.2]
  input  [8:0] io_a, // @[:@23304.4]
  output [7:0] io_b // @[:@23304.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@23317.4]
endmodule
module x316_x11( // @[:@23319.2]
  input  [7:0] io_a, // @[:@23322.4]
  input  [7:0] io_b, // @[:@23322.4]
  output [7:0] io_result // @[:@23322.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@23330.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@23330.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@23337.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@23337.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@23347.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@23347.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@23335.4 Math.scala 713:14:@23336.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@23342.4 Math.scala 713:14:@23343.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@23344.4]
  __75 _ ( // @[Math.scala 709:24:@23330.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __75 __1 ( // @[Math.scala 709:24:@23337.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_46 fix2fixBox ( // @[Math.scala 141:30:@23347.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@23335.4 Math.scala 713:14:@23336.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@23342.4 Math.scala 713:14:@23343.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@23344.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@23355.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@23333.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@23340.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@23350.4]
endmodule
module RetimeWrapper_273( // @[:@23853.2]
  input        clock, // @[:@23854.4]
  input        reset, // @[:@23855.4]
  input        io_flow, // @[:@23856.4]
  input  [7:0] io_in, // @[:@23856.4]
  output [7:0] io_out // @[:@23856.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23858.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23858.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23858.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23858.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23858.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23858.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@23858.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23871.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23870.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@23869.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23868.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23867.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23865.4]
endmodule
module x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@23969.2]
  input          clock, // @[:@23970.4]
  input          reset, // @[:@23971.4]
  output         io_in_x206_TVALID, // @[:@23972.4]
  input          io_in_x206_TREADY, // @[:@23972.4]
  output [255:0] io_in_x206_TDATA, // @[:@23972.4]
  output         io_in_x205_TREADY, // @[:@23972.4]
  input  [255:0] io_in_x205_TDATA, // @[:@23972.4]
  input  [7:0]   io_in_x205_TID, // @[:@23972.4]
  input  [7:0]   io_in_x205_TDEST, // @[:@23972.4]
  input          io_sigsIn_backpressure, // @[:@23972.4]
  input          io_sigsIn_datapathEn, // @[:@23972.4]
  input          io_sigsIn_break, // @[:@23972.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@23972.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@23972.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@23972.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@23972.4]
  input          io_rr // @[:@23972.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@23986.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@23986.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@23998.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@23998.4]
  wire  x218_lb_0_clock; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_reset; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_8_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_8_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_8_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_8_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_8_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_8_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_7_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_7_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_7_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_7_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_7_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_7_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_6_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_6_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_6_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_6_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_6_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_6_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_5_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_5_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_5_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_5_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_5_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_5_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_4_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_4_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_4_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_4_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_4_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_4_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_3_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_3_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_3_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_3_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_3_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_3_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_2_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_2_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_2_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_2_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_2_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_2_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_1_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_1_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_1_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_1_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_1_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_1_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_rPort_0_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_rPort_0_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_rPort_0_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_0_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_rPort_0_backpressure; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_rPort_0_output_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [1:0] x218_lb_0_io_wPort_0_banks_1; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [2:0] x218_lb_0_io_wPort_0_banks_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [8:0] x218_lb_0_io_wPort_0_ofs_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire [7:0] x218_lb_0_io_wPort_0_data_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  x218_lb_0_io_wPort_0_en_0; // @[m_x218_lb_0.scala 35:17:@24008.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@24088.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@24088.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@24088.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@24088.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@24088.4]
  wire  x396_sum_1_clock; // @[Math.scala 150:24:@24184.4]
  wire  x396_sum_1_reset; // @[Math.scala 150:24:@24184.4]
  wire [31:0] x396_sum_1_io_a; // @[Math.scala 150:24:@24184.4]
  wire [31:0] x396_sum_1_io_b; // @[Math.scala 150:24:@24184.4]
  wire  x396_sum_1_io_flow; // @[Math.scala 150:24:@24184.4]
  wire [31:0] x396_sum_1_io_result; // @[Math.scala 150:24:@24184.4]
  wire  x399_sum_1_clock; // @[Math.scala 150:24:@24214.4]
  wire  x399_sum_1_reset; // @[Math.scala 150:24:@24214.4]
  wire [31:0] x399_sum_1_io_a; // @[Math.scala 150:24:@24214.4]
  wire [31:0] x399_sum_1_io_b; // @[Math.scala 150:24:@24214.4]
  wire  x399_sum_1_io_flow; // @[Math.scala 150:24:@24214.4]
  wire [31:0] x399_sum_1_io_result; // @[Math.scala 150:24:@24214.4]
  wire  x402_sum_1_clock; // @[Math.scala 150:24:@24244.4]
  wire  x402_sum_1_reset; // @[Math.scala 150:24:@24244.4]
  wire [31:0] x402_sum_1_io_a; // @[Math.scala 150:24:@24244.4]
  wire [31:0] x402_sum_1_io_b; // @[Math.scala 150:24:@24244.4]
  wire  x402_sum_1_io_flow; // @[Math.scala 150:24:@24244.4]
  wire [31:0] x402_sum_1_io_result; // @[Math.scala 150:24:@24244.4]
  wire  x405_sum_1_clock; // @[Math.scala 150:24:@24274.4]
  wire  x405_sum_1_reset; // @[Math.scala 150:24:@24274.4]
  wire [31:0] x405_sum_1_io_a; // @[Math.scala 150:24:@24274.4]
  wire [31:0] x405_sum_1_io_b; // @[Math.scala 150:24:@24274.4]
  wire  x405_sum_1_io_flow; // @[Math.scala 150:24:@24274.4]
  wire [31:0] x405_sum_1_io_result; // @[Math.scala 150:24:@24274.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@24290.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@24290.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@24290.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@24290.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@24290.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@24307.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@24307.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@24307.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@24307.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@24307.4]
  wire  x408_sum_1_clock; // @[Math.scala 150:24:@24320.4]
  wire  x408_sum_1_reset; // @[Math.scala 150:24:@24320.4]
  wire [31:0] x408_sum_1_io_a; // @[Math.scala 150:24:@24320.4]
  wire [31:0] x408_sum_1_io_b; // @[Math.scala 150:24:@24320.4]
  wire  x408_sum_1_io_flow; // @[Math.scala 150:24:@24320.4]
  wire [31:0] x408_sum_1_io_result; // @[Math.scala 150:24:@24320.4]
  wire  x411_sum_1_clock; // @[Math.scala 150:24:@24350.4]
  wire  x411_sum_1_reset; // @[Math.scala 150:24:@24350.4]
  wire [31:0] x411_sum_1_io_a; // @[Math.scala 150:24:@24350.4]
  wire [31:0] x411_sum_1_io_b; // @[Math.scala 150:24:@24350.4]
  wire  x411_sum_1_io_flow; // @[Math.scala 150:24:@24350.4]
  wire [31:0] x411_sum_1_io_result; // @[Math.scala 150:24:@24350.4]
  wire  x414_sub_1_clock; // @[Math.scala 191:24:@24376.4]
  wire  x414_sub_1_reset; // @[Math.scala 191:24:@24376.4]
  wire [31:0] x414_sub_1_io_a; // @[Math.scala 191:24:@24376.4]
  wire [31:0] x414_sub_1_io_b; // @[Math.scala 191:24:@24376.4]
  wire  x414_sub_1_io_flow; // @[Math.scala 191:24:@24376.4]
  wire [31:0] x414_sub_1_io_result; // @[Math.scala 191:24:@24376.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@24386.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@24386.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@24386.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@24386.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@24386.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@24395.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@24395.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@24395.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@24395.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@24395.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@24404.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@24404.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@24404.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@24404.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@24404.4]
  wire  x232_div_1_clock; // @[Math.scala 327:24:@24427.4]
  wire  x232_div_1_reset; // @[Math.scala 327:24:@24427.4]
  wire [31:0] x232_div_1_io_a; // @[Math.scala 327:24:@24427.4]
  wire  x232_div_1_io_flow; // @[Math.scala 327:24:@24427.4]
  wire [31:0] x232_div_1_io_result; // @[Math.scala 327:24:@24427.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@24437.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@24437.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@24437.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@24437.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@24437.4]
  wire  x416_1_clock; // @[Math.scala 849:24:@24448.4]
  wire  x416_1_reset; // @[Math.scala 849:24:@24448.4]
  wire [31:0] x416_1_io_m0; // @[Math.scala 849:24:@24448.4]
  wire [31:0] x416_1_io_add; // @[Math.scala 849:24:@24448.4]
  wire  x416_1_io_flow; // @[Math.scala 849:24:@24448.4]
  wire [31:0] x416_1_io_result; // @[Math.scala 849:24:@24448.4]
  wire [31:0] cast_x416_io_b; // @[Math.scala 709:24:@24457.4]
  wire [31:0] cast_x416_io_result; // @[Math.scala 709:24:@24457.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@24466.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@24466.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@24466.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@24466.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@24466.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@24475.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@24475.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@24475.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@24475.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@24475.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@24484.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@24484.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@24493.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@24493.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@24493.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@24493.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@24493.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@24502.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@24502.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@24502.4]
  wire [7:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@24502.4]
  wire [7:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@24502.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@24513.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@24513.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@24513.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@24513.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@24513.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@24534.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@24534.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@24534.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@24534.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@24534.4]
  wire  x236_1_clock; // @[Math.scala 366:24:@24547.4]
  wire  x236_1_reset; // @[Math.scala 366:24:@24547.4]
  wire [31:0] x236_1_io_a; // @[Math.scala 366:24:@24547.4]
  wire  x236_1_io_flow; // @[Math.scala 366:24:@24547.4]
  wire [31:0] x236_1_io_result; // @[Math.scala 366:24:@24547.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@24562.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@24562.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@24562.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@24562.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@24562.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@24571.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@24571.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@24585.4]
  wire  x243_mul_1_clock; // @[Math.scala 262:24:@24622.4]
  wire  x243_mul_1_reset; // @[Math.scala 262:24:@24622.4]
  wire [31:0] x243_mul_1_io_a; // @[Math.scala 262:24:@24622.4]
  wire  x243_mul_1_io_flow; // @[Math.scala 262:24:@24622.4]
  wire [31:0] x243_mul_1_io_result; // @[Math.scala 262:24:@24622.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@24632.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@24632.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@24632.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@24632.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@24632.4]
  wire  x244_sum_1_clock; // @[Math.scala 150:24:@24641.4]
  wire  x244_sum_1_reset; // @[Math.scala 150:24:@24641.4]
  wire [31:0] x244_sum_1_io_a; // @[Math.scala 150:24:@24641.4]
  wire [31:0] x244_sum_1_io_b; // @[Math.scala 150:24:@24641.4]
  wire  x244_sum_1_io_flow; // @[Math.scala 150:24:@24641.4]
  wire [31:0] x244_sum_1_io_result; // @[Math.scala 150:24:@24641.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@24651.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@24651.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@24651.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@24651.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@24651.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@24660.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@24660.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@24669.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@24669.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@24669.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@24669.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@24669.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@24678.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@24678.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@24678.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@24678.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@24678.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@24696.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@24696.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@24696.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@24696.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@24696.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@24708.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@24708.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@24708.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@24708.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@24708.4]
  wire  x247_rdcol_1_clock; // @[Math.scala 191:24:@24731.4]
  wire  x247_rdcol_1_reset; // @[Math.scala 191:24:@24731.4]
  wire [31:0] x247_rdcol_1_io_a; // @[Math.scala 191:24:@24731.4]
  wire [31:0] x247_rdcol_1_io_b; // @[Math.scala 191:24:@24731.4]
  wire  x247_rdcol_1_io_flow; // @[Math.scala 191:24:@24731.4]
  wire [31:0] x247_rdcol_1_io_result; // @[Math.scala 191:24:@24731.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@24746.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@24746.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@24746.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@24746.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@24746.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@24755.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@24755.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@24755.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@24755.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@24755.4]
  wire  x420_sum_1_clock; // @[Math.scala 150:24:@24790.4]
  wire  x420_sum_1_reset; // @[Math.scala 150:24:@24790.4]
  wire [31:0] x420_sum_1_io_a; // @[Math.scala 150:24:@24790.4]
  wire [31:0] x420_sum_1_io_b; // @[Math.scala 150:24:@24790.4]
  wire  x420_sum_1_io_flow; // @[Math.scala 150:24:@24790.4]
  wire [31:0] x420_sum_1_io_result; // @[Math.scala 150:24:@24790.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@24806.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@24806.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@24806.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@24806.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@24806.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@24823.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@24823.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@24823.4]
  wire  x423_sum_1_clock; // @[Math.scala 150:24:@24836.4]
  wire  x423_sum_1_reset; // @[Math.scala 150:24:@24836.4]
  wire [31:0] x423_sum_1_io_a; // @[Math.scala 150:24:@24836.4]
  wire [31:0] x423_sum_1_io_b; // @[Math.scala 150:24:@24836.4]
  wire  x423_sum_1_io_flow; // @[Math.scala 150:24:@24836.4]
  wire [31:0] x423_sum_1_io_result; // @[Math.scala 150:24:@24836.4]
  wire  x426_sum_1_clock; // @[Math.scala 150:24:@24866.4]
  wire  x426_sum_1_reset; // @[Math.scala 150:24:@24866.4]
  wire [31:0] x426_sum_1_io_a; // @[Math.scala 150:24:@24866.4]
  wire [31:0] x426_sum_1_io_b; // @[Math.scala 150:24:@24866.4]
  wire  x426_sum_1_io_flow; // @[Math.scala 150:24:@24866.4]
  wire [31:0] x426_sum_1_io_result; // @[Math.scala 150:24:@24866.4]
  wire  x429_sum_1_clock; // @[Math.scala 150:24:@24896.4]
  wire  x429_sum_1_reset; // @[Math.scala 150:24:@24896.4]
  wire [31:0] x429_sum_1_io_a; // @[Math.scala 150:24:@24896.4]
  wire [31:0] x429_sum_1_io_b; // @[Math.scala 150:24:@24896.4]
  wire  x429_sum_1_io_flow; // @[Math.scala 150:24:@24896.4]
  wire [31:0] x429_sum_1_io_result; // @[Math.scala 150:24:@24896.4]
  wire  x432_sum_1_clock; // @[Math.scala 150:24:@24926.4]
  wire  x432_sum_1_reset; // @[Math.scala 150:24:@24926.4]
  wire [31:0] x432_sum_1_io_a; // @[Math.scala 150:24:@24926.4]
  wire [31:0] x432_sum_1_io_b; // @[Math.scala 150:24:@24926.4]
  wire  x432_sum_1_io_flow; // @[Math.scala 150:24:@24926.4]
  wire [31:0] x432_sum_1_io_result; // @[Math.scala 150:24:@24926.4]
  wire  x435_sum_1_clock; // @[Math.scala 150:24:@24956.4]
  wire  x435_sum_1_reset; // @[Math.scala 150:24:@24956.4]
  wire [31:0] x435_sum_1_io_a; // @[Math.scala 150:24:@24956.4]
  wire [31:0] x435_sum_1_io_b; // @[Math.scala 150:24:@24956.4]
  wire  x435_sum_1_io_flow; // @[Math.scala 150:24:@24956.4]
  wire [31:0] x435_sum_1_io_result; // @[Math.scala 150:24:@24956.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@24971.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@24971.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@24971.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@24971.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@24971.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@24985.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@24985.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@24985.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@24985.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@24985.4]
  wire  x438_sub_1_clock; // @[Math.scala 191:24:@24996.4]
  wire  x438_sub_1_reset; // @[Math.scala 191:24:@24996.4]
  wire [31:0] x438_sub_1_io_a; // @[Math.scala 191:24:@24996.4]
  wire [31:0] x438_sub_1_io_b; // @[Math.scala 191:24:@24996.4]
  wire  x438_sub_1_io_flow; // @[Math.scala 191:24:@24996.4]
  wire [31:0] x438_sub_1_io_result; // @[Math.scala 191:24:@24996.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@25006.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@25006.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@25006.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@25006.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@25006.4]
  wire  x252_div_1_clock; // @[Math.scala 327:24:@25020.4]
  wire  x252_div_1_reset; // @[Math.scala 327:24:@25020.4]
  wire [31:0] x252_div_1_io_a; // @[Math.scala 327:24:@25020.4]
  wire  x252_div_1_io_flow; // @[Math.scala 327:24:@25020.4]
  wire [31:0] x252_div_1_io_result; // @[Math.scala 327:24:@25020.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@25030.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@25030.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@25030.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@25030.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@25030.4]
  wire  x253_sum_1_clock; // @[Math.scala 150:24:@25041.4]
  wire  x253_sum_1_reset; // @[Math.scala 150:24:@25041.4]
  wire [31:0] x253_sum_1_io_a; // @[Math.scala 150:24:@25041.4]
  wire [31:0] x253_sum_1_io_b; // @[Math.scala 150:24:@25041.4]
  wire  x253_sum_1_io_flow; // @[Math.scala 150:24:@25041.4]
  wire [31:0] x253_sum_1_io_result; // @[Math.scala 150:24:@25041.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@25051.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@25051.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@25051.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@25051.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@25051.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@25060.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@25060.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@25069.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@25069.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@25069.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@25069.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@25069.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@25081.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@25081.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@25081.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@25081.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@25081.4]
  wire  x256_rdcol_1_clock; // @[Math.scala 191:24:@25104.4]
  wire  x256_rdcol_1_reset; // @[Math.scala 191:24:@25104.4]
  wire [31:0] x256_rdcol_1_io_a; // @[Math.scala 191:24:@25104.4]
  wire [31:0] x256_rdcol_1_io_b; // @[Math.scala 191:24:@25104.4]
  wire  x256_rdcol_1_io_flow; // @[Math.scala 191:24:@25104.4]
  wire [31:0] x256_rdcol_1_io_result; // @[Math.scala 191:24:@25104.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@25119.4]
  wire  x442_sum_1_clock; // @[Math.scala 150:24:@25154.4]
  wire  x442_sum_1_reset; // @[Math.scala 150:24:@25154.4]
  wire [31:0] x442_sum_1_io_a; // @[Math.scala 150:24:@25154.4]
  wire [31:0] x442_sum_1_io_b; // @[Math.scala 150:24:@25154.4]
  wire  x442_sum_1_io_flow; // @[Math.scala 150:24:@25154.4]
  wire [31:0] x442_sum_1_io_result; // @[Math.scala 150:24:@25154.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@25170.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@25170.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@25170.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@25170.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@25170.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@25187.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@25187.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@25187.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@25187.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@25187.4]
  wire  x445_sum_1_clock; // @[Math.scala 150:24:@25200.4]
  wire  x445_sum_1_reset; // @[Math.scala 150:24:@25200.4]
  wire [31:0] x445_sum_1_io_a; // @[Math.scala 150:24:@25200.4]
  wire [31:0] x445_sum_1_io_b; // @[Math.scala 150:24:@25200.4]
  wire  x445_sum_1_io_flow; // @[Math.scala 150:24:@25200.4]
  wire [31:0] x445_sum_1_io_result; // @[Math.scala 150:24:@25200.4]
  wire  x448_sum_1_clock; // @[Math.scala 150:24:@25230.4]
  wire  x448_sum_1_reset; // @[Math.scala 150:24:@25230.4]
  wire [31:0] x448_sum_1_io_a; // @[Math.scala 150:24:@25230.4]
  wire [31:0] x448_sum_1_io_b; // @[Math.scala 150:24:@25230.4]
  wire  x448_sum_1_io_flow; // @[Math.scala 150:24:@25230.4]
  wire [31:0] x448_sum_1_io_result; // @[Math.scala 150:24:@25230.4]
  wire  x451_sum_1_clock; // @[Math.scala 150:24:@25260.4]
  wire  x451_sum_1_reset; // @[Math.scala 150:24:@25260.4]
  wire [31:0] x451_sum_1_io_a; // @[Math.scala 150:24:@25260.4]
  wire [31:0] x451_sum_1_io_b; // @[Math.scala 150:24:@25260.4]
  wire  x451_sum_1_io_flow; // @[Math.scala 150:24:@25260.4]
  wire [31:0] x451_sum_1_io_result; // @[Math.scala 150:24:@25260.4]
  wire  x454_sum_1_clock; // @[Math.scala 150:24:@25290.4]
  wire  x454_sum_1_reset; // @[Math.scala 150:24:@25290.4]
  wire [31:0] x454_sum_1_io_a; // @[Math.scala 150:24:@25290.4]
  wire [31:0] x454_sum_1_io_b; // @[Math.scala 150:24:@25290.4]
  wire  x454_sum_1_io_flow; // @[Math.scala 150:24:@25290.4]
  wire [31:0] x454_sum_1_io_result; // @[Math.scala 150:24:@25290.4]
  wire  x457_sum_1_clock; // @[Math.scala 150:24:@25320.4]
  wire  x457_sum_1_reset; // @[Math.scala 150:24:@25320.4]
  wire [31:0] x457_sum_1_io_a; // @[Math.scala 150:24:@25320.4]
  wire [31:0] x457_sum_1_io_b; // @[Math.scala 150:24:@25320.4]
  wire  x457_sum_1_io_flow; // @[Math.scala 150:24:@25320.4]
  wire [31:0] x457_sum_1_io_result; // @[Math.scala 150:24:@25320.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@25335.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@25335.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@25335.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@25335.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@25335.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@25349.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@25349.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@25349.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@25349.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@25349.4]
  wire  x460_sub_1_clock; // @[Math.scala 191:24:@25360.4]
  wire  x460_sub_1_reset; // @[Math.scala 191:24:@25360.4]
  wire [31:0] x460_sub_1_io_a; // @[Math.scala 191:24:@25360.4]
  wire [31:0] x460_sub_1_io_b; // @[Math.scala 191:24:@25360.4]
  wire  x460_sub_1_io_flow; // @[Math.scala 191:24:@25360.4]
  wire [31:0] x460_sub_1_io_result; // @[Math.scala 191:24:@25360.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@25370.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@25370.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@25370.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@25370.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@25370.4]
  wire  x261_div_1_clock; // @[Math.scala 327:24:@25384.4]
  wire  x261_div_1_reset; // @[Math.scala 327:24:@25384.4]
  wire [31:0] x261_div_1_io_a; // @[Math.scala 327:24:@25384.4]
  wire  x261_div_1_io_flow; // @[Math.scala 327:24:@25384.4]
  wire [31:0] x261_div_1_io_result; // @[Math.scala 327:24:@25384.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@25394.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@25394.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@25394.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@25394.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@25394.4]
  wire  x262_sum_1_clock; // @[Math.scala 150:24:@25403.4]
  wire  x262_sum_1_reset; // @[Math.scala 150:24:@25403.4]
  wire [31:0] x262_sum_1_io_a; // @[Math.scala 150:24:@25403.4]
  wire [31:0] x262_sum_1_io_b; // @[Math.scala 150:24:@25403.4]
  wire  x262_sum_1_io_flow; // @[Math.scala 150:24:@25403.4]
  wire [31:0] x262_sum_1_io_result; // @[Math.scala 150:24:@25403.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@25413.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@25413.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@25413.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@25413.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@25413.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@25422.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@25422.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@25422.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@25422.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@25422.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@25431.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@25431.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@25443.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@25443.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@25443.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@25443.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@25443.4]
  wire  x265_rdrow_1_clock; // @[Math.scala 191:24:@25466.4]
  wire  x265_rdrow_1_reset; // @[Math.scala 191:24:@25466.4]
  wire [31:0] x265_rdrow_1_io_a; // @[Math.scala 191:24:@25466.4]
  wire [31:0] x265_rdrow_1_io_b; // @[Math.scala 191:24:@25466.4]
  wire  x265_rdrow_1_io_flow; // @[Math.scala 191:24:@25466.4]
  wire [31:0] x265_rdrow_1_io_result; // @[Math.scala 191:24:@25466.4]
  wire  x266_1_clock; // @[Math.scala 366:24:@25478.4]
  wire  x266_1_reset; // @[Math.scala 366:24:@25478.4]
  wire [31:0] x266_1_io_a; // @[Math.scala 366:24:@25478.4]
  wire  x266_1_io_flow; // @[Math.scala 366:24:@25478.4]
  wire [31:0] x266_1_io_result; // @[Math.scala 366:24:@25478.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@25493.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@25493.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@25493.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@25493.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@25493.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@25502.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@25502.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@25502.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@25502.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@25502.4]
  wire  x272_mul_1_clock; // @[Math.scala 262:24:@25541.4]
  wire  x272_mul_1_reset; // @[Math.scala 262:24:@25541.4]
  wire [31:0] x272_mul_1_io_a; // @[Math.scala 262:24:@25541.4]
  wire  x272_mul_1_io_flow; // @[Math.scala 262:24:@25541.4]
  wire [31:0] x272_mul_1_io_result; // @[Math.scala 262:24:@25541.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@25551.4]
  wire [31:0] RetimeWrapper_50_io_in; // @[package.scala 93:22:@25551.4]
  wire [31:0] RetimeWrapper_50_io_out; // @[package.scala 93:22:@25551.4]
  wire  x273_sum_1_clock; // @[Math.scala 150:24:@25560.4]
  wire  x273_sum_1_reset; // @[Math.scala 150:24:@25560.4]
  wire [31:0] x273_sum_1_io_a; // @[Math.scala 150:24:@25560.4]
  wire [31:0] x273_sum_1_io_b; // @[Math.scala 150:24:@25560.4]
  wire  x273_sum_1_io_flow; // @[Math.scala 150:24:@25560.4]
  wire [31:0] x273_sum_1_io_result; // @[Math.scala 150:24:@25560.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@25570.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@25570.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@25570.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@25570.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@25570.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@25579.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@25579.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@25579.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@25579.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@25579.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@25588.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@25588.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@25600.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@25600.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@25600.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@25600.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@25600.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@25627.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@25627.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@25627.4]
  wire [31:0] RetimeWrapper_55_io_in; // @[package.scala 93:22:@25627.4]
  wire [31:0] RetimeWrapper_55_io_out; // @[package.scala 93:22:@25627.4]
  wire  x278_sum_1_clock; // @[Math.scala 150:24:@25636.4]
  wire  x278_sum_1_reset; // @[Math.scala 150:24:@25636.4]
  wire [31:0] x278_sum_1_io_a; // @[Math.scala 150:24:@25636.4]
  wire [31:0] x278_sum_1_io_b; // @[Math.scala 150:24:@25636.4]
  wire  x278_sum_1_io_flow; // @[Math.scala 150:24:@25636.4]
  wire [31:0] x278_sum_1_io_result; // @[Math.scala 150:24:@25636.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@25646.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@25646.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@25646.4]
  wire [31:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@25646.4]
  wire [31:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@25646.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@25667.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@25667.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@25667.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@25667.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@25667.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@25694.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@25694.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@25694.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@25694.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@25694.4]
  wire  x283_sum_1_clock; // @[Math.scala 150:24:@25703.4]
  wire  x283_sum_1_reset; // @[Math.scala 150:24:@25703.4]
  wire [31:0] x283_sum_1_io_a; // @[Math.scala 150:24:@25703.4]
  wire [31:0] x283_sum_1_io_b; // @[Math.scala 150:24:@25703.4]
  wire  x283_sum_1_io_flow; // @[Math.scala 150:24:@25703.4]
  wire [31:0] x283_sum_1_io_result; // @[Math.scala 150:24:@25703.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@25713.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@25713.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@25713.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@25713.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@25713.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@25722.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@25722.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@25722.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@25722.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@25722.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@25734.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@25734.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@25734.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@25734.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@25734.4]
  wire  x286_rdrow_1_clock; // @[Math.scala 191:24:@25757.4]
  wire  x286_rdrow_1_reset; // @[Math.scala 191:24:@25757.4]
  wire [31:0] x286_rdrow_1_io_a; // @[Math.scala 191:24:@25757.4]
  wire [31:0] x286_rdrow_1_io_b; // @[Math.scala 191:24:@25757.4]
  wire  x286_rdrow_1_io_flow; // @[Math.scala 191:24:@25757.4]
  wire [31:0] x286_rdrow_1_io_result; // @[Math.scala 191:24:@25757.4]
  wire  x287_1_clock; // @[Math.scala 366:24:@25769.4]
  wire  x287_1_reset; // @[Math.scala 366:24:@25769.4]
  wire [31:0] x287_1_io_a; // @[Math.scala 366:24:@25769.4]
  wire  x287_1_io_flow; // @[Math.scala 366:24:@25769.4]
  wire [31:0] x287_1_io_result; // @[Math.scala 366:24:@25769.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@25784.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@25784.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@25784.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@25784.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@25784.4]
  wire  x293_mul_1_clock; // @[Math.scala 262:24:@25821.4]
  wire  x293_mul_1_reset; // @[Math.scala 262:24:@25821.4]
  wire [31:0] x293_mul_1_io_a; // @[Math.scala 262:24:@25821.4]
  wire  x293_mul_1_io_flow; // @[Math.scala 262:24:@25821.4]
  wire [31:0] x293_mul_1_io_result; // @[Math.scala 262:24:@25821.4]
  wire  x294_sum_1_clock; // @[Math.scala 150:24:@25831.4]
  wire  x294_sum_1_reset; // @[Math.scala 150:24:@25831.4]
  wire [31:0] x294_sum_1_io_a; // @[Math.scala 150:24:@25831.4]
  wire [31:0] x294_sum_1_io_b; // @[Math.scala 150:24:@25831.4]
  wire  x294_sum_1_io_flow; // @[Math.scala 150:24:@25831.4]
  wire [31:0] x294_sum_1_io_result; // @[Math.scala 150:24:@25831.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@25841.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@25841.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@25841.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@25841.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@25841.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@25850.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@25850.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@25850.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@25850.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@25850.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@25859.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@25859.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@25859.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@25859.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@25859.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@25871.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@25871.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@25871.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@25871.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@25871.4]
  wire  x299_sum_1_clock; // @[Math.scala 150:24:@25898.4]
  wire  x299_sum_1_reset; // @[Math.scala 150:24:@25898.4]
  wire [31:0] x299_sum_1_io_a; // @[Math.scala 150:24:@25898.4]
  wire [31:0] x299_sum_1_io_b; // @[Math.scala 150:24:@25898.4]
  wire  x299_sum_1_io_flow; // @[Math.scala 150:24:@25898.4]
  wire [31:0] x299_sum_1_io_result; // @[Math.scala 150:24:@25898.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@25908.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@25908.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@25908.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@25908.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@25908.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@25917.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@25917.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@25917.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@25917.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@25917.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@25929.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@25929.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@25929.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@25929.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@25929.4]
  wire  x304_sum_1_clock; // @[Math.scala 150:24:@25956.4]
  wire  x304_sum_1_reset; // @[Math.scala 150:24:@25956.4]
  wire [31:0] x304_sum_1_io_a; // @[Math.scala 150:24:@25956.4]
  wire [31:0] x304_sum_1_io_b; // @[Math.scala 150:24:@25956.4]
  wire  x304_sum_1_io_flow; // @[Math.scala 150:24:@25956.4]
  wire [31:0] x304_sum_1_io_result; // @[Math.scala 150:24:@25956.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@25975.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@25975.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@25975.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@25975.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@25975.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@25987.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@25987.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@25987.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@25987.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@25987.4]
  wire  x312_x11_1_clock; // @[Math.scala 150:24:@26035.4]
  wire  x312_x11_1_reset; // @[Math.scala 150:24:@26035.4]
  wire [7:0] x312_x11_1_io_a; // @[Math.scala 150:24:@26035.4]
  wire [7:0] x312_x11_1_io_b; // @[Math.scala 150:24:@26035.4]
  wire  x312_x11_1_io_flow; // @[Math.scala 150:24:@26035.4]
  wire [7:0] x312_x11_1_io_result; // @[Math.scala 150:24:@26035.4]
  wire  x313_x12_1_clock; // @[Math.scala 150:24:@26045.4]
  wire  x313_x12_1_reset; // @[Math.scala 150:24:@26045.4]
  wire [7:0] x313_x12_1_io_a; // @[Math.scala 150:24:@26045.4]
  wire [7:0] x313_x12_1_io_b; // @[Math.scala 150:24:@26045.4]
  wire  x313_x12_1_io_flow; // @[Math.scala 150:24:@26045.4]
  wire [7:0] x313_x12_1_io_result; // @[Math.scala 150:24:@26045.4]
  wire  x314_x11_1_clock; // @[Math.scala 150:24:@26055.4]
  wire  x314_x11_1_reset; // @[Math.scala 150:24:@26055.4]
  wire [7:0] x314_x11_1_io_a; // @[Math.scala 150:24:@26055.4]
  wire [7:0] x314_x11_1_io_b; // @[Math.scala 150:24:@26055.4]
  wire  x314_x11_1_io_flow; // @[Math.scala 150:24:@26055.4]
  wire [7:0] x314_x11_1_io_result; // @[Math.scala 150:24:@26055.4]
  wire  x315_x12_1_clock; // @[Math.scala 150:24:@26065.4]
  wire  x315_x12_1_reset; // @[Math.scala 150:24:@26065.4]
  wire [7:0] x315_x12_1_io_a; // @[Math.scala 150:24:@26065.4]
  wire [7:0] x315_x12_1_io_b; // @[Math.scala 150:24:@26065.4]
  wire  x315_x12_1_io_flow; // @[Math.scala 150:24:@26065.4]
  wire [7:0] x315_x12_1_io_result; // @[Math.scala 150:24:@26065.4]
  wire [7:0] x316_x11_1_io_a; // @[Math.scala 150:24:@26075.4]
  wire [7:0] x316_x11_1_io_b; // @[Math.scala 150:24:@26075.4]
  wire [7:0] x316_x11_1_io_result; // @[Math.scala 150:24:@26075.4]
  wire [7:0] x317_x12_1_io_a; // @[Math.scala 150:24:@26085.4]
  wire [7:0] x317_x12_1_io_b; // @[Math.scala 150:24:@26085.4]
  wire [7:0] x317_x12_1_io_result; // @[Math.scala 150:24:@26085.4]
  wire [7:0] x318_x11_1_io_a; // @[Math.scala 150:24:@26095.4]
  wire [7:0] x318_x11_1_io_b; // @[Math.scala 150:24:@26095.4]
  wire [7:0] x318_x11_1_io_result; // @[Math.scala 150:24:@26095.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@26105.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@26105.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@26105.4]
  wire [7:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@26105.4]
  wire [7:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@26105.4]
  wire [7:0] x319_sum_1_io_a; // @[Math.scala 150:24:@26114.4]
  wire [7:0] x319_sum_1_io_b; // @[Math.scala 150:24:@26114.4]
  wire [7:0] x319_sum_1_io_result; // @[Math.scala 150:24:@26114.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@26128.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@26128.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@26128.4]
  wire [7:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@26128.4]
  wire [7:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@26128.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@26142.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@26142.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@26142.4]
  wire [7:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@26142.4]
  wire [7:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@26142.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@26151.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@26151.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@26151.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@26151.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@26151.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@26160.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@26160.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@26160.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@26160.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@26160.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@26169.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@26169.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@26169.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@26169.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@26169.4]
  wire  b216; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 62:18:@24006.4]
  wire  b217; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 63:18:@24007.4]
  wire  _T_206; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 68:30:@24076.4]
  wire  _T_207; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 68:37:@24077.4]
  wire  _T_211; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 70:76:@24082.4]
  wire  _T_212; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 70:62:@24083.4]
  wire  _T_214; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 70:101:@24084.4]
  wire [31:0] b214_number; // @[Math.scala 712:22:@23991.4 Math.scala 713:14:@23992.4]
  wire [31:0] _T_240; // @[Math.scala 499:52:@24107.4]
  wire  x223; // @[Math.scala 499:44:@24115.4]
  wire  x224; // @[Math.scala 499:44:@24122.4]
  wire  x225; // @[Math.scala 499:44:@24129.4]
  wire [31:0] _T_287; // @[Mux.scala 19:72:@24141.4]
  wire [31:0] _T_289; // @[Mux.scala 19:72:@24142.4]
  wire [31:0] _T_291; // @[Mux.scala 19:72:@24143.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@24145.4]
  wire [31:0] x226_number; // @[Mux.scala 19:72:@24146.4]
  wire [31:0] _T_305; // @[Math.scala 406:49:@24156.4]
  wire [31:0] _T_307; // @[Math.scala 406:56:@24158.4]
  wire [31:0] _T_308; // @[Math.scala 406:56:@24159.4]
  wire [31:0] b215_number; // @[Math.scala 712:22:@24003.4 Math.scala 713:14:@24004.4]
  wire  _T_313; // @[FixedPoint.scala 50:25:@24165.4]
  wire [15:0] _T_317; // @[Bitwise.scala 72:12:@24167.4]
  wire [15:0] _T_318; // @[FixedPoint.scala 18:52:@24168.4]
  wire [31:0] _T_327; // @[Math.scala 406:49:@24176.4]
  wire [31:0] _T_329; // @[Math.scala 406:56:@24178.4]
  wire [31:0] _T_330; // @[Math.scala 406:56:@24179.4]
  wire [31:0] x396_sum_number; // @[Math.scala 154:22:@24190.4 Math.scala 155:14:@24191.4]
  wire  _T_338; // @[FixedPoint.scala 50:25:@24195.4]
  wire [7:0] _T_342; // @[Bitwise.scala 72:12:@24197.4]
  wire [23:0] _T_343; // @[FixedPoint.scala 18:52:@24198.4]
  wire [31:0] _T_352; // @[Math.scala 406:49:@24206.4]
  wire [31:0] _T_354; // @[Math.scala 406:56:@24208.4]
  wire [31:0] _T_355; // @[Math.scala 406:56:@24209.4]
  wire [31:0] x399_sum_number; // @[Math.scala 154:22:@24220.4 Math.scala 155:14:@24221.4]
  wire  _T_363; // @[FixedPoint.scala 50:25:@24225.4]
  wire [3:0] _T_367; // @[Bitwise.scala 72:12:@24227.4]
  wire [27:0] _T_368; // @[FixedPoint.scala 18:52:@24228.4]
  wire [31:0] _T_377; // @[Math.scala 406:49:@24236.4]
  wire [31:0] _T_379; // @[Math.scala 406:56:@24238.4]
  wire [31:0] _T_380; // @[Math.scala 406:56:@24239.4]
  wire [31:0] x402_sum_number; // @[Math.scala 154:22:@24250.4 Math.scala 155:14:@24251.4]
  wire  _T_388; // @[FixedPoint.scala 50:25:@24255.4]
  wire [1:0] _T_392; // @[Bitwise.scala 72:12:@24257.4]
  wire [29:0] _T_393; // @[FixedPoint.scala 18:52:@24258.4]
  wire [31:0] _T_402; // @[Math.scala 406:49:@24266.4]
  wire [31:0] _T_404; // @[Math.scala 406:56:@24268.4]
  wire [31:0] _T_405; // @[Math.scala 406:56:@24269.4]
  wire [31:0] x405_sum_number; // @[Math.scala 154:22:@24280.4 Math.scala 155:14:@24281.4]
  wire  _T_413; // @[FixedPoint.scala 50:25:@24285.4]
  wire [1:0] _T_417; // @[Bitwise.scala 72:12:@24287.4]
  wire [29:0] _T_418; // @[FixedPoint.scala 18:52:@24288.4]
  wire [31:0] _T_429; // @[Math.scala 406:49:@24303.4]
  wire [31:0] _T_431; // @[Math.scala 406:56:@24305.4]
  wire [31:0] _T_432; // @[Math.scala 406:56:@24306.4]
  wire [31:0] _T_436; // @[package.scala 96:25:@24314.4]
  wire [31:0] x408_sum_number; // @[Math.scala 154:22:@24326.4 Math.scala 155:14:@24327.4]
  wire  _T_444; // @[FixedPoint.scala 50:25:@24331.4]
  wire [1:0] _T_448; // @[Bitwise.scala 72:12:@24333.4]
  wire [29:0] _T_449; // @[FixedPoint.scala 18:52:@24334.4]
  wire [31:0] _T_458; // @[Math.scala 406:49:@24342.4]
  wire [31:0] _T_460; // @[Math.scala 406:56:@24344.4]
  wire [31:0] _T_461; // @[Math.scala 406:56:@24345.4]
  wire [31:0] x411_sum_number; // @[Math.scala 154:22:@24356.4 Math.scala 155:14:@24357.4]
  wire [31:0] _T_471; // @[Math.scala 465:37:@24362.4]
  wire  x466_x412_D1; // @[package.scala 96:25:@24400.4 package.scala 96:25:@24401.4]
  wire [31:0] x467_x411_sum_D1_number; // @[package.scala 96:25:@24409.4 package.scala 96:25:@24410.4]
  wire [31:0] x414_sub_number; // @[Math.scala 195:22:@24382.4 Math.scala 196:14:@24383.4]
  wire  _T_503; // @[FixedPoint.scala 50:25:@24417.4]
  wire [1:0] _T_507; // @[Bitwise.scala 72:12:@24419.4]
  wire [29:0] _T_508; // @[FixedPoint.scala 18:52:@24420.4]
  wire  _T_546; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:101:@24510.4]
  wire  _T_550; // @[package.scala 96:25:@24518.4 package.scala 96:25:@24519.4]
  wire  _T_552; // @[implicits.scala 55:10:@24520.4]
  wire  _T_553; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:118:@24521.4]
  wire  _T_555; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:207:@24523.4]
  wire  _T_556; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:226:@24524.4]
  wire  x470_b216_D26; // @[package.scala 96:25:@24480.4 package.scala 96:25:@24481.4]
  wire  _T_557; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:252:@24525.4]
  wire  x469_b217_D26; // @[package.scala 96:25:@24471.4 package.scala 96:25:@24472.4]
  wire [31:0] x474_b214_D28_number; // @[package.scala 96:25:@24539.4 package.scala 96:25:@24540.4]
  wire [31:0] _T_576; // @[Math.scala 465:37:@24559.4]
  wire [31:0] x475_b215_D28_number; // @[package.scala 96:25:@24576.4 package.scala 96:25:@24577.4]
  wire [31:0] _T_589; // @[Math.scala 465:37:@24582.4]
  wire  x237; // @[package.scala 96:25:@24567.4 package.scala 96:25:@24568.4]
  wire  x238; // @[package.scala 96:25:@24590.4 package.scala 96:25:@24591.4]
  wire  x239; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 186:24:@24594.4]
  wire [31:0] x236_number; // @[Math.scala 370:22:@24553.4 Math.scala 371:14:@24554.4]
  wire [31:0] _T_605; // @[Math.scala 406:49:@24603.4]
  wire [31:0] _T_607; // @[Math.scala 406:56:@24605.4]
  wire [31:0] _T_608; // @[Math.scala 406:56:@24606.4]
  wire  _T_613; // @[FixedPoint.scala 50:25:@24612.4]
  wire [1:0] _T_617; // @[Bitwise.scala 72:12:@24614.4]
  wire [29:0] _T_618; // @[FixedPoint.scala 18:52:@24615.4]
  wire  _T_662; // @[package.scala 96:25:@24713.4 package.scala 96:25:@24714.4]
  wire  _T_664; // @[implicits.scala 55:10:@24715.4]
  wire  _T_665; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 215:194:@24716.4]
  wire  x481_x240_D26; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  wire  _T_666; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 215:283:@24717.4]
  wire  x479_b216_D55; // @[package.scala 96:25:@24674.4 package.scala 96:25:@24675.4]
  wire  _T_667; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 215:291:@24718.4]
  wire  x477_b217_D55; // @[package.scala 96:25:@24656.4 package.scala 96:25:@24657.4]
  wire [31:0] x247_rdcol_number; // @[Math.scala 195:22:@24737.4 Math.scala 196:14:@24738.4]
  wire [31:0] _T_682; // @[Math.scala 465:37:@24743.4]
  wire  x483_x237_D1; // @[package.scala 96:25:@24760.4 package.scala 96:25:@24761.4]
  wire  x248; // @[package.scala 96:25:@24751.4 package.scala 96:25:@24752.4]
  wire  x249; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 225:24:@24764.4]
  wire  _T_697; // @[FixedPoint.scala 50:25:@24771.4]
  wire [15:0] _T_701; // @[Bitwise.scala 72:12:@24773.4]
  wire [15:0] _T_702; // @[FixedPoint.scala 18:52:@24774.4]
  wire [31:0] _T_713; // @[Math.scala 406:56:@24784.4]
  wire [31:0] _T_714; // @[Math.scala 406:56:@24785.4]
  wire [31:0] x420_sum_number; // @[Math.scala 154:22:@24796.4 Math.scala 155:14:@24797.4]
  wire  _T_722; // @[FixedPoint.scala 50:25:@24801.4]
  wire [7:0] _T_726; // @[Bitwise.scala 72:12:@24803.4]
  wire [23:0] _T_727; // @[FixedPoint.scala 18:52:@24804.4]
  wire [31:0] _T_738; // @[Math.scala 406:49:@24819.4]
  wire [31:0] _T_740; // @[Math.scala 406:56:@24821.4]
  wire [31:0] _T_741; // @[Math.scala 406:56:@24822.4]
  wire [31:0] _T_745; // @[package.scala 96:25:@24830.4]
  wire [31:0] x423_sum_number; // @[Math.scala 154:22:@24842.4 Math.scala 155:14:@24843.4]
  wire  _T_753; // @[FixedPoint.scala 50:25:@24847.4]
  wire [3:0] _T_757; // @[Bitwise.scala 72:12:@24849.4]
  wire [27:0] _T_758; // @[FixedPoint.scala 18:52:@24850.4]
  wire [31:0] _T_767; // @[Math.scala 406:49:@24858.4]
  wire [31:0] _T_769; // @[Math.scala 406:56:@24860.4]
  wire [31:0] _T_770; // @[Math.scala 406:56:@24861.4]
  wire [31:0] x426_sum_number; // @[Math.scala 154:22:@24872.4 Math.scala 155:14:@24873.4]
  wire  _T_778; // @[FixedPoint.scala 50:25:@24877.4]
  wire [1:0] _T_782; // @[Bitwise.scala 72:12:@24879.4]
  wire [29:0] _T_783; // @[FixedPoint.scala 18:52:@24880.4]
  wire [31:0] _T_792; // @[Math.scala 406:49:@24888.4]
  wire [31:0] _T_794; // @[Math.scala 406:56:@24890.4]
  wire [31:0] _T_795; // @[Math.scala 406:56:@24891.4]
  wire [31:0] x429_sum_number; // @[Math.scala 154:22:@24902.4 Math.scala 155:14:@24903.4]
  wire  _T_803; // @[FixedPoint.scala 50:25:@24907.4]
  wire [1:0] _T_807; // @[Bitwise.scala 72:12:@24909.4]
  wire [29:0] _T_808; // @[FixedPoint.scala 18:52:@24910.4]
  wire [31:0] _T_817; // @[Math.scala 406:49:@24918.4]
  wire [31:0] _T_819; // @[Math.scala 406:56:@24920.4]
  wire [31:0] _T_820; // @[Math.scala 406:56:@24921.4]
  wire [31:0] x432_sum_number; // @[Math.scala 154:22:@24932.4 Math.scala 155:14:@24933.4]
  wire  _T_828; // @[FixedPoint.scala 50:25:@24937.4]
  wire [1:0] _T_832; // @[Bitwise.scala 72:12:@24939.4]
  wire [29:0] _T_833; // @[FixedPoint.scala 18:52:@24940.4]
  wire [31:0] _T_842; // @[Math.scala 406:49:@24948.4]
  wire [31:0] _T_844; // @[Math.scala 406:56:@24950.4]
  wire [31:0] _T_845; // @[Math.scala 406:56:@24951.4]
  wire [31:0] x435_sum_number; // @[Math.scala 154:22:@24962.4 Math.scala 155:14:@24963.4]
  wire [31:0] _T_855; // @[Math.scala 465:37:@24968.4]
  wire  x436; // @[package.scala 96:25:@24976.4 package.scala 96:25:@24977.4]
  wire [31:0] x484_x435_sum_D1_number; // @[package.scala 96:25:@25011.4 package.scala 96:25:@25012.4]
  wire [31:0] x438_sub_number; // @[Math.scala 195:22:@25002.4 Math.scala 196:14:@25003.4]
  wire  _T_917; // @[package.scala 96:25:@25086.4 package.scala 96:25:@25087.4]
  wire  _T_919; // @[implicits.scala 55:10:@25088.4]
  wire  _T_920; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:194:@25089.4]
  wire  x488_x250_D25; // @[package.scala 96:25:@25074.4 package.scala 96:25:@25075.4]
  wire  _T_921; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:283:@25090.4]
  wire  _T_922; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:291:@25091.4]
  wire [31:0] x256_rdcol_number; // @[Math.scala 195:22:@25110.4 Math.scala 196:14:@25111.4]
  wire [31:0] _T_937; // @[Math.scala 465:37:@25116.4]
  wire  x257; // @[package.scala 96:25:@25124.4 package.scala 96:25:@25125.4]
  wire  x258; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 306:59:@25128.4]
  wire  _T_949; // @[FixedPoint.scala 50:25:@25135.4]
  wire [15:0] _T_953; // @[Bitwise.scala 72:12:@25137.4]
  wire [15:0] _T_954; // @[FixedPoint.scala 18:52:@25138.4]
  wire [31:0] _T_965; // @[Math.scala 406:56:@25148.4]
  wire [31:0] _T_966; // @[Math.scala 406:56:@25149.4]
  wire [31:0] x442_sum_number; // @[Math.scala 154:22:@25160.4 Math.scala 155:14:@25161.4]
  wire  _T_974; // @[FixedPoint.scala 50:25:@25165.4]
  wire [7:0] _T_978; // @[Bitwise.scala 72:12:@25167.4]
  wire [23:0] _T_979; // @[FixedPoint.scala 18:52:@25168.4]
  wire [31:0] _T_990; // @[Math.scala 406:49:@25183.4]
  wire [31:0] _T_992; // @[Math.scala 406:56:@25185.4]
  wire [31:0] _T_993; // @[Math.scala 406:56:@25186.4]
  wire [31:0] _T_997; // @[package.scala 96:25:@25194.4]
  wire [31:0] x445_sum_number; // @[Math.scala 154:22:@25206.4 Math.scala 155:14:@25207.4]
  wire  _T_1005; // @[FixedPoint.scala 50:25:@25211.4]
  wire [3:0] _T_1009; // @[Bitwise.scala 72:12:@25213.4]
  wire [27:0] _T_1010; // @[FixedPoint.scala 18:52:@25214.4]
  wire [31:0] _T_1019; // @[Math.scala 406:49:@25222.4]
  wire [31:0] _T_1021; // @[Math.scala 406:56:@25224.4]
  wire [31:0] _T_1022; // @[Math.scala 406:56:@25225.4]
  wire [31:0] x448_sum_number; // @[Math.scala 154:22:@25236.4 Math.scala 155:14:@25237.4]
  wire  _T_1030; // @[FixedPoint.scala 50:25:@25241.4]
  wire [1:0] _T_1034; // @[Bitwise.scala 72:12:@25243.4]
  wire [29:0] _T_1035; // @[FixedPoint.scala 18:52:@25244.4]
  wire [31:0] _T_1044; // @[Math.scala 406:49:@25252.4]
  wire [31:0] _T_1046; // @[Math.scala 406:56:@25254.4]
  wire [31:0] _T_1047; // @[Math.scala 406:56:@25255.4]
  wire [31:0] x451_sum_number; // @[Math.scala 154:22:@25266.4 Math.scala 155:14:@25267.4]
  wire  _T_1055; // @[FixedPoint.scala 50:25:@25271.4]
  wire [1:0] _T_1059; // @[Bitwise.scala 72:12:@25273.4]
  wire [29:0] _T_1060; // @[FixedPoint.scala 18:52:@25274.4]
  wire [31:0] _T_1069; // @[Math.scala 406:49:@25282.4]
  wire [31:0] _T_1071; // @[Math.scala 406:56:@25284.4]
  wire [31:0] _T_1072; // @[Math.scala 406:56:@25285.4]
  wire [31:0] x454_sum_number; // @[Math.scala 154:22:@25296.4 Math.scala 155:14:@25297.4]
  wire  _T_1080; // @[FixedPoint.scala 50:25:@25301.4]
  wire [1:0] _T_1084; // @[Bitwise.scala 72:12:@25303.4]
  wire [29:0] _T_1085; // @[FixedPoint.scala 18:52:@25304.4]
  wire [31:0] _T_1094; // @[Math.scala 406:49:@25312.4]
  wire [31:0] _T_1096; // @[Math.scala 406:56:@25314.4]
  wire [31:0] _T_1097; // @[Math.scala 406:56:@25315.4]
  wire [31:0] x457_sum_number; // @[Math.scala 154:22:@25326.4 Math.scala 155:14:@25327.4]
  wire [31:0] _T_1107; // @[Math.scala 465:37:@25332.4]
  wire  x458; // @[package.scala 96:25:@25340.4 package.scala 96:25:@25341.4]
  wire [31:0] x489_x457_sum_D1_number; // @[package.scala 96:25:@25375.4 package.scala 96:25:@25376.4]
  wire [31:0] x460_sub_number; // @[Math.scala 195:22:@25366.4 Math.scala 196:14:@25367.4]
  wire  _T_1167; // @[package.scala 96:25:@25448.4 package.scala 96:25:@25449.4]
  wire  _T_1169; // @[implicits.scala 55:10:@25450.4]
  wire  _T_1170; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 371:194:@25451.4]
  wire  x492_x259_D25; // @[package.scala 96:25:@25427.4 package.scala 96:25:@25428.4]
  wire  _T_1171; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 371:283:@25452.4]
  wire  _T_1172; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 371:291:@25453.4]
  wire [31:0] x265_rdrow_number; // @[Math.scala 195:22:@25472.4 Math.scala 196:14:@25473.4]
  wire [31:0] _T_1194; // @[Math.scala 465:37:@25490.4]
  wire  x267; // @[package.scala 96:25:@25498.4 package.scala 96:25:@25499.4]
  wire  x494_x238_D1; // @[package.scala 96:25:@25507.4 package.scala 96:25:@25508.4]
  wire  x268; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 383:24:@25511.4]
  wire [31:0] x266_number; // @[Math.scala 370:22:@25484.4 Math.scala 371:14:@25485.4]
  wire [31:0] _T_1213; // @[Math.scala 406:49:@25520.4]
  wire [31:0] _T_1215; // @[Math.scala 406:56:@25522.4]
  wire [31:0] _T_1216; // @[Math.scala 406:56:@25523.4]
  wire  _T_1221; // @[FixedPoint.scala 50:25:@25529.4]
  wire [1:0] _T_1225; // @[Bitwise.scala 72:12:@25531.4]
  wire [29:0] _T_1226; // @[FixedPoint.scala 18:52:@25532.4]
  wire  _T_1263; // @[package.scala 96:25:@25605.4 package.scala 96:25:@25606.4]
  wire  _T_1265; // @[implicits.scala 55:10:@25607.4]
  wire  _T_1266; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:194:@25608.4]
  wire  x496_x269_D25; // @[package.scala 96:25:@25575.4 package.scala 96:25:@25576.4]
  wire  _T_1267; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:283:@25609.4]
  wire  _T_1268; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:291:@25610.4]
  wire  x276; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 418:59:@25621.4]
  wire  _T_1298; // @[package.scala 96:25:@25672.4 package.scala 96:25:@25673.4]
  wire  _T_1300; // @[implicits.scala 55:10:@25674.4]
  wire  _T_1301; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:194:@25675.4]
  wire  x501_x277_D25; // @[package.scala 96:25:@25660.4 package.scala 96:25:@25661.4]
  wire  _T_1302; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:283:@25676.4]
  wire  _T_1303; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:291:@25677.4]
  wire  x281; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 437:59:@25688.4]
  wire  _T_1333; // @[package.scala 96:25:@25739.4 package.scala 96:25:@25740.4]
  wire  _T_1335; // @[implicits.scala 55:10:@25741.4]
  wire  _T_1336; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:194:@25742.4]
  wire  x503_x282_D25; // @[package.scala 96:25:@25718.4 package.scala 96:25:@25719.4]
  wire  _T_1337; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:283:@25743.4]
  wire  _T_1338; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:291:@25744.4]
  wire [31:0] x286_rdrow_number; // @[Math.scala 195:22:@25763.4 Math.scala 196:14:@25764.4]
  wire [31:0] _T_1360; // @[Math.scala 465:37:@25781.4]
  wire  x288; // @[package.scala 96:25:@25789.4 package.scala 96:25:@25790.4]
  wire  x289; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 462:24:@25793.4]
  wire [31:0] x287_number; // @[Math.scala 370:22:@25775.4 Math.scala 371:14:@25776.4]
  wire [31:0] _T_1376; // @[Math.scala 406:49:@25802.4]
  wire [31:0] _T_1378; // @[Math.scala 406:56:@25804.4]
  wire [31:0] _T_1379; // @[Math.scala 406:56:@25805.4]
  wire  _T_1384; // @[FixedPoint.scala 50:25:@25811.4]
  wire [1:0] _T_1388; // @[Bitwise.scala 72:12:@25813.4]
  wire [29:0] _T_1389; // @[FixedPoint.scala 18:52:@25814.4]
  wire  _T_1421; // @[package.scala 96:25:@25876.4 package.scala 96:25:@25877.4]
  wire  _T_1423; // @[implicits.scala 55:10:@25878.4]
  wire  _T_1424; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 483:194:@25879.4]
  wire  x506_x290_D25; // @[package.scala 96:25:@25855.4 package.scala 96:25:@25856.4]
  wire  _T_1425; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 483:283:@25880.4]
  wire  _T_1426; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 483:291:@25881.4]
  wire  x297; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 487:24:@25892.4]
  wire  _T_1453; // @[package.scala 96:25:@25934.4 package.scala 96:25:@25935.4]
  wire  _T_1455; // @[implicits.scala 55:10:@25936.4]
  wire  _T_1456; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:194:@25937.4]
  wire  x508_x298_D25; // @[package.scala 96:25:@25913.4 package.scala 96:25:@25914.4]
  wire  _T_1457; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:283:@25938.4]
  wire  _T_1458; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:291:@25939.4]
  wire  x302; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 504:24:@25950.4]
  wire  _T_1485; // @[package.scala 96:25:@25992.4 package.scala 96:25:@25993.4]
  wire  _T_1487; // @[implicits.scala 55:10:@25994.4]
  wire  _T_1488; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 523:194:@25995.4]
  wire  x510_x303_D25; // @[package.scala 96:25:@25971.4 package.scala 96:25:@25972.4]
  wire  _T_1489; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 523:283:@25996.4]
  wire  _T_1490; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 523:326:@25997.4]
  wire [7:0] x254_rd_0_number; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 294:29:@25077.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:408:@25098.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@26011.4]
  wire [8:0] _T_1498; // @[Math.scala 450:32:@26011.4]
  wire [7:0] x274_rd_0_number; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 410:29:@25596.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:408:@25617.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@26016.4]
  wire [8:0] _T_1502; // @[Math.scala 450:32:@26016.4]
  wire [7:0] x279_rd_0_number; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 429:29:@25663.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:408:@25684.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@26021.4]
  wire [9:0] _T_1506; // @[Math.scala 450:32:@26021.4]
  wire [7:0] x284_rd_0_number; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 448:29:@25730.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:408:@25751.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@26026.4]
  wire [8:0] _T_1510; // @[Math.scala 450:32:@26026.4]
  wire [7:0] x300_rd_0_number; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 496:29:@25925.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:408:@25946.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@26031.4]
  wire [8:0] _T_1514; // @[Math.scala 450:32:@26031.4]
  wire [7:0] x319_sum_number; // @[Math.scala 154:22:@26120.4 Math.scala 155:14:@26121.4]
  wire [3:0] _T_1550; // @[FixedPoint.scala 18:52:@26126.4]
  wire  _T_1573; // @[package.scala 96:25:@26174.4 package.scala 96:25:@26175.4]
  wire  _T_1575; // @[implicits.scala 55:10:@26176.4]
  wire  x513_b216_D62; // @[package.scala 96:25:@26156.4 package.scala 96:25:@26157.4]
  wire  _T_1576; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 567:117:@26177.4]
  wire  x514_b217_D62; // @[package.scala 96:25:@26165.4 package.scala 96:25:@26166.4]
  wire  _T_1577; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 567:123:@26178.4]
  wire [31:0] x416_number; // @[Math.scala 712:22:@24462.4 Math.scala 713:14:@24463.4]
  wire [31:0] x471_x393_D26_number; // @[package.scala 96:25:@24489.4 package.scala 96:25:@24490.4]
  wire [31:0] x472_x415_D18_number; // @[package.scala 96:25:@24498.4 package.scala 96:25:@24499.4]
  wire [31:0] x478_x417_D11_number; // @[package.scala 96:25:@24665.4 package.scala 96:25:@24666.4]
  wire [31:0] x480_x244_sum_D4_number; // @[package.scala 96:25:@24683.4 package.scala 96:25:@24684.4]
  wire [31:0] x482_x415_D47_number; // @[package.scala 96:25:@24701.4 package.scala 96:25:@24702.4]
  wire [31:0] x486_x253_sum_D4_number; // @[package.scala 96:25:@25056.4 package.scala 96:25:@25057.4]
  wire [31:0] x487_x439_D18_number; // @[package.scala 96:25:@25065.4 package.scala 96:25:@25066.4]
  wire [31:0] x491_x461_D18_number; // @[package.scala 96:25:@25418.4 package.scala 96:25:@25419.4]
  wire [31:0] x493_x262_sum_D4_number; // @[package.scala 96:25:@25436.4 package.scala 96:25:@25437.4]
  wire [31:0] x497_x462_D10_number; // @[package.scala 96:25:@25584.4 package.scala 96:25:@25585.4]
  wire [31:0] x498_x273_sum_D3_number; // @[package.scala 96:25:@25593.4 package.scala 96:25:@25594.4]
  wire [31:0] x500_x278_sum_D3_number; // @[package.scala 96:25:@25651.4 package.scala 96:25:@25652.4]
  wire [31:0] x504_x283_sum_D3_number; // @[package.scala 96:25:@25727.4 package.scala 96:25:@25728.4]
  wire [31:0] x505_x463_D10_number; // @[package.scala 96:25:@25846.4 package.scala 96:25:@25847.4]
  wire [31:0] x507_x294_sum_D3_number; // @[package.scala 96:25:@25864.4 package.scala 96:25:@25865.4]
  wire [31:0] x509_x299_sum_D3_number; // @[package.scala 96:25:@25922.4 package.scala 96:25:@25923.4]
  wire [31:0] x511_x304_sum_D3_number; // @[package.scala 96:25:@25980.4 package.scala 96:25:@25981.4]
  _ _ ( // @[Math.scala 709:24:@23986.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@23998.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x218_lb_0 x218_lb_0 ( // @[m_x218_lb_0.scala 35:17:@24008.4]
    .clock(x218_lb_0_clock),
    .reset(x218_lb_0_reset),
    .io_rPort_8_banks_1(x218_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x218_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x218_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x218_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x218_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x218_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x218_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x218_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x218_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x218_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x218_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x218_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x218_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x218_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x218_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x218_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x218_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x218_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x218_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x218_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x218_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x218_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x218_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x218_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x218_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x218_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x218_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x218_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x218_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x218_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x218_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x218_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x218_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x218_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x218_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x218_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x218_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x218_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x218_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x218_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x218_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x218_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x218_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x218_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x218_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x218_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x218_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x218_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x218_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x218_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x218_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x218_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x218_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x218_lb_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x218_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x218_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x218_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x218_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x218_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_140 RetimeWrapper ( // @[package.scala 93:22:@24088.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x396_sum x396_sum_1 ( // @[Math.scala 150:24:@24184.4]
    .clock(x396_sum_1_clock),
    .reset(x396_sum_1_reset),
    .io_a(x396_sum_1_io_a),
    .io_b(x396_sum_1_io_b),
    .io_flow(x396_sum_1_io_flow),
    .io_result(x396_sum_1_io_result)
  );
  x396_sum x399_sum_1 ( // @[Math.scala 150:24:@24214.4]
    .clock(x399_sum_1_clock),
    .reset(x399_sum_1_reset),
    .io_a(x399_sum_1_io_a),
    .io_b(x399_sum_1_io_b),
    .io_flow(x399_sum_1_io_flow),
    .io_result(x399_sum_1_io_result)
  );
  x396_sum x402_sum_1 ( // @[Math.scala 150:24:@24244.4]
    .clock(x402_sum_1_clock),
    .reset(x402_sum_1_reset),
    .io_a(x402_sum_1_io_a),
    .io_b(x402_sum_1_io_b),
    .io_flow(x402_sum_1_io_flow),
    .io_result(x402_sum_1_io_result)
  );
  x396_sum x405_sum_1 ( // @[Math.scala 150:24:@24274.4]
    .clock(x405_sum_1_clock),
    .reset(x405_sum_1_reset),
    .io_a(x405_sum_1_io_a),
    .io_b(x405_sum_1_io_b),
    .io_flow(x405_sum_1_io_flow),
    .io_result(x405_sum_1_io_result)
  );
  RetimeWrapper_141 RetimeWrapper_1 ( // @[package.scala 93:22:@24290.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_141 RetimeWrapper_2 ( // @[package.scala 93:22:@24307.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x396_sum x408_sum_1 ( // @[Math.scala 150:24:@24320.4]
    .clock(x408_sum_1_clock),
    .reset(x408_sum_1_reset),
    .io_a(x408_sum_1_io_a),
    .io_b(x408_sum_1_io_b),
    .io_flow(x408_sum_1_io_flow),
    .io_result(x408_sum_1_io_result)
  );
  x396_sum x411_sum_1 ( // @[Math.scala 150:24:@24350.4]
    .clock(x411_sum_1_clock),
    .reset(x411_sum_1_reset),
    .io_a(x411_sum_1_io_a),
    .io_b(x411_sum_1_io_b),
    .io_flow(x411_sum_1_io_flow),
    .io_result(x411_sum_1_io_result)
  );
  x414_sub x414_sub_1 ( // @[Math.scala 191:24:@24376.4]
    .clock(x414_sub_1_clock),
    .reset(x414_sub_1_reset),
    .io_a(x414_sub_1_io_a),
    .io_b(x414_sub_1_io_b),
    .io_flow(x414_sub_1_io_flow),
    .io_result(x414_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@24386.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@24395.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_141 RetimeWrapper_5 ( // @[package.scala 93:22:@24404.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x232_div x232_div_1 ( // @[Math.scala 327:24:@24427.4]
    .clock(x232_div_1_clock),
    .reset(x232_div_1_reset),
    .io_a(x232_div_1_io_a),
    .io_flow(x232_div_1_io_flow),
    .io_result(x232_div_1_io_result)
  );
  RetimeWrapper_153 RetimeWrapper_6 ( // @[package.scala 93:22:@24437.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x416 x416_1 ( // @[Math.scala 849:24:@24448.4]
    .clock(x416_1_clock),
    .reset(x416_1_reset),
    .io_m0(x416_1_io_m0),
    .io_add(x416_1_io_add),
    .io_flow(x416_1_io_flow),
    .io_result(x416_1_io_result)
  );
  _ cast_x416 ( // @[Math.scala 709:24:@24457.4]
    .io_b(cast_x416_io_b),
    .io_result(cast_x416_io_result)
  );
  RetimeWrapper_159 RetimeWrapper_7 ( // @[package.scala 93:22:@24466.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_159 RetimeWrapper_8 ( // @[package.scala 93:22:@24475.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_161 RetimeWrapper_9 ( // @[package.scala 93:22:@24484.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_162 RetimeWrapper_10 ( // @[package.scala 93:22:@24493.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_163 RetimeWrapper_11 ( // @[package.scala 93:22:@24502.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_159 RetimeWrapper_12 ( // @[package.scala 93:22:@24513.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_13 ( // @[package.scala 93:22:@24534.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x236 x236_1 ( // @[Math.scala 366:24:@24547.4]
    .clock(x236_1_clock),
    .reset(x236_1_reset),
    .io_a(x236_1_io_a),
    .io_flow(x236_1_io_flow),
    .io_result(x236_1_io_result)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@24562.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_15 ( // @[package.scala 93:22:@24571.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@24585.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  fmamul_x416 x243_mul_1 ( // @[Math.scala 262:24:@24622.4]
    .clock(x243_mul_1_clock),
    .reset(x243_mul_1_reset),
    .io_a(x243_mul_1_io_a),
    .io_flow(x243_mul_1_io_flow),
    .io_result(x243_mul_1_io_result)
  );
  RetimeWrapper_173 RetimeWrapper_17 ( // @[package.scala 93:22:@24632.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x396_sum x244_sum_1 ( // @[Math.scala 150:24:@24641.4]
    .clock(x244_sum_1_clock),
    .reset(x244_sum_1_reset),
    .io_a(x244_sum_1_io_a),
    .io_b(x244_sum_1_io_b),
    .io_flow(x244_sum_1_io_flow),
    .io_result(x244_sum_1_io_result)
  );
  RetimeWrapper_175 RetimeWrapper_18 ( // @[package.scala 93:22:@24651.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_176 RetimeWrapper_19 ( // @[package.scala 93:22:@24660.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_20 ( // @[package.scala 93:22:@24669.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_178 RetimeWrapper_21 ( // @[package.scala 93:22:@24678.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_159 RetimeWrapper_22 ( // @[package.scala 93:22:@24687.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_180 RetimeWrapper_23 ( // @[package.scala 93:22:@24696.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_24 ( // @[package.scala 93:22:@24708.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x414_sub x247_rdcol_1 ( // @[Math.scala 191:24:@24731.4]
    .clock(x247_rdcol_1_clock),
    .reset(x247_rdcol_1_reset),
    .io_a(x247_rdcol_1_io_a),
    .io_b(x247_rdcol_1_io_b),
    .io_flow(x247_rdcol_1_io_flow),
    .io_result(x247_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@24746.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@24755.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  x396_sum x420_sum_1 ( // @[Math.scala 150:24:@24790.4]
    .clock(x420_sum_1_clock),
    .reset(x420_sum_1_reset),
    .io_a(x420_sum_1_io_a),
    .io_b(x420_sum_1_io_b),
    .io_flow(x420_sum_1_io_flow),
    .io_result(x420_sum_1_io_result)
  );
  RetimeWrapper_141 RetimeWrapper_27 ( // @[package.scala 93:22:@24806.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_141 RetimeWrapper_28 ( // @[package.scala 93:22:@24823.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x396_sum x423_sum_1 ( // @[Math.scala 150:24:@24836.4]
    .clock(x423_sum_1_clock),
    .reset(x423_sum_1_reset),
    .io_a(x423_sum_1_io_a),
    .io_b(x423_sum_1_io_b),
    .io_flow(x423_sum_1_io_flow),
    .io_result(x423_sum_1_io_result)
  );
  x396_sum x426_sum_1 ( // @[Math.scala 150:24:@24866.4]
    .clock(x426_sum_1_clock),
    .reset(x426_sum_1_reset),
    .io_a(x426_sum_1_io_a),
    .io_b(x426_sum_1_io_b),
    .io_flow(x426_sum_1_io_flow),
    .io_result(x426_sum_1_io_result)
  );
  x396_sum x429_sum_1 ( // @[Math.scala 150:24:@24896.4]
    .clock(x429_sum_1_clock),
    .reset(x429_sum_1_reset),
    .io_a(x429_sum_1_io_a),
    .io_b(x429_sum_1_io_b),
    .io_flow(x429_sum_1_io_flow),
    .io_result(x429_sum_1_io_result)
  );
  x396_sum x432_sum_1 ( // @[Math.scala 150:24:@24926.4]
    .clock(x432_sum_1_clock),
    .reset(x432_sum_1_reset),
    .io_a(x432_sum_1_io_a),
    .io_b(x432_sum_1_io_b),
    .io_flow(x432_sum_1_io_flow),
    .io_result(x432_sum_1_io_result)
  );
  x396_sum x435_sum_1 ( // @[Math.scala 150:24:@24956.4]
    .clock(x435_sum_1_clock),
    .reset(x435_sum_1_reset),
    .io_a(x435_sum_1_io_a),
    .io_b(x435_sum_1_io_b),
    .io_flow(x435_sum_1_io_flow),
    .io_result(x435_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@24971.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper RetimeWrapper_30 ( // @[package.scala 93:22:@24985.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x414_sub x438_sub_1 ( // @[Math.scala 191:24:@24996.4]
    .clock(x438_sub_1_clock),
    .reset(x438_sub_1_reset),
    .io_a(x438_sub_1_io_a),
    .io_b(x438_sub_1_io_b),
    .io_flow(x438_sub_1_io_flow),
    .io_result(x438_sub_1_io_result)
  );
  RetimeWrapper_141 RetimeWrapper_31 ( // @[package.scala 93:22:@25006.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x232_div x252_div_1 ( // @[Math.scala 327:24:@25020.4]
    .clock(x252_div_1_clock),
    .reset(x252_div_1_reset),
    .io_a(x252_div_1_io_a),
    .io_flow(x252_div_1_io_flow),
    .io_result(x252_div_1_io_result)
  );
  RetimeWrapper_141 RetimeWrapper_32 ( // @[package.scala 93:22:@25030.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x396_sum x253_sum_1 ( // @[Math.scala 150:24:@25041.4]
    .clock(x253_sum_1_clock),
    .reset(x253_sum_1_reset),
    .io_a(x253_sum_1_io_a),
    .io_b(x253_sum_1_io_b),
    .io_flow(x253_sum_1_io_flow),
    .io_result(x253_sum_1_io_result)
  );
  RetimeWrapper_178 RetimeWrapper_33 ( // @[package.scala 93:22:@25051.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_162 RetimeWrapper_34 ( // @[package.scala 93:22:@25060.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_202 RetimeWrapper_35 ( // @[package.scala 93:22:@25069.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_36 ( // @[package.scala 93:22:@25081.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x414_sub x256_rdcol_1 ( // @[Math.scala 191:24:@25104.4]
    .clock(x256_rdcol_1_clock),
    .reset(x256_rdcol_1_reset),
    .io_a(x256_rdcol_1_io_a),
    .io_b(x256_rdcol_1_io_b),
    .io_flow(x256_rdcol_1_io_flow),
    .io_result(x256_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_37 ( // @[package.scala 93:22:@25119.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x396_sum x442_sum_1 ( // @[Math.scala 150:24:@25154.4]
    .clock(x442_sum_1_clock),
    .reset(x442_sum_1_reset),
    .io_a(x442_sum_1_io_a),
    .io_b(x442_sum_1_io_b),
    .io_flow(x442_sum_1_io_flow),
    .io_result(x442_sum_1_io_result)
  );
  RetimeWrapper_141 RetimeWrapper_38 ( // @[package.scala 93:22:@25170.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_141 RetimeWrapper_39 ( // @[package.scala 93:22:@25187.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x396_sum x445_sum_1 ( // @[Math.scala 150:24:@25200.4]
    .clock(x445_sum_1_clock),
    .reset(x445_sum_1_reset),
    .io_a(x445_sum_1_io_a),
    .io_b(x445_sum_1_io_b),
    .io_flow(x445_sum_1_io_flow),
    .io_result(x445_sum_1_io_result)
  );
  x396_sum x448_sum_1 ( // @[Math.scala 150:24:@25230.4]
    .clock(x448_sum_1_clock),
    .reset(x448_sum_1_reset),
    .io_a(x448_sum_1_io_a),
    .io_b(x448_sum_1_io_b),
    .io_flow(x448_sum_1_io_flow),
    .io_result(x448_sum_1_io_result)
  );
  x396_sum x451_sum_1 ( // @[Math.scala 150:24:@25260.4]
    .clock(x451_sum_1_clock),
    .reset(x451_sum_1_reset),
    .io_a(x451_sum_1_io_a),
    .io_b(x451_sum_1_io_b),
    .io_flow(x451_sum_1_io_flow),
    .io_result(x451_sum_1_io_result)
  );
  x396_sum x454_sum_1 ( // @[Math.scala 150:24:@25290.4]
    .clock(x454_sum_1_clock),
    .reset(x454_sum_1_reset),
    .io_a(x454_sum_1_io_a),
    .io_b(x454_sum_1_io_b),
    .io_flow(x454_sum_1_io_flow),
    .io_result(x454_sum_1_io_result)
  );
  x396_sum x457_sum_1 ( // @[Math.scala 150:24:@25320.4]
    .clock(x457_sum_1_clock),
    .reset(x457_sum_1_reset),
    .io_a(x457_sum_1_io_a),
    .io_b(x457_sum_1_io_b),
    .io_flow(x457_sum_1_io_flow),
    .io_result(x457_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_40 ( // @[package.scala 93:22:@25335.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@25349.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  x414_sub x460_sub_1 ( // @[Math.scala 191:24:@25360.4]
    .clock(x460_sub_1_clock),
    .reset(x460_sub_1_reset),
    .io_a(x460_sub_1_io_a),
    .io_b(x460_sub_1_io_b),
    .io_flow(x460_sub_1_io_flow),
    .io_result(x460_sub_1_io_result)
  );
  RetimeWrapper_141 RetimeWrapper_42 ( // @[package.scala 93:22:@25370.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  x232_div x261_div_1 ( // @[Math.scala 327:24:@25384.4]
    .clock(x261_div_1_clock),
    .reset(x261_div_1_reset),
    .io_a(x261_div_1_io_a),
    .io_flow(x261_div_1_io_flow),
    .io_result(x261_div_1_io_result)
  );
  RetimeWrapper_141 RetimeWrapper_43 ( // @[package.scala 93:22:@25394.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x396_sum x262_sum_1 ( // @[Math.scala 150:24:@25403.4]
    .clock(x262_sum_1_clock),
    .reset(x262_sum_1_reset),
    .io_a(x262_sum_1_io_a),
    .io_b(x262_sum_1_io_b),
    .io_flow(x262_sum_1_io_flow),
    .io_result(x262_sum_1_io_result)
  );
  RetimeWrapper_162 RetimeWrapper_44 ( // @[package.scala 93:22:@25413.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_202 RetimeWrapper_45 ( // @[package.scala 93:22:@25422.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_178 RetimeWrapper_46 ( // @[package.scala 93:22:@25431.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_47 ( // @[package.scala 93:22:@25443.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  x414_sub x265_rdrow_1 ( // @[Math.scala 191:24:@25466.4]
    .clock(x265_rdrow_1_clock),
    .reset(x265_rdrow_1_reset),
    .io_a(x265_rdrow_1_io_a),
    .io_b(x265_rdrow_1_io_b),
    .io_flow(x265_rdrow_1_io_flow),
    .io_result(x265_rdrow_1_io_result)
  );
  x236 x266_1 ( // @[Math.scala 366:24:@25478.4]
    .clock(x266_1_clock),
    .reset(x266_1_reset),
    .io_a(x266_1_io_a),
    .io_flow(x266_1_io_flow),
    .io_result(x266_1_io_result)
  );
  RetimeWrapper RetimeWrapper_48 ( // @[package.scala 93:22:@25493.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper RetimeWrapper_49 ( // @[package.scala 93:22:@25502.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  fmamul_x416 x272_mul_1 ( // @[Math.scala 262:24:@25541.4]
    .clock(x272_mul_1_clock),
    .reset(x272_mul_1_reset),
    .io_a(x272_mul_1_io_a),
    .io_flow(x272_mul_1_io_flow),
    .io_result(x272_mul_1_io_result)
  );
  RetimeWrapper_232 RetimeWrapper_50 ( // @[package.scala 93:22:@25551.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x396_sum x273_sum_1 ( // @[Math.scala 150:24:@25560.4]
    .clock(x273_sum_1_clock),
    .reset(x273_sum_1_reset),
    .io_a(x273_sum_1_io_a),
    .io_b(x273_sum_1_io_b),
    .io_flow(x273_sum_1_io_flow),
    .io_result(x273_sum_1_io_result)
  );
  RetimeWrapper_202 RetimeWrapper_51 ( // @[package.scala 93:22:@25570.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_235 RetimeWrapper_52 ( // @[package.scala 93:22:@25579.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_236 RetimeWrapper_53 ( // @[package.scala 93:22:@25588.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_54 ( // @[package.scala 93:22:@25600.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_238 RetimeWrapper_55 ( // @[package.scala 93:22:@25627.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x396_sum x278_sum_1 ( // @[Math.scala 150:24:@25636.4]
    .clock(x278_sum_1_clock),
    .reset(x278_sum_1_reset),
    .io_a(x278_sum_1_io_a),
    .io_b(x278_sum_1_io_b),
    .io_flow(x278_sum_1_io_flow),
    .io_result(x278_sum_1_io_result)
  );
  RetimeWrapper_236 RetimeWrapper_56 ( // @[package.scala 93:22:@25646.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_202 RetimeWrapper_57 ( // @[package.scala 93:22:@25655.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_58 ( // @[package.scala 93:22:@25667.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_238 RetimeWrapper_59 ( // @[package.scala 93:22:@25694.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  x396_sum x283_sum_1 ( // @[Math.scala 150:24:@25703.4]
    .clock(x283_sum_1_clock),
    .reset(x283_sum_1_reset),
    .io_a(x283_sum_1_io_a),
    .io_b(x283_sum_1_io_b),
    .io_flow(x283_sum_1_io_flow),
    .io_result(x283_sum_1_io_result)
  );
  RetimeWrapper_202 RetimeWrapper_60 ( // @[package.scala 93:22:@25713.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_236 RetimeWrapper_61 ( // @[package.scala 93:22:@25722.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_62 ( // @[package.scala 93:22:@25734.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x414_sub x286_rdrow_1 ( // @[Math.scala 191:24:@25757.4]
    .clock(x286_rdrow_1_clock),
    .reset(x286_rdrow_1_reset),
    .io_a(x286_rdrow_1_io_a),
    .io_b(x286_rdrow_1_io_b),
    .io_flow(x286_rdrow_1_io_flow),
    .io_result(x286_rdrow_1_io_result)
  );
  x236 x287_1 ( // @[Math.scala 366:24:@25769.4]
    .clock(x287_1_clock),
    .reset(x287_1_reset),
    .io_a(x287_1_io_a),
    .io_flow(x287_1_io_flow),
    .io_result(x287_1_io_result)
  );
  RetimeWrapper RetimeWrapper_63 ( // @[package.scala 93:22:@25784.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  fmamul_x416 x293_mul_1 ( // @[Math.scala 262:24:@25821.4]
    .clock(x293_mul_1_clock),
    .reset(x293_mul_1_reset),
    .io_a(x293_mul_1_io_a),
    .io_flow(x293_mul_1_io_flow),
    .io_result(x293_mul_1_io_result)
  );
  x396_sum x294_sum_1 ( // @[Math.scala 150:24:@25831.4]
    .clock(x294_sum_1_clock),
    .reset(x294_sum_1_reset),
    .io_a(x294_sum_1_io_a),
    .io_b(x294_sum_1_io_b),
    .io_flow(x294_sum_1_io_flow),
    .io_result(x294_sum_1_io_result)
  );
  RetimeWrapper_235 RetimeWrapper_64 ( // @[package.scala 93:22:@25841.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_202 RetimeWrapper_65 ( // @[package.scala 93:22:@25850.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_236 RetimeWrapper_66 ( // @[package.scala 93:22:@25859.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_67 ( // @[package.scala 93:22:@25871.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x396_sum x299_sum_1 ( // @[Math.scala 150:24:@25898.4]
    .clock(x299_sum_1_clock),
    .reset(x299_sum_1_reset),
    .io_a(x299_sum_1_io_a),
    .io_b(x299_sum_1_io_b),
    .io_flow(x299_sum_1_io_flow),
    .io_result(x299_sum_1_io_result)
  );
  RetimeWrapper_202 RetimeWrapper_68 ( // @[package.scala 93:22:@25908.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_236 RetimeWrapper_69 ( // @[package.scala 93:22:@25917.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_70 ( // @[package.scala 93:22:@25929.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  x396_sum x304_sum_1 ( // @[Math.scala 150:24:@25956.4]
    .clock(x304_sum_1_clock),
    .reset(x304_sum_1_reset),
    .io_a(x304_sum_1_io_a),
    .io_b(x304_sum_1_io_b),
    .io_flow(x304_sum_1_io_flow),
    .io_result(x304_sum_1_io_result)
  );
  RetimeWrapper_202 RetimeWrapper_71 ( // @[package.scala 93:22:@25966.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_236 RetimeWrapper_72 ( // @[package.scala 93:22:@25975.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_175 RetimeWrapper_73 ( // @[package.scala 93:22:@25987.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x312_x11 x312_x11_1 ( // @[Math.scala 150:24:@26035.4]
    .clock(x312_x11_1_clock),
    .reset(x312_x11_1_reset),
    .io_a(x312_x11_1_io_a),
    .io_b(x312_x11_1_io_b),
    .io_flow(x312_x11_1_io_flow),
    .io_result(x312_x11_1_io_result)
  );
  x312_x11 x313_x12_1 ( // @[Math.scala 150:24:@26045.4]
    .clock(x313_x12_1_clock),
    .reset(x313_x12_1_reset),
    .io_a(x313_x12_1_io_a),
    .io_b(x313_x12_1_io_b),
    .io_flow(x313_x12_1_io_flow),
    .io_result(x313_x12_1_io_result)
  );
  x312_x11 x314_x11_1 ( // @[Math.scala 150:24:@26055.4]
    .clock(x314_x11_1_clock),
    .reset(x314_x11_1_reset),
    .io_a(x314_x11_1_io_a),
    .io_b(x314_x11_1_io_b),
    .io_flow(x314_x11_1_io_flow),
    .io_result(x314_x11_1_io_result)
  );
  x312_x11 x315_x12_1 ( // @[Math.scala 150:24:@26065.4]
    .clock(x315_x12_1_clock),
    .reset(x315_x12_1_reset),
    .io_a(x315_x12_1_io_a),
    .io_b(x315_x12_1_io_b),
    .io_flow(x315_x12_1_io_flow),
    .io_result(x315_x12_1_io_result)
  );
  x316_x11 x316_x11_1 ( // @[Math.scala 150:24:@26075.4]
    .io_a(x316_x11_1_io_a),
    .io_b(x316_x11_1_io_b),
    .io_result(x316_x11_1_io_result)
  );
  x316_x11 x317_x12_1 ( // @[Math.scala 150:24:@26085.4]
    .io_a(x317_x12_1_io_a),
    .io_b(x317_x12_1_io_b),
    .io_result(x317_x12_1_io_result)
  );
  x316_x11 x318_x11_1 ( // @[Math.scala 150:24:@26095.4]
    .io_a(x318_x11_1_io_a),
    .io_b(x318_x11_1_io_b),
    .io_result(x318_x11_1_io_result)
  );
  RetimeWrapper_140 RetimeWrapper_74 ( // @[package.scala 93:22:@26105.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x316_x11 x319_sum_1 ( // @[Math.scala 150:24:@26114.4]
    .io_a(x319_sum_1_io_a),
    .io_b(x319_sum_1_io_b),
    .io_result(x319_sum_1_io_result)
  );
  RetimeWrapper_140 RetimeWrapper_75 ( // @[package.scala 93:22:@26128.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_273 RetimeWrapper_76 ( // @[package.scala 93:22:@26142.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_77 ( // @[package.scala 93:22:@26151.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_78 ( // @[package.scala 93:22:@26160.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_79 ( // @[package.scala 93:22:@26169.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  assign b216 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 62:18:@24006.4]
  assign b217 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 63:18:@24007.4]
  assign _T_206 = b216 & b217; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 68:30:@24076.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 68:37:@24077.4]
  assign _T_211 = io_in_x205_TID == 8'h0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 70:76:@24082.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 70:62:@24083.4]
  assign _T_214 = io_in_x205_TDEST == 8'h0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 70:101:@24084.4]
  assign b214_number = __io_result; // @[Math.scala 712:22:@23991.4 Math.scala 713:14:@23992.4]
  assign _T_240 = $signed(b214_number); // @[Math.scala 499:52:@24107.4]
  assign x223 = $signed(32'sh1) == $signed(_T_240); // @[Math.scala 499:44:@24115.4]
  assign x224 = $signed(32'sh2) == $signed(_T_240); // @[Math.scala 499:44:@24122.4]
  assign x225 = $signed(32'sh3) == $signed(_T_240); // @[Math.scala 499:44:@24129.4]
  assign _T_287 = x223 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@24141.4]
  assign _T_289 = x224 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@24142.4]
  assign _T_291 = x225 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@24143.4]
  assign _T_293 = _T_287 | _T_289; // @[Mux.scala 19:72:@24145.4]
  assign x226_number = _T_293 | _T_291; // @[Mux.scala 19:72:@24146.4]
  assign _T_305 = $signed(x226_number); // @[Math.scala 406:49:@24156.4]
  assign _T_307 = $signed(_T_305) & $signed(32'sh3); // @[Math.scala 406:56:@24158.4]
  assign _T_308 = $signed(_T_307); // @[Math.scala 406:56:@24159.4]
  assign b215_number = __1_io_result; // @[Math.scala 712:22:@24003.4 Math.scala 713:14:@24004.4]
  assign _T_313 = b215_number[31]; // @[FixedPoint.scala 50:25:@24165.4]
  assign _T_317 = _T_313 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@24167.4]
  assign _T_318 = b215_number[31:16]; // @[FixedPoint.scala 18:52:@24168.4]
  assign _T_327 = $signed(b215_number); // @[Math.scala 406:49:@24176.4]
  assign _T_329 = $signed(_T_327) & $signed(32'shffff); // @[Math.scala 406:56:@24178.4]
  assign _T_330 = $signed(_T_329); // @[Math.scala 406:56:@24179.4]
  assign x396_sum_number = x396_sum_1_io_result; // @[Math.scala 154:22:@24190.4 Math.scala 155:14:@24191.4]
  assign _T_338 = x396_sum_number[31]; // @[FixedPoint.scala 50:25:@24195.4]
  assign _T_342 = _T_338 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@24197.4]
  assign _T_343 = x396_sum_number[31:8]; // @[FixedPoint.scala 18:52:@24198.4]
  assign _T_352 = $signed(x396_sum_number); // @[Math.scala 406:49:@24206.4]
  assign _T_354 = $signed(_T_352) & $signed(32'shff); // @[Math.scala 406:56:@24208.4]
  assign _T_355 = $signed(_T_354); // @[Math.scala 406:56:@24209.4]
  assign x399_sum_number = x399_sum_1_io_result; // @[Math.scala 154:22:@24220.4 Math.scala 155:14:@24221.4]
  assign _T_363 = x399_sum_number[31]; // @[FixedPoint.scala 50:25:@24225.4]
  assign _T_367 = _T_363 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@24227.4]
  assign _T_368 = x399_sum_number[31:4]; // @[FixedPoint.scala 18:52:@24228.4]
  assign _T_377 = $signed(x399_sum_number); // @[Math.scala 406:49:@24236.4]
  assign _T_379 = $signed(_T_377) & $signed(32'shf); // @[Math.scala 406:56:@24238.4]
  assign _T_380 = $signed(_T_379); // @[Math.scala 406:56:@24239.4]
  assign x402_sum_number = x402_sum_1_io_result; // @[Math.scala 154:22:@24250.4 Math.scala 155:14:@24251.4]
  assign _T_388 = x402_sum_number[31]; // @[FixedPoint.scala 50:25:@24255.4]
  assign _T_392 = _T_388 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24257.4]
  assign _T_393 = x402_sum_number[31:2]; // @[FixedPoint.scala 18:52:@24258.4]
  assign _T_402 = $signed(x402_sum_number); // @[Math.scala 406:49:@24266.4]
  assign _T_404 = $signed(_T_402) & $signed(32'sh3); // @[Math.scala 406:56:@24268.4]
  assign _T_405 = $signed(_T_404); // @[Math.scala 406:56:@24269.4]
  assign x405_sum_number = x405_sum_1_io_result; // @[Math.scala 154:22:@24280.4 Math.scala 155:14:@24281.4]
  assign _T_413 = x405_sum_number[31]; // @[FixedPoint.scala 50:25:@24285.4]
  assign _T_417 = _T_413 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24287.4]
  assign _T_418 = x405_sum_number[31:2]; // @[FixedPoint.scala 18:52:@24288.4]
  assign _T_429 = $signed(x405_sum_number); // @[Math.scala 406:49:@24303.4]
  assign _T_431 = $signed(_T_429) & $signed(32'sh3); // @[Math.scala 406:56:@24305.4]
  assign _T_432 = $signed(_T_431); // @[Math.scala 406:56:@24306.4]
  assign _T_436 = $signed(RetimeWrapper_2_io_out); // @[package.scala 96:25:@24314.4]
  assign x408_sum_number = x408_sum_1_io_result; // @[Math.scala 154:22:@24326.4 Math.scala 155:14:@24327.4]
  assign _T_444 = x408_sum_number[31]; // @[FixedPoint.scala 50:25:@24331.4]
  assign _T_448 = _T_444 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24333.4]
  assign _T_449 = x408_sum_number[31:2]; // @[FixedPoint.scala 18:52:@24334.4]
  assign _T_458 = $signed(x408_sum_number); // @[Math.scala 406:49:@24342.4]
  assign _T_460 = $signed(_T_458) & $signed(32'sh3); // @[Math.scala 406:56:@24344.4]
  assign _T_461 = $signed(_T_460); // @[Math.scala 406:56:@24345.4]
  assign x411_sum_number = x411_sum_1_io_result; // @[Math.scala 154:22:@24356.4 Math.scala 155:14:@24357.4]
  assign _T_471 = $signed(x411_sum_number); // @[Math.scala 465:37:@24362.4]
  assign x466_x412_D1 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@24400.4 package.scala 96:25:@24401.4]
  assign x467_x411_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@24409.4 package.scala 96:25:@24410.4]
  assign x414_sub_number = x414_sub_1_io_result; // @[Math.scala 195:22:@24382.4 Math.scala 196:14:@24383.4]
  assign _T_503 = x226_number[31]; // @[FixedPoint.scala 50:25:@24417.4]
  assign _T_507 = _T_503 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24419.4]
  assign _T_508 = x226_number[31:2]; // @[FixedPoint.scala 18:52:@24420.4]
  assign _T_546 = ~ io_sigsIn_break; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:101:@24510.4]
  assign _T_550 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@24518.4 package.scala 96:25:@24519.4]
  assign _T_552 = io_rr ? _T_550 : 1'h0; // @[implicits.scala 55:10:@24520.4]
  assign _T_553 = _T_546 & _T_552; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:118:@24521.4]
  assign _T_555 = _T_553 & _T_546; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:207:@24523.4]
  assign _T_556 = _T_555 & io_sigsIn_backpressure; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:226:@24524.4]
  assign x470_b216_D26 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@24480.4 package.scala 96:25:@24481.4]
  assign _T_557 = _T_556 & x470_b216_D26; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 165:252:@24525.4]
  assign x469_b217_D26 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@24471.4 package.scala 96:25:@24472.4]
  assign x474_b214_D28_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@24539.4 package.scala 96:25:@24540.4]
  assign _T_576 = $signed(x474_b214_D28_number); // @[Math.scala 465:37:@24559.4]
  assign x475_b215_D28_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@24576.4 package.scala 96:25:@24577.4]
  assign _T_589 = $signed(x475_b215_D28_number); // @[Math.scala 465:37:@24582.4]
  assign x237 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@24567.4 package.scala 96:25:@24568.4]
  assign x238 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@24590.4 package.scala 96:25:@24591.4]
  assign x239 = x237 | x238; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 186:24:@24594.4]
  assign x236_number = x236_1_io_result; // @[Math.scala 370:22:@24553.4 Math.scala 371:14:@24554.4]
  assign _T_605 = $signed(x236_number); // @[Math.scala 406:49:@24603.4]
  assign _T_607 = $signed(_T_605) & $signed(32'sh3); // @[Math.scala 406:56:@24605.4]
  assign _T_608 = $signed(_T_607); // @[Math.scala 406:56:@24606.4]
  assign _T_613 = x236_number[31]; // @[FixedPoint.scala 50:25:@24612.4]
  assign _T_617 = _T_613 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24614.4]
  assign _T_618 = x236_number[31:2]; // @[FixedPoint.scala 18:52:@24615.4]
  assign _T_662 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@24713.4 package.scala 96:25:@24714.4]
  assign _T_664 = io_rr ? _T_662 : 1'h0; // @[implicits.scala 55:10:@24715.4]
  assign _T_665 = _T_546 & _T_664; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 215:194:@24716.4]
  assign x481_x240_D26 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  assign _T_666 = _T_665 & x481_x240_D26; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 215:283:@24717.4]
  assign x479_b216_D55 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@24674.4 package.scala 96:25:@24675.4]
  assign _T_667 = _T_666 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 215:291:@24718.4]
  assign x477_b217_D55 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@24656.4 package.scala 96:25:@24657.4]
  assign x247_rdcol_number = x247_rdcol_1_io_result; // @[Math.scala 195:22:@24737.4 Math.scala 196:14:@24738.4]
  assign _T_682 = $signed(x247_rdcol_number); // @[Math.scala 465:37:@24743.4]
  assign x483_x237_D1 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@24760.4 package.scala 96:25:@24761.4]
  assign x248 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@24751.4 package.scala 96:25:@24752.4]
  assign x249 = x483_x237_D1 | x248; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 225:24:@24764.4]
  assign _T_697 = x247_rdcol_number[31]; // @[FixedPoint.scala 50:25:@24771.4]
  assign _T_701 = _T_697 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@24773.4]
  assign _T_702 = x247_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@24774.4]
  assign _T_713 = $signed(_T_682) & $signed(32'shffff); // @[Math.scala 406:56:@24784.4]
  assign _T_714 = $signed(_T_713); // @[Math.scala 406:56:@24785.4]
  assign x420_sum_number = x420_sum_1_io_result; // @[Math.scala 154:22:@24796.4 Math.scala 155:14:@24797.4]
  assign _T_722 = x420_sum_number[31]; // @[FixedPoint.scala 50:25:@24801.4]
  assign _T_726 = _T_722 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@24803.4]
  assign _T_727 = x420_sum_number[31:8]; // @[FixedPoint.scala 18:52:@24804.4]
  assign _T_738 = $signed(x420_sum_number); // @[Math.scala 406:49:@24819.4]
  assign _T_740 = $signed(_T_738) & $signed(32'shff); // @[Math.scala 406:56:@24821.4]
  assign _T_741 = $signed(_T_740); // @[Math.scala 406:56:@24822.4]
  assign _T_745 = $signed(RetimeWrapper_28_io_out); // @[package.scala 96:25:@24830.4]
  assign x423_sum_number = x423_sum_1_io_result; // @[Math.scala 154:22:@24842.4 Math.scala 155:14:@24843.4]
  assign _T_753 = x423_sum_number[31]; // @[FixedPoint.scala 50:25:@24847.4]
  assign _T_757 = _T_753 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@24849.4]
  assign _T_758 = x423_sum_number[31:4]; // @[FixedPoint.scala 18:52:@24850.4]
  assign _T_767 = $signed(x423_sum_number); // @[Math.scala 406:49:@24858.4]
  assign _T_769 = $signed(_T_767) & $signed(32'shf); // @[Math.scala 406:56:@24860.4]
  assign _T_770 = $signed(_T_769); // @[Math.scala 406:56:@24861.4]
  assign x426_sum_number = x426_sum_1_io_result; // @[Math.scala 154:22:@24872.4 Math.scala 155:14:@24873.4]
  assign _T_778 = x426_sum_number[31]; // @[FixedPoint.scala 50:25:@24877.4]
  assign _T_782 = _T_778 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24879.4]
  assign _T_783 = x426_sum_number[31:2]; // @[FixedPoint.scala 18:52:@24880.4]
  assign _T_792 = $signed(x426_sum_number); // @[Math.scala 406:49:@24888.4]
  assign _T_794 = $signed(_T_792) & $signed(32'sh3); // @[Math.scala 406:56:@24890.4]
  assign _T_795 = $signed(_T_794); // @[Math.scala 406:56:@24891.4]
  assign x429_sum_number = x429_sum_1_io_result; // @[Math.scala 154:22:@24902.4 Math.scala 155:14:@24903.4]
  assign _T_803 = x429_sum_number[31]; // @[FixedPoint.scala 50:25:@24907.4]
  assign _T_807 = _T_803 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24909.4]
  assign _T_808 = x429_sum_number[31:2]; // @[FixedPoint.scala 18:52:@24910.4]
  assign _T_817 = $signed(x429_sum_number); // @[Math.scala 406:49:@24918.4]
  assign _T_819 = $signed(_T_817) & $signed(32'sh3); // @[Math.scala 406:56:@24920.4]
  assign _T_820 = $signed(_T_819); // @[Math.scala 406:56:@24921.4]
  assign x432_sum_number = x432_sum_1_io_result; // @[Math.scala 154:22:@24932.4 Math.scala 155:14:@24933.4]
  assign _T_828 = x432_sum_number[31]; // @[FixedPoint.scala 50:25:@24937.4]
  assign _T_832 = _T_828 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24939.4]
  assign _T_833 = x432_sum_number[31:2]; // @[FixedPoint.scala 18:52:@24940.4]
  assign _T_842 = $signed(x432_sum_number); // @[Math.scala 406:49:@24948.4]
  assign _T_844 = $signed(_T_842) & $signed(32'sh3); // @[Math.scala 406:56:@24950.4]
  assign _T_845 = $signed(_T_844); // @[Math.scala 406:56:@24951.4]
  assign x435_sum_number = x435_sum_1_io_result; // @[Math.scala 154:22:@24962.4 Math.scala 155:14:@24963.4]
  assign _T_855 = $signed(x435_sum_number); // @[Math.scala 465:37:@24968.4]
  assign x436 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@24976.4 package.scala 96:25:@24977.4]
  assign x484_x435_sum_D1_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@25011.4 package.scala 96:25:@25012.4]
  assign x438_sub_number = x438_sub_1_io_result; // @[Math.scala 195:22:@25002.4 Math.scala 196:14:@25003.4]
  assign _T_917 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@25086.4 package.scala 96:25:@25087.4]
  assign _T_919 = io_rr ? _T_917 : 1'h0; // @[implicits.scala 55:10:@25088.4]
  assign _T_920 = _T_546 & _T_919; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:194:@25089.4]
  assign x488_x250_D25 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@25074.4 package.scala 96:25:@25075.4]
  assign _T_921 = _T_920 & x488_x250_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:283:@25090.4]
  assign _T_922 = _T_921 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:291:@25091.4]
  assign x256_rdcol_number = x256_rdcol_1_io_result; // @[Math.scala 195:22:@25110.4 Math.scala 196:14:@25111.4]
  assign _T_937 = $signed(x256_rdcol_number); // @[Math.scala 465:37:@25116.4]
  assign x257 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@25124.4 package.scala 96:25:@25125.4]
  assign x258 = x483_x237_D1 | x257; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 306:59:@25128.4]
  assign _T_949 = x256_rdcol_number[31]; // @[FixedPoint.scala 50:25:@25135.4]
  assign _T_953 = _T_949 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@25137.4]
  assign _T_954 = x256_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@25138.4]
  assign _T_965 = $signed(_T_937) & $signed(32'shffff); // @[Math.scala 406:56:@25148.4]
  assign _T_966 = $signed(_T_965); // @[Math.scala 406:56:@25149.4]
  assign x442_sum_number = x442_sum_1_io_result; // @[Math.scala 154:22:@25160.4 Math.scala 155:14:@25161.4]
  assign _T_974 = x442_sum_number[31]; // @[FixedPoint.scala 50:25:@25165.4]
  assign _T_978 = _T_974 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@25167.4]
  assign _T_979 = x442_sum_number[31:8]; // @[FixedPoint.scala 18:52:@25168.4]
  assign _T_990 = $signed(x442_sum_number); // @[Math.scala 406:49:@25183.4]
  assign _T_992 = $signed(_T_990) & $signed(32'shff); // @[Math.scala 406:56:@25185.4]
  assign _T_993 = $signed(_T_992); // @[Math.scala 406:56:@25186.4]
  assign _T_997 = $signed(RetimeWrapper_39_io_out); // @[package.scala 96:25:@25194.4]
  assign x445_sum_number = x445_sum_1_io_result; // @[Math.scala 154:22:@25206.4 Math.scala 155:14:@25207.4]
  assign _T_1005 = x445_sum_number[31]; // @[FixedPoint.scala 50:25:@25211.4]
  assign _T_1009 = _T_1005 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@25213.4]
  assign _T_1010 = x445_sum_number[31:4]; // @[FixedPoint.scala 18:52:@25214.4]
  assign _T_1019 = $signed(x445_sum_number); // @[Math.scala 406:49:@25222.4]
  assign _T_1021 = $signed(_T_1019) & $signed(32'shf); // @[Math.scala 406:56:@25224.4]
  assign _T_1022 = $signed(_T_1021); // @[Math.scala 406:56:@25225.4]
  assign x448_sum_number = x448_sum_1_io_result; // @[Math.scala 154:22:@25236.4 Math.scala 155:14:@25237.4]
  assign _T_1030 = x448_sum_number[31]; // @[FixedPoint.scala 50:25:@25241.4]
  assign _T_1034 = _T_1030 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25243.4]
  assign _T_1035 = x448_sum_number[31:2]; // @[FixedPoint.scala 18:52:@25244.4]
  assign _T_1044 = $signed(x448_sum_number); // @[Math.scala 406:49:@25252.4]
  assign _T_1046 = $signed(_T_1044) & $signed(32'sh3); // @[Math.scala 406:56:@25254.4]
  assign _T_1047 = $signed(_T_1046); // @[Math.scala 406:56:@25255.4]
  assign x451_sum_number = x451_sum_1_io_result; // @[Math.scala 154:22:@25266.4 Math.scala 155:14:@25267.4]
  assign _T_1055 = x451_sum_number[31]; // @[FixedPoint.scala 50:25:@25271.4]
  assign _T_1059 = _T_1055 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25273.4]
  assign _T_1060 = x451_sum_number[31:2]; // @[FixedPoint.scala 18:52:@25274.4]
  assign _T_1069 = $signed(x451_sum_number); // @[Math.scala 406:49:@25282.4]
  assign _T_1071 = $signed(_T_1069) & $signed(32'sh3); // @[Math.scala 406:56:@25284.4]
  assign _T_1072 = $signed(_T_1071); // @[Math.scala 406:56:@25285.4]
  assign x454_sum_number = x454_sum_1_io_result; // @[Math.scala 154:22:@25296.4 Math.scala 155:14:@25297.4]
  assign _T_1080 = x454_sum_number[31]; // @[FixedPoint.scala 50:25:@25301.4]
  assign _T_1084 = _T_1080 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25303.4]
  assign _T_1085 = x454_sum_number[31:2]; // @[FixedPoint.scala 18:52:@25304.4]
  assign _T_1094 = $signed(x454_sum_number); // @[Math.scala 406:49:@25312.4]
  assign _T_1096 = $signed(_T_1094) & $signed(32'sh3); // @[Math.scala 406:56:@25314.4]
  assign _T_1097 = $signed(_T_1096); // @[Math.scala 406:56:@25315.4]
  assign x457_sum_number = x457_sum_1_io_result; // @[Math.scala 154:22:@25326.4 Math.scala 155:14:@25327.4]
  assign _T_1107 = $signed(x457_sum_number); // @[Math.scala 465:37:@25332.4]
  assign x458 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@25340.4 package.scala 96:25:@25341.4]
  assign x489_x457_sum_D1_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@25375.4 package.scala 96:25:@25376.4]
  assign x460_sub_number = x460_sub_1_io_result; // @[Math.scala 195:22:@25366.4 Math.scala 196:14:@25367.4]
  assign _T_1167 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@25448.4 package.scala 96:25:@25449.4]
  assign _T_1169 = io_rr ? _T_1167 : 1'h0; // @[implicits.scala 55:10:@25450.4]
  assign _T_1170 = _T_546 & _T_1169; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 371:194:@25451.4]
  assign x492_x259_D25 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@25427.4 package.scala 96:25:@25428.4]
  assign _T_1171 = _T_1170 & x492_x259_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 371:283:@25452.4]
  assign _T_1172 = _T_1171 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 371:291:@25453.4]
  assign x265_rdrow_number = x265_rdrow_1_io_result; // @[Math.scala 195:22:@25472.4 Math.scala 196:14:@25473.4]
  assign _T_1194 = $signed(x265_rdrow_number); // @[Math.scala 465:37:@25490.4]
  assign x267 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@25498.4 package.scala 96:25:@25499.4]
  assign x494_x238_D1 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@25507.4 package.scala 96:25:@25508.4]
  assign x268 = x267 | x494_x238_D1; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 383:24:@25511.4]
  assign x266_number = x266_1_io_result; // @[Math.scala 370:22:@25484.4 Math.scala 371:14:@25485.4]
  assign _T_1213 = $signed(x266_number); // @[Math.scala 406:49:@25520.4]
  assign _T_1215 = $signed(_T_1213) & $signed(32'sh3); // @[Math.scala 406:56:@25522.4]
  assign _T_1216 = $signed(_T_1215); // @[Math.scala 406:56:@25523.4]
  assign _T_1221 = x266_number[31]; // @[FixedPoint.scala 50:25:@25529.4]
  assign _T_1225 = _T_1221 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25531.4]
  assign _T_1226 = x266_number[31:2]; // @[FixedPoint.scala 18:52:@25532.4]
  assign _T_1263 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@25605.4 package.scala 96:25:@25606.4]
  assign _T_1265 = io_rr ? _T_1263 : 1'h0; // @[implicits.scala 55:10:@25607.4]
  assign _T_1266 = _T_546 & _T_1265; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:194:@25608.4]
  assign x496_x269_D25 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@25575.4 package.scala 96:25:@25576.4]
  assign _T_1267 = _T_1266 & x496_x269_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:283:@25609.4]
  assign _T_1268 = _T_1267 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:291:@25610.4]
  assign x276 = x267 | x248; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 418:59:@25621.4]
  assign _T_1298 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@25672.4 package.scala 96:25:@25673.4]
  assign _T_1300 = io_rr ? _T_1298 : 1'h0; // @[implicits.scala 55:10:@25674.4]
  assign _T_1301 = _T_546 & _T_1300; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:194:@25675.4]
  assign x501_x277_D25 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@25660.4 package.scala 96:25:@25661.4]
  assign _T_1302 = _T_1301 & x501_x277_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:283:@25676.4]
  assign _T_1303 = _T_1302 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:291:@25677.4]
  assign x281 = x267 | x257; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 437:59:@25688.4]
  assign _T_1333 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@25739.4 package.scala 96:25:@25740.4]
  assign _T_1335 = io_rr ? _T_1333 : 1'h0; // @[implicits.scala 55:10:@25741.4]
  assign _T_1336 = _T_546 & _T_1335; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:194:@25742.4]
  assign x503_x282_D25 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@25718.4 package.scala 96:25:@25719.4]
  assign _T_1337 = _T_1336 & x503_x282_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:283:@25743.4]
  assign _T_1338 = _T_1337 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:291:@25744.4]
  assign x286_rdrow_number = x286_rdrow_1_io_result; // @[Math.scala 195:22:@25763.4 Math.scala 196:14:@25764.4]
  assign _T_1360 = $signed(x286_rdrow_number); // @[Math.scala 465:37:@25781.4]
  assign x288 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@25789.4 package.scala 96:25:@25790.4]
  assign x289 = x288 | x494_x238_D1; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 462:24:@25793.4]
  assign x287_number = x287_1_io_result; // @[Math.scala 370:22:@25775.4 Math.scala 371:14:@25776.4]
  assign _T_1376 = $signed(x287_number); // @[Math.scala 406:49:@25802.4]
  assign _T_1378 = $signed(_T_1376) & $signed(32'sh3); // @[Math.scala 406:56:@25804.4]
  assign _T_1379 = $signed(_T_1378); // @[Math.scala 406:56:@25805.4]
  assign _T_1384 = x287_number[31]; // @[FixedPoint.scala 50:25:@25811.4]
  assign _T_1388 = _T_1384 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25813.4]
  assign _T_1389 = x287_number[31:2]; // @[FixedPoint.scala 18:52:@25814.4]
  assign _T_1421 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@25876.4 package.scala 96:25:@25877.4]
  assign _T_1423 = io_rr ? _T_1421 : 1'h0; // @[implicits.scala 55:10:@25878.4]
  assign _T_1424 = _T_546 & _T_1423; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 483:194:@25879.4]
  assign x506_x290_D25 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@25855.4 package.scala 96:25:@25856.4]
  assign _T_1425 = _T_1424 & x506_x290_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 483:283:@25880.4]
  assign _T_1426 = _T_1425 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 483:291:@25881.4]
  assign x297 = x288 | x248; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 487:24:@25892.4]
  assign _T_1453 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@25934.4 package.scala 96:25:@25935.4]
  assign _T_1455 = io_rr ? _T_1453 : 1'h0; // @[implicits.scala 55:10:@25936.4]
  assign _T_1456 = _T_546 & _T_1455; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:194:@25937.4]
  assign x508_x298_D25 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@25913.4 package.scala 96:25:@25914.4]
  assign _T_1457 = _T_1456 & x508_x298_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:283:@25938.4]
  assign _T_1458 = _T_1457 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:291:@25939.4]
  assign x302 = x288 | x257; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 504:24:@25950.4]
  assign _T_1485 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@25992.4 package.scala 96:25:@25993.4]
  assign _T_1487 = io_rr ? _T_1485 : 1'h0; // @[implicits.scala 55:10:@25994.4]
  assign _T_1488 = _T_546 & _T_1487; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 523:194:@25995.4]
  assign x510_x303_D25 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@25971.4 package.scala 96:25:@25972.4]
  assign _T_1489 = _T_1488 & x510_x303_D25; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 523:283:@25996.4]
  assign _T_1490 = _T_1489 & x479_b216_D55; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 523:326:@25997.4]
  assign x254_rd_0_number = x218_lb_0_io_rPort_8_output_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 294:29:@25077.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 298:408:@25098.4]
  assign _GEN_0 = {{1'd0}, x254_rd_0_number}; // @[Math.scala 450:32:@26011.4]
  assign _T_1498 = _GEN_0 << 1; // @[Math.scala 450:32:@26011.4]
  assign x274_rd_0_number = x218_lb_0_io_rPort_2_output_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 410:29:@25596.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 414:408:@25617.4]
  assign _GEN_1 = {{1'd0}, x274_rd_0_number}; // @[Math.scala 450:32:@26016.4]
  assign _T_1502 = _GEN_1 << 1; // @[Math.scala 450:32:@26016.4]
  assign x279_rd_0_number = x218_lb_0_io_rPort_1_output_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 429:29:@25663.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 433:408:@25684.4]
  assign _GEN_2 = {{2'd0}, x279_rd_0_number}; // @[Math.scala 450:32:@26021.4]
  assign _T_1506 = _GEN_2 << 2; // @[Math.scala 450:32:@26021.4]
  assign x284_rd_0_number = x218_lb_0_io_rPort_0_output_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 448:29:@25730.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 452:408:@25751.4]
  assign _GEN_3 = {{1'd0}, x284_rd_0_number}; // @[Math.scala 450:32:@26026.4]
  assign _T_1510 = _GEN_3 << 1; // @[Math.scala 450:32:@26026.4]
  assign x300_rd_0_number = x218_lb_0_io_rPort_6_output_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 496:29:@25925.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 500:408:@25946.4]
  assign _GEN_4 = {{1'd0}, x300_rd_0_number}; // @[Math.scala 450:32:@26031.4]
  assign _T_1514 = _GEN_4 << 1; // @[Math.scala 450:32:@26031.4]
  assign x319_sum_number = x319_sum_1_io_result; // @[Math.scala 154:22:@26120.4 Math.scala 155:14:@26121.4]
  assign _T_1550 = x319_sum_number[7:4]; // @[FixedPoint.scala 18:52:@26126.4]
  assign _T_1573 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@26174.4 package.scala 96:25:@26175.4]
  assign _T_1575 = io_rr ? _T_1573 : 1'h0; // @[implicits.scala 55:10:@26176.4]
  assign x513_b216_D62 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@26156.4 package.scala 96:25:@26157.4]
  assign _T_1576 = _T_1575 & x513_b216_D62; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 567:117:@26177.4]
  assign x514_b217_D62 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@26165.4 package.scala 96:25:@26166.4]
  assign _T_1577 = _T_1576 & x514_b217_D62; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 567:123:@26178.4]
  assign x416_number = cast_x416_io_result; // @[Math.scala 712:22:@24462.4 Math.scala 713:14:@24463.4]
  assign x471_x393_D26_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@24489.4 package.scala 96:25:@24490.4]
  assign x472_x415_D18_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@24498.4 package.scala 96:25:@24499.4]
  assign x478_x417_D11_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@24665.4 package.scala 96:25:@24666.4]
  assign x480_x244_sum_D4_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@24683.4 package.scala 96:25:@24684.4]
  assign x482_x415_D47_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@24701.4 package.scala 96:25:@24702.4]
  assign x486_x253_sum_D4_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@25056.4 package.scala 96:25:@25057.4]
  assign x487_x439_D18_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@25065.4 package.scala 96:25:@25066.4]
  assign x491_x461_D18_number = RetimeWrapper_44_io_out; // @[package.scala 96:25:@25418.4 package.scala 96:25:@25419.4]
  assign x493_x262_sum_D4_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@25436.4 package.scala 96:25:@25437.4]
  assign x497_x462_D10_number = RetimeWrapper_52_io_out; // @[package.scala 96:25:@25584.4 package.scala 96:25:@25585.4]
  assign x498_x273_sum_D3_number = RetimeWrapper_53_io_out; // @[package.scala 96:25:@25593.4 package.scala 96:25:@25594.4]
  assign x500_x278_sum_D3_number = RetimeWrapper_56_io_out; // @[package.scala 96:25:@25651.4 package.scala 96:25:@25652.4]
  assign x504_x283_sum_D3_number = RetimeWrapper_61_io_out; // @[package.scala 96:25:@25727.4 package.scala 96:25:@25728.4]
  assign x505_x463_D10_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@25846.4 package.scala 96:25:@25847.4]
  assign x507_x294_sum_D3_number = RetimeWrapper_66_io_out; // @[package.scala 96:25:@25864.4 package.scala 96:25:@25865.4]
  assign x509_x299_sum_D3_number = RetimeWrapper_69_io_out; // @[package.scala 96:25:@25922.4 package.scala 96:25:@25923.4]
  assign x511_x304_sum_D3_number = RetimeWrapper_72_io_out; // @[package.scala 96:25:@25980.4 package.scala 96:25:@25981.4]
  assign io_in_x206_TVALID = _T_1577 & io_sigsIn_backpressure; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 567:22:@26180.4]
  assign io_in_x206_TDATA = {{248'd0}, RetimeWrapper_76_io_out}; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 568:24:@26181.4]
  assign io_in_x205_TREADY = _T_212 & _T_214; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 68:22:@24078.4 sm_x325_inr_Foreach_SAMPLER_BOX.scala 70:22:@24086.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@23989.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@24001.4]
  assign x218_lb_0_clock = clock; // @[:@24009.4]
  assign x218_lb_0_reset = reset; // @[:@24010.4]
  assign x218_lb_0_io_rPort_8_banks_1 = x487_x439_D18_number[1:0]; // @[MemInterfaceType.scala 106:58:@25094.4]
  assign x218_lb_0_io_rPort_8_banks_0 = x478_x417_D11_number[2:0]; // @[MemInterfaceType.scala 106:58:@25093.4]
  assign x218_lb_0_io_rPort_8_ofs_0 = x486_x253_sum_D4_number[8:0]; // @[MemInterfaceType.scala 107:54:@25095.4]
  assign x218_lb_0_io_rPort_8_en_0 = _T_922 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@25097.4]
  assign x218_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25096.4]
  assign x218_lb_0_io_rPort_7_banks_1 = x491_x461_D18_number[1:0]; // @[MemInterfaceType.scala 106:58:@26000.4]
  assign x218_lb_0_io_rPort_7_banks_0 = x505_x463_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@25999.4]
  assign x218_lb_0_io_rPort_7_ofs_0 = x511_x304_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@26001.4]
  assign x218_lb_0_io_rPort_7_en_0 = _T_1490 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@26003.4]
  assign x218_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26002.4]
  assign x218_lb_0_io_rPort_6_banks_1 = x487_x439_D18_number[1:0]; // @[MemInterfaceType.scala 106:58:@25942.4]
  assign x218_lb_0_io_rPort_6_banks_0 = x505_x463_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@25941.4]
  assign x218_lb_0_io_rPort_6_ofs_0 = x509_x299_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25943.4]
  assign x218_lb_0_io_rPort_6_en_0 = _T_1458 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@25945.4]
  assign x218_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25944.4]
  assign x218_lb_0_io_rPort_5_banks_1 = x491_x461_D18_number[1:0]; // @[MemInterfaceType.scala 106:58:@25456.4]
  assign x218_lb_0_io_rPort_5_banks_0 = x478_x417_D11_number[2:0]; // @[MemInterfaceType.scala 106:58:@25455.4]
  assign x218_lb_0_io_rPort_5_ofs_0 = x493_x262_sum_D4_number[8:0]; // @[MemInterfaceType.scala 107:54:@25457.4]
  assign x218_lb_0_io_rPort_5_en_0 = _T_1172 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@25459.4]
  assign x218_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25458.4]
  assign x218_lb_0_io_rPort_4_banks_1 = x482_x415_D47_number[1:0]; // @[MemInterfaceType.scala 106:58:@25884.4]
  assign x218_lb_0_io_rPort_4_banks_0 = x505_x463_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@25883.4]
  assign x218_lb_0_io_rPort_4_ofs_0 = x507_x294_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25885.4]
  assign x218_lb_0_io_rPort_4_en_0 = _T_1426 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@25887.4]
  assign x218_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25886.4]
  assign x218_lb_0_io_rPort_3_banks_1 = x482_x415_D47_number[1:0]; // @[MemInterfaceType.scala 106:58:@24721.4]
  assign x218_lb_0_io_rPort_3_banks_0 = x478_x417_D11_number[2:0]; // @[MemInterfaceType.scala 106:58:@24720.4]
  assign x218_lb_0_io_rPort_3_ofs_0 = x480_x244_sum_D4_number[8:0]; // @[MemInterfaceType.scala 107:54:@24722.4]
  assign x218_lb_0_io_rPort_3_en_0 = _T_667 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@24724.4]
  assign x218_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24723.4]
  assign x218_lb_0_io_rPort_2_banks_1 = x482_x415_D47_number[1:0]; // @[MemInterfaceType.scala 106:58:@25613.4]
  assign x218_lb_0_io_rPort_2_banks_0 = x497_x462_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@25612.4]
  assign x218_lb_0_io_rPort_2_ofs_0 = x498_x273_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25614.4]
  assign x218_lb_0_io_rPort_2_en_0 = _T_1268 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@25616.4]
  assign x218_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25615.4]
  assign x218_lb_0_io_rPort_1_banks_1 = x487_x439_D18_number[1:0]; // @[MemInterfaceType.scala 106:58:@25680.4]
  assign x218_lb_0_io_rPort_1_banks_0 = x497_x462_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@25679.4]
  assign x218_lb_0_io_rPort_1_ofs_0 = x500_x278_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25681.4]
  assign x218_lb_0_io_rPort_1_en_0 = _T_1303 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@25683.4]
  assign x218_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25682.4]
  assign x218_lb_0_io_rPort_0_banks_1 = x491_x461_D18_number[1:0]; // @[MemInterfaceType.scala 106:58:@25747.4]
  assign x218_lb_0_io_rPort_0_banks_0 = x497_x462_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@25746.4]
  assign x218_lb_0_io_rPort_0_ofs_0 = x504_x283_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25748.4]
  assign x218_lb_0_io_rPort_0_en_0 = _T_1338 & x477_b217_D55; // @[MemInterfaceType.scala 110:79:@25750.4]
  assign x218_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25749.4]
  assign x218_lb_0_io_wPort_0_banks_1 = x472_x415_D18_number[1:0]; // @[MemInterfaceType.scala 88:58:@24528.4]
  assign x218_lb_0_io_wPort_0_banks_0 = x471_x393_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@24527.4]
  assign x218_lb_0_io_wPort_0_ofs_0 = x416_number[8:0]; // @[MemInterfaceType.scala 89:54:@24529.4]
  assign x218_lb_0_io_wPort_0_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@24530.4]
  assign x218_lb_0_io_wPort_0_en_0 = _T_557 & x469_b217_D26; // @[MemInterfaceType.scala 93:57:@24532.4]
  assign RetimeWrapper_clock = clock; // @[:@24089.4]
  assign RetimeWrapper_reset = reset; // @[:@24090.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24092.4]
  assign RetimeWrapper_io_in = io_in_x205_TDATA[7:0]; // @[package.scala 94:16:@24091.4]
  assign x396_sum_1_clock = clock; // @[:@24185.4]
  assign x396_sum_1_reset = reset; // @[:@24186.4]
  assign x396_sum_1_io_a = {_T_317,_T_318}; // @[Math.scala 151:17:@24187.4]
  assign x396_sum_1_io_b = $unsigned(_T_330); // @[Math.scala 152:17:@24188.4]
  assign x396_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24189.4]
  assign x399_sum_1_clock = clock; // @[:@24215.4]
  assign x399_sum_1_reset = reset; // @[:@24216.4]
  assign x399_sum_1_io_a = {_T_342,_T_343}; // @[Math.scala 151:17:@24217.4]
  assign x399_sum_1_io_b = $unsigned(_T_355); // @[Math.scala 152:17:@24218.4]
  assign x399_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24219.4]
  assign x402_sum_1_clock = clock; // @[:@24245.4]
  assign x402_sum_1_reset = reset; // @[:@24246.4]
  assign x402_sum_1_io_a = {_T_367,_T_368}; // @[Math.scala 151:17:@24247.4]
  assign x402_sum_1_io_b = $unsigned(_T_380); // @[Math.scala 152:17:@24248.4]
  assign x402_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24249.4]
  assign x405_sum_1_clock = clock; // @[:@24275.4]
  assign x405_sum_1_reset = reset; // @[:@24276.4]
  assign x405_sum_1_io_a = {_T_392,_T_393}; // @[Math.scala 151:17:@24277.4]
  assign x405_sum_1_io_b = $unsigned(_T_405); // @[Math.scala 152:17:@24278.4]
  assign x405_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24279.4]
  assign RetimeWrapper_1_clock = clock; // @[:@24291.4]
  assign RetimeWrapper_1_reset = reset; // @[:@24292.4]
  assign RetimeWrapper_1_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24294.4]
  assign RetimeWrapper_1_io_in = {_T_417,_T_418}; // @[package.scala 94:16:@24293.4]
  assign RetimeWrapper_2_clock = clock; // @[:@24308.4]
  assign RetimeWrapper_2_reset = reset; // @[:@24309.4]
  assign RetimeWrapper_2_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24312.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_432); // @[package.scala 94:16:@24311.4]
  assign x408_sum_1_clock = clock; // @[:@24321.4]
  assign x408_sum_1_reset = reset; // @[:@24322.4]
  assign x408_sum_1_io_a = RetimeWrapper_1_io_out; // @[Math.scala 151:17:@24323.4]
  assign x408_sum_1_io_b = $unsigned(_T_436); // @[Math.scala 152:17:@24324.4]
  assign x408_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24325.4]
  assign x411_sum_1_clock = clock; // @[:@24351.4]
  assign x411_sum_1_reset = reset; // @[:@24352.4]
  assign x411_sum_1_io_a = {_T_448,_T_449}; // @[Math.scala 151:17:@24353.4]
  assign x411_sum_1_io_b = $unsigned(_T_461); // @[Math.scala 152:17:@24354.4]
  assign x411_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24355.4]
  assign x414_sub_1_clock = clock; // @[:@24377.4]
  assign x414_sub_1_reset = reset; // @[:@24378.4]
  assign x414_sub_1_io_a = x411_sum_1_io_result; // @[Math.scala 192:17:@24379.4]
  assign x414_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@24380.4]
  assign x414_sub_1_io_flow = io_in_x206_TREADY; // @[Math.scala 194:20:@24381.4]
  assign RetimeWrapper_3_clock = clock; // @[:@24387.4]
  assign RetimeWrapper_3_reset = reset; // @[:@24388.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24390.4]
  assign RetimeWrapper_3_io_in = $signed(_T_471) < $signed(32'sh6); // @[package.scala 94:16:@24389.4]
  assign RetimeWrapper_4_clock = clock; // @[:@24396.4]
  assign RetimeWrapper_4_reset = reset; // @[:@24397.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24399.4]
  assign RetimeWrapper_4_io_in = $signed(_T_471) < $signed(32'sh3); // @[package.scala 94:16:@24398.4]
  assign RetimeWrapper_5_clock = clock; // @[:@24405.4]
  assign RetimeWrapper_5_reset = reset; // @[:@24406.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24408.4]
  assign RetimeWrapper_5_io_in = x411_sum_1_io_result; // @[package.scala 94:16:@24407.4]
  assign x232_div_1_clock = clock; // @[:@24428.4]
  assign x232_div_1_reset = reset; // @[:@24429.4]
  assign x232_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@24430.4]
  assign x232_div_1_io_flow = io_in_x206_TREADY; // @[Math.scala 330:20:@24432.4]
  assign RetimeWrapper_6_clock = clock; // @[:@24438.4]
  assign RetimeWrapper_6_reset = reset; // @[:@24439.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24441.4]
  assign RetimeWrapper_6_io_in = {_T_507,_T_508}; // @[package.scala 94:16:@24440.4]
  assign x416_1_clock = clock; // @[:@24449.4]
  assign x416_1_reset = reset; // @[:@24450.4]
  assign x416_1_io_m0 = RetimeWrapper_6_io_out; // @[Math.scala 850:18:@24451.4]
  assign x416_1_io_add = x232_div_1_io_result; // @[Math.scala 852:19:@24453.4]
  assign x416_1_io_flow = io_in_x206_TREADY; // @[Math.scala 853:20:@24454.4]
  assign cast_x416_io_b = x416_1_io_result; // @[Math.scala 710:17:@24460.4]
  assign RetimeWrapper_7_clock = clock; // @[:@24467.4]
  assign RetimeWrapper_7_reset = reset; // @[:@24468.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24470.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@24469.4]
  assign RetimeWrapper_8_clock = clock; // @[:@24476.4]
  assign RetimeWrapper_8_reset = reset; // @[:@24477.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24479.4]
  assign RetimeWrapper_8_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@24478.4]
  assign RetimeWrapper_9_clock = clock; // @[:@24485.4]
  assign RetimeWrapper_9_reset = reset; // @[:@24486.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24488.4]
  assign RetimeWrapper_9_io_in = $unsigned(_T_308); // @[package.scala 94:16:@24487.4]
  assign RetimeWrapper_10_clock = clock; // @[:@24494.4]
  assign RetimeWrapper_10_reset = reset; // @[:@24495.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24497.4]
  assign RetimeWrapper_10_io_in = x466_x412_D1 ? x467_x411_sum_D1_number : x414_sub_number; // @[package.scala 94:16:@24496.4]
  assign RetimeWrapper_11_clock = clock; // @[:@24503.4]
  assign RetimeWrapper_11_reset = reset; // @[:@24504.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24506.4]
  assign RetimeWrapper_11_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@24505.4]
  assign RetimeWrapper_12_clock = clock; // @[:@24514.4]
  assign RetimeWrapper_12_reset = reset; // @[:@24515.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24517.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24516.4]
  assign RetimeWrapper_13_clock = clock; // @[:@24535.4]
  assign RetimeWrapper_13_reset = reset; // @[:@24536.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24538.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@24537.4]
  assign x236_1_clock = clock; // @[:@24548.4]
  assign x236_1_reset = reset; // @[:@24549.4]
  assign x236_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 367:17:@24550.4]
  assign x236_1_io_flow = io_in_x206_TREADY; // @[Math.scala 369:20:@24552.4]
  assign RetimeWrapper_14_clock = clock; // @[:@24563.4]
  assign RetimeWrapper_14_reset = reset; // @[:@24564.4]
  assign RetimeWrapper_14_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24566.4]
  assign RetimeWrapper_14_io_in = $signed(_T_576) < $signed(32'sh0); // @[package.scala 94:16:@24565.4]
  assign RetimeWrapper_15_clock = clock; // @[:@24572.4]
  assign RetimeWrapper_15_reset = reset; // @[:@24573.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24575.4]
  assign RetimeWrapper_15_io_in = __1_io_result; // @[package.scala 94:16:@24574.4]
  assign RetimeWrapper_16_clock = clock; // @[:@24586.4]
  assign RetimeWrapper_16_reset = reset; // @[:@24587.4]
  assign RetimeWrapper_16_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24589.4]
  assign RetimeWrapper_16_io_in = $signed(_T_589) < $signed(32'sh0); // @[package.scala 94:16:@24588.4]
  assign x243_mul_1_clock = clock; // @[:@24623.4]
  assign x243_mul_1_reset = reset; // @[:@24624.4]
  assign x243_mul_1_io_a = {_T_617,_T_618}; // @[Math.scala 263:17:@24625.4]
  assign x243_mul_1_io_flow = io_in_x206_TREADY; // @[Math.scala 265:20:@24627.4]
  assign RetimeWrapper_17_clock = clock; // @[:@24633.4]
  assign RetimeWrapper_17_reset = reset; // @[:@24634.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24636.4]
  assign RetimeWrapper_17_io_in = x232_div_1_io_result; // @[package.scala 94:16:@24635.4]
  assign x244_sum_1_clock = clock; // @[:@24642.4]
  assign x244_sum_1_reset = reset; // @[:@24643.4]
  assign x244_sum_1_io_a = x243_mul_1_io_result; // @[Math.scala 151:17:@24644.4]
  assign x244_sum_1_io_b = RetimeWrapper_17_io_out; // @[Math.scala 152:17:@24645.4]
  assign x244_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24646.4]
  assign RetimeWrapper_18_clock = clock; // @[:@24652.4]
  assign RetimeWrapper_18_reset = reset; // @[:@24653.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24655.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@24654.4]
  assign RetimeWrapper_19_clock = clock; // @[:@24661.4]
  assign RetimeWrapper_19_reset = reset; // @[:@24662.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24664.4]
  assign RetimeWrapper_19_io_in = $unsigned(_T_608); // @[package.scala 94:16:@24663.4]
  assign RetimeWrapper_20_clock = clock; // @[:@24670.4]
  assign RetimeWrapper_20_reset = reset; // @[:@24671.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24673.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@24672.4]
  assign RetimeWrapper_21_clock = clock; // @[:@24679.4]
  assign RetimeWrapper_21_reset = reset; // @[:@24680.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24682.4]
  assign RetimeWrapper_21_io_in = x244_sum_1_io_result; // @[package.scala 94:16:@24681.4]
  assign RetimeWrapper_22_clock = clock; // @[:@24688.4]
  assign RetimeWrapper_22_reset = reset; // @[:@24689.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24691.4]
  assign RetimeWrapper_22_io_in = ~ x239; // @[package.scala 94:16:@24690.4]
  assign RetimeWrapper_23_clock = clock; // @[:@24697.4]
  assign RetimeWrapper_23_reset = reset; // @[:@24698.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24700.4]
  assign RetimeWrapper_23_io_in = x466_x412_D1 ? x467_x411_sum_D1_number : x414_sub_number; // @[package.scala 94:16:@24699.4]
  assign RetimeWrapper_24_clock = clock; // @[:@24709.4]
  assign RetimeWrapper_24_reset = reset; // @[:@24710.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24712.4]
  assign RetimeWrapper_24_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24711.4]
  assign x247_rdcol_1_clock = clock; // @[:@24732.4]
  assign x247_rdcol_1_reset = reset; // @[:@24733.4]
  assign x247_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@24734.4]
  assign x247_rdcol_1_io_b = 32'h1; // @[Math.scala 193:17:@24735.4]
  assign x247_rdcol_1_io_flow = io_in_x206_TREADY; // @[Math.scala 194:20:@24736.4]
  assign RetimeWrapper_25_clock = clock; // @[:@24747.4]
  assign RetimeWrapper_25_reset = reset; // @[:@24748.4]
  assign RetimeWrapper_25_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24750.4]
  assign RetimeWrapper_25_io_in = $signed(_T_682) < $signed(32'sh0); // @[package.scala 94:16:@24749.4]
  assign RetimeWrapper_26_clock = clock; // @[:@24756.4]
  assign RetimeWrapper_26_reset = reset; // @[:@24757.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24759.4]
  assign RetimeWrapper_26_io_in = RetimeWrapper_14_io_out; // @[package.scala 94:16:@24758.4]
  assign x420_sum_1_clock = clock; // @[:@24791.4]
  assign x420_sum_1_reset = reset; // @[:@24792.4]
  assign x420_sum_1_io_a = {_T_701,_T_702}; // @[Math.scala 151:17:@24793.4]
  assign x420_sum_1_io_b = $unsigned(_T_714); // @[Math.scala 152:17:@24794.4]
  assign x420_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24795.4]
  assign RetimeWrapper_27_clock = clock; // @[:@24807.4]
  assign RetimeWrapper_27_reset = reset; // @[:@24808.4]
  assign RetimeWrapper_27_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24810.4]
  assign RetimeWrapper_27_io_in = {_T_726,_T_727}; // @[package.scala 94:16:@24809.4]
  assign RetimeWrapper_28_clock = clock; // @[:@24824.4]
  assign RetimeWrapper_28_reset = reset; // @[:@24825.4]
  assign RetimeWrapper_28_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24828.4]
  assign RetimeWrapper_28_io_in = $unsigned(_T_741); // @[package.scala 94:16:@24827.4]
  assign x423_sum_1_clock = clock; // @[:@24837.4]
  assign x423_sum_1_reset = reset; // @[:@24838.4]
  assign x423_sum_1_io_a = RetimeWrapper_27_io_out; // @[Math.scala 151:17:@24839.4]
  assign x423_sum_1_io_b = $unsigned(_T_745); // @[Math.scala 152:17:@24840.4]
  assign x423_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24841.4]
  assign x426_sum_1_clock = clock; // @[:@24867.4]
  assign x426_sum_1_reset = reset; // @[:@24868.4]
  assign x426_sum_1_io_a = {_T_757,_T_758}; // @[Math.scala 151:17:@24869.4]
  assign x426_sum_1_io_b = $unsigned(_T_770); // @[Math.scala 152:17:@24870.4]
  assign x426_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24871.4]
  assign x429_sum_1_clock = clock; // @[:@24897.4]
  assign x429_sum_1_reset = reset; // @[:@24898.4]
  assign x429_sum_1_io_a = {_T_782,_T_783}; // @[Math.scala 151:17:@24899.4]
  assign x429_sum_1_io_b = $unsigned(_T_795); // @[Math.scala 152:17:@24900.4]
  assign x429_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24901.4]
  assign x432_sum_1_clock = clock; // @[:@24927.4]
  assign x432_sum_1_reset = reset; // @[:@24928.4]
  assign x432_sum_1_io_a = {_T_807,_T_808}; // @[Math.scala 151:17:@24929.4]
  assign x432_sum_1_io_b = $unsigned(_T_820); // @[Math.scala 152:17:@24930.4]
  assign x432_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24931.4]
  assign x435_sum_1_clock = clock; // @[:@24957.4]
  assign x435_sum_1_reset = reset; // @[:@24958.4]
  assign x435_sum_1_io_a = {_T_832,_T_833}; // @[Math.scala 151:17:@24959.4]
  assign x435_sum_1_io_b = $unsigned(_T_845); // @[Math.scala 152:17:@24960.4]
  assign x435_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@24961.4]
  assign RetimeWrapper_29_clock = clock; // @[:@24972.4]
  assign RetimeWrapper_29_reset = reset; // @[:@24973.4]
  assign RetimeWrapper_29_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24975.4]
  assign RetimeWrapper_29_io_in = $signed(_T_855) < $signed(32'sh3); // @[package.scala 94:16:@24974.4]
  assign RetimeWrapper_30_clock = clock; // @[:@24986.4]
  assign RetimeWrapper_30_reset = reset; // @[:@24987.4]
  assign RetimeWrapper_30_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@24989.4]
  assign RetimeWrapper_30_io_in = $signed(_T_855) < $signed(32'sh6); // @[package.scala 94:16:@24988.4]
  assign x438_sub_1_clock = clock; // @[:@24997.4]
  assign x438_sub_1_reset = reset; // @[:@24998.4]
  assign x438_sub_1_io_a = x435_sum_1_io_result; // @[Math.scala 192:17:@24999.4]
  assign x438_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@25000.4]
  assign x438_sub_1_io_flow = io_in_x206_TREADY; // @[Math.scala 194:20:@25001.4]
  assign RetimeWrapper_31_clock = clock; // @[:@25007.4]
  assign RetimeWrapper_31_reset = reset; // @[:@25008.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25010.4]
  assign RetimeWrapper_31_io_in = x435_sum_1_io_result; // @[package.scala 94:16:@25009.4]
  assign x252_div_1_clock = clock; // @[:@25021.4]
  assign x252_div_1_reset = reset; // @[:@25022.4]
  assign x252_div_1_io_a = x247_rdcol_1_io_result; // @[Math.scala 328:17:@25023.4]
  assign x252_div_1_io_flow = io_in_x206_TREADY; // @[Math.scala 330:20:@25025.4]
  assign RetimeWrapper_32_clock = clock; // @[:@25031.4]
  assign RetimeWrapper_32_reset = reset; // @[:@25032.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25034.4]
  assign RetimeWrapper_32_io_in = x252_div_1_io_result; // @[package.scala 94:16:@25033.4]
  assign x253_sum_1_clock = clock; // @[:@25042.4]
  assign x253_sum_1_reset = reset; // @[:@25043.4]
  assign x253_sum_1_io_a = x243_mul_1_io_result; // @[Math.scala 151:17:@25044.4]
  assign x253_sum_1_io_b = RetimeWrapper_32_io_out; // @[Math.scala 152:17:@25045.4]
  assign x253_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25046.4]
  assign RetimeWrapper_33_clock = clock; // @[:@25052.4]
  assign RetimeWrapper_33_reset = reset; // @[:@25053.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25055.4]
  assign RetimeWrapper_33_io_in = x253_sum_1_io_result; // @[package.scala 94:16:@25054.4]
  assign RetimeWrapper_34_clock = clock; // @[:@25061.4]
  assign RetimeWrapper_34_reset = reset; // @[:@25062.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25064.4]
  assign RetimeWrapper_34_io_in = x436 ? x484_x435_sum_D1_number : x438_sub_number; // @[package.scala 94:16:@25063.4]
  assign RetimeWrapper_35_clock = clock; // @[:@25070.4]
  assign RetimeWrapper_35_reset = reset; // @[:@25071.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25073.4]
  assign RetimeWrapper_35_io_in = ~ x249; // @[package.scala 94:16:@25072.4]
  assign RetimeWrapper_36_clock = clock; // @[:@25082.4]
  assign RetimeWrapper_36_reset = reset; // @[:@25083.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25085.4]
  assign RetimeWrapper_36_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25084.4]
  assign x256_rdcol_1_clock = clock; // @[:@25105.4]
  assign x256_rdcol_1_reset = reset; // @[:@25106.4]
  assign x256_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@25107.4]
  assign x256_rdcol_1_io_b = 32'h2; // @[Math.scala 193:17:@25108.4]
  assign x256_rdcol_1_io_flow = io_in_x206_TREADY; // @[Math.scala 194:20:@25109.4]
  assign RetimeWrapper_37_clock = clock; // @[:@25120.4]
  assign RetimeWrapper_37_reset = reset; // @[:@25121.4]
  assign RetimeWrapper_37_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@25123.4]
  assign RetimeWrapper_37_io_in = $signed(_T_937) < $signed(32'sh0); // @[package.scala 94:16:@25122.4]
  assign x442_sum_1_clock = clock; // @[:@25155.4]
  assign x442_sum_1_reset = reset; // @[:@25156.4]
  assign x442_sum_1_io_a = {_T_953,_T_954}; // @[Math.scala 151:17:@25157.4]
  assign x442_sum_1_io_b = $unsigned(_T_966); // @[Math.scala 152:17:@25158.4]
  assign x442_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25159.4]
  assign RetimeWrapper_38_clock = clock; // @[:@25171.4]
  assign RetimeWrapper_38_reset = reset; // @[:@25172.4]
  assign RetimeWrapper_38_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@25174.4]
  assign RetimeWrapper_38_io_in = {_T_978,_T_979}; // @[package.scala 94:16:@25173.4]
  assign RetimeWrapper_39_clock = clock; // @[:@25188.4]
  assign RetimeWrapper_39_reset = reset; // @[:@25189.4]
  assign RetimeWrapper_39_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@25192.4]
  assign RetimeWrapper_39_io_in = $unsigned(_T_993); // @[package.scala 94:16:@25191.4]
  assign x445_sum_1_clock = clock; // @[:@25201.4]
  assign x445_sum_1_reset = reset; // @[:@25202.4]
  assign x445_sum_1_io_a = RetimeWrapper_38_io_out; // @[Math.scala 151:17:@25203.4]
  assign x445_sum_1_io_b = $unsigned(_T_997); // @[Math.scala 152:17:@25204.4]
  assign x445_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25205.4]
  assign x448_sum_1_clock = clock; // @[:@25231.4]
  assign x448_sum_1_reset = reset; // @[:@25232.4]
  assign x448_sum_1_io_a = {_T_1009,_T_1010}; // @[Math.scala 151:17:@25233.4]
  assign x448_sum_1_io_b = $unsigned(_T_1022); // @[Math.scala 152:17:@25234.4]
  assign x448_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25235.4]
  assign x451_sum_1_clock = clock; // @[:@25261.4]
  assign x451_sum_1_reset = reset; // @[:@25262.4]
  assign x451_sum_1_io_a = {_T_1034,_T_1035}; // @[Math.scala 151:17:@25263.4]
  assign x451_sum_1_io_b = $unsigned(_T_1047); // @[Math.scala 152:17:@25264.4]
  assign x451_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25265.4]
  assign x454_sum_1_clock = clock; // @[:@25291.4]
  assign x454_sum_1_reset = reset; // @[:@25292.4]
  assign x454_sum_1_io_a = {_T_1059,_T_1060}; // @[Math.scala 151:17:@25293.4]
  assign x454_sum_1_io_b = $unsigned(_T_1072); // @[Math.scala 152:17:@25294.4]
  assign x454_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25295.4]
  assign x457_sum_1_clock = clock; // @[:@25321.4]
  assign x457_sum_1_reset = reset; // @[:@25322.4]
  assign x457_sum_1_io_a = {_T_1084,_T_1085}; // @[Math.scala 151:17:@25323.4]
  assign x457_sum_1_io_b = $unsigned(_T_1097); // @[Math.scala 152:17:@25324.4]
  assign x457_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25325.4]
  assign RetimeWrapper_40_clock = clock; // @[:@25336.4]
  assign RetimeWrapper_40_reset = reset; // @[:@25337.4]
  assign RetimeWrapper_40_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@25339.4]
  assign RetimeWrapper_40_io_in = $signed(_T_1107) < $signed(32'sh3); // @[package.scala 94:16:@25338.4]
  assign RetimeWrapper_41_clock = clock; // @[:@25350.4]
  assign RetimeWrapper_41_reset = reset; // @[:@25351.4]
  assign RetimeWrapper_41_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@25353.4]
  assign RetimeWrapper_41_io_in = $signed(_T_1107) < $signed(32'sh6); // @[package.scala 94:16:@25352.4]
  assign x460_sub_1_clock = clock; // @[:@25361.4]
  assign x460_sub_1_reset = reset; // @[:@25362.4]
  assign x460_sub_1_io_a = x457_sum_1_io_result; // @[Math.scala 192:17:@25363.4]
  assign x460_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@25364.4]
  assign x460_sub_1_io_flow = io_in_x206_TREADY; // @[Math.scala 194:20:@25365.4]
  assign RetimeWrapper_42_clock = clock; // @[:@25371.4]
  assign RetimeWrapper_42_reset = reset; // @[:@25372.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25374.4]
  assign RetimeWrapper_42_io_in = x457_sum_1_io_result; // @[package.scala 94:16:@25373.4]
  assign x261_div_1_clock = clock; // @[:@25385.4]
  assign x261_div_1_reset = reset; // @[:@25386.4]
  assign x261_div_1_io_a = x256_rdcol_1_io_result; // @[Math.scala 328:17:@25387.4]
  assign x261_div_1_io_flow = io_in_x206_TREADY; // @[Math.scala 330:20:@25389.4]
  assign RetimeWrapper_43_clock = clock; // @[:@25395.4]
  assign RetimeWrapper_43_reset = reset; // @[:@25396.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25398.4]
  assign RetimeWrapper_43_io_in = x261_div_1_io_result; // @[package.scala 94:16:@25397.4]
  assign x262_sum_1_clock = clock; // @[:@25404.4]
  assign x262_sum_1_reset = reset; // @[:@25405.4]
  assign x262_sum_1_io_a = x243_mul_1_io_result; // @[Math.scala 151:17:@25406.4]
  assign x262_sum_1_io_b = RetimeWrapper_43_io_out; // @[Math.scala 152:17:@25407.4]
  assign x262_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25408.4]
  assign RetimeWrapper_44_clock = clock; // @[:@25414.4]
  assign RetimeWrapper_44_reset = reset; // @[:@25415.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25417.4]
  assign RetimeWrapper_44_io_in = x458 ? x489_x457_sum_D1_number : x460_sub_number; // @[package.scala 94:16:@25416.4]
  assign RetimeWrapper_45_clock = clock; // @[:@25423.4]
  assign RetimeWrapper_45_reset = reset; // @[:@25424.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25426.4]
  assign RetimeWrapper_45_io_in = ~ x258; // @[package.scala 94:16:@25425.4]
  assign RetimeWrapper_46_clock = clock; // @[:@25432.4]
  assign RetimeWrapper_46_reset = reset; // @[:@25433.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25435.4]
  assign RetimeWrapper_46_io_in = x262_sum_1_io_result; // @[package.scala 94:16:@25434.4]
  assign RetimeWrapper_47_clock = clock; // @[:@25444.4]
  assign RetimeWrapper_47_reset = reset; // @[:@25445.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25447.4]
  assign RetimeWrapper_47_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25446.4]
  assign x265_rdrow_1_clock = clock; // @[:@25467.4]
  assign x265_rdrow_1_reset = reset; // @[:@25468.4]
  assign x265_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@25469.4]
  assign x265_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@25470.4]
  assign x265_rdrow_1_io_flow = io_in_x206_TREADY; // @[Math.scala 194:20:@25471.4]
  assign x266_1_clock = clock; // @[:@25479.4]
  assign x266_1_reset = reset; // @[:@25480.4]
  assign x266_1_io_a = x265_rdrow_1_io_result; // @[Math.scala 367:17:@25481.4]
  assign x266_1_io_flow = io_in_x206_TREADY; // @[Math.scala 369:20:@25483.4]
  assign RetimeWrapper_48_clock = clock; // @[:@25494.4]
  assign RetimeWrapper_48_reset = reset; // @[:@25495.4]
  assign RetimeWrapper_48_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@25497.4]
  assign RetimeWrapper_48_io_in = $signed(_T_1194) < $signed(32'sh0); // @[package.scala 94:16:@25496.4]
  assign RetimeWrapper_49_clock = clock; // @[:@25503.4]
  assign RetimeWrapper_49_reset = reset; // @[:@25504.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25506.4]
  assign RetimeWrapper_49_io_in = RetimeWrapper_16_io_out; // @[package.scala 94:16:@25505.4]
  assign x272_mul_1_clock = clock; // @[:@25542.4]
  assign x272_mul_1_reset = reset; // @[:@25543.4]
  assign x272_mul_1_io_a = {_T_1225,_T_1226}; // @[Math.scala 263:17:@25544.4]
  assign x272_mul_1_io_flow = io_in_x206_TREADY; // @[Math.scala 265:20:@25546.4]
  assign RetimeWrapper_50_clock = clock; // @[:@25552.4]
  assign RetimeWrapper_50_reset = reset; // @[:@25553.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25555.4]
  assign RetimeWrapper_50_io_in = x232_div_1_io_result; // @[package.scala 94:16:@25554.4]
  assign x273_sum_1_clock = clock; // @[:@25561.4]
  assign x273_sum_1_reset = reset; // @[:@25562.4]
  assign x273_sum_1_io_a = x272_mul_1_io_result; // @[Math.scala 151:17:@25563.4]
  assign x273_sum_1_io_b = RetimeWrapper_50_io_out; // @[Math.scala 152:17:@25564.4]
  assign x273_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25565.4]
  assign RetimeWrapper_51_clock = clock; // @[:@25571.4]
  assign RetimeWrapper_51_reset = reset; // @[:@25572.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25574.4]
  assign RetimeWrapper_51_io_in = ~ x268; // @[package.scala 94:16:@25573.4]
  assign RetimeWrapper_52_clock = clock; // @[:@25580.4]
  assign RetimeWrapper_52_reset = reset; // @[:@25581.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25583.4]
  assign RetimeWrapper_52_io_in = $unsigned(_T_1216); // @[package.scala 94:16:@25582.4]
  assign RetimeWrapper_53_clock = clock; // @[:@25589.4]
  assign RetimeWrapper_53_reset = reset; // @[:@25590.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25592.4]
  assign RetimeWrapper_53_io_in = x273_sum_1_io_result; // @[package.scala 94:16:@25591.4]
  assign RetimeWrapper_54_clock = clock; // @[:@25601.4]
  assign RetimeWrapper_54_reset = reset; // @[:@25602.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25604.4]
  assign RetimeWrapper_54_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25603.4]
  assign RetimeWrapper_55_clock = clock; // @[:@25628.4]
  assign RetimeWrapper_55_reset = reset; // @[:@25629.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25631.4]
  assign RetimeWrapper_55_io_in = x252_div_1_io_result; // @[package.scala 94:16:@25630.4]
  assign x278_sum_1_clock = clock; // @[:@25637.4]
  assign x278_sum_1_reset = reset; // @[:@25638.4]
  assign x278_sum_1_io_a = x272_mul_1_io_result; // @[Math.scala 151:17:@25639.4]
  assign x278_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@25640.4]
  assign x278_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25641.4]
  assign RetimeWrapper_56_clock = clock; // @[:@25647.4]
  assign RetimeWrapper_56_reset = reset; // @[:@25648.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25650.4]
  assign RetimeWrapper_56_io_in = x278_sum_1_io_result; // @[package.scala 94:16:@25649.4]
  assign RetimeWrapper_57_clock = clock; // @[:@25656.4]
  assign RetimeWrapper_57_reset = reset; // @[:@25657.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25659.4]
  assign RetimeWrapper_57_io_in = ~ x276; // @[package.scala 94:16:@25658.4]
  assign RetimeWrapper_58_clock = clock; // @[:@25668.4]
  assign RetimeWrapper_58_reset = reset; // @[:@25669.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25671.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25670.4]
  assign RetimeWrapper_59_clock = clock; // @[:@25695.4]
  assign RetimeWrapper_59_reset = reset; // @[:@25696.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25698.4]
  assign RetimeWrapper_59_io_in = x261_div_1_io_result; // @[package.scala 94:16:@25697.4]
  assign x283_sum_1_clock = clock; // @[:@25704.4]
  assign x283_sum_1_reset = reset; // @[:@25705.4]
  assign x283_sum_1_io_a = x272_mul_1_io_result; // @[Math.scala 151:17:@25706.4]
  assign x283_sum_1_io_b = RetimeWrapper_59_io_out; // @[Math.scala 152:17:@25707.4]
  assign x283_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25708.4]
  assign RetimeWrapper_60_clock = clock; // @[:@25714.4]
  assign RetimeWrapper_60_reset = reset; // @[:@25715.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25717.4]
  assign RetimeWrapper_60_io_in = ~ x281; // @[package.scala 94:16:@25716.4]
  assign RetimeWrapper_61_clock = clock; // @[:@25723.4]
  assign RetimeWrapper_61_reset = reset; // @[:@25724.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25726.4]
  assign RetimeWrapper_61_io_in = x283_sum_1_io_result; // @[package.scala 94:16:@25725.4]
  assign RetimeWrapper_62_clock = clock; // @[:@25735.4]
  assign RetimeWrapper_62_reset = reset; // @[:@25736.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25738.4]
  assign RetimeWrapper_62_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25737.4]
  assign x286_rdrow_1_clock = clock; // @[:@25758.4]
  assign x286_rdrow_1_reset = reset; // @[:@25759.4]
  assign x286_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@25760.4]
  assign x286_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@25761.4]
  assign x286_rdrow_1_io_flow = io_in_x206_TREADY; // @[Math.scala 194:20:@25762.4]
  assign x287_1_clock = clock; // @[:@25770.4]
  assign x287_1_reset = reset; // @[:@25771.4]
  assign x287_1_io_a = x286_rdrow_1_io_result; // @[Math.scala 367:17:@25772.4]
  assign x287_1_io_flow = io_in_x206_TREADY; // @[Math.scala 369:20:@25774.4]
  assign RetimeWrapper_63_clock = clock; // @[:@25785.4]
  assign RetimeWrapper_63_reset = reset; // @[:@25786.4]
  assign RetimeWrapper_63_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@25788.4]
  assign RetimeWrapper_63_io_in = $signed(_T_1360) < $signed(32'sh0); // @[package.scala 94:16:@25787.4]
  assign x293_mul_1_clock = clock; // @[:@25822.4]
  assign x293_mul_1_reset = reset; // @[:@25823.4]
  assign x293_mul_1_io_a = {_T_1388,_T_1389}; // @[Math.scala 263:17:@25824.4]
  assign x293_mul_1_io_flow = io_in_x206_TREADY; // @[Math.scala 265:20:@25826.4]
  assign x294_sum_1_clock = clock; // @[:@25832.4]
  assign x294_sum_1_reset = reset; // @[:@25833.4]
  assign x294_sum_1_io_a = x293_mul_1_io_result; // @[Math.scala 151:17:@25834.4]
  assign x294_sum_1_io_b = RetimeWrapper_50_io_out; // @[Math.scala 152:17:@25835.4]
  assign x294_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25836.4]
  assign RetimeWrapper_64_clock = clock; // @[:@25842.4]
  assign RetimeWrapper_64_reset = reset; // @[:@25843.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25845.4]
  assign RetimeWrapper_64_io_in = $unsigned(_T_1379); // @[package.scala 94:16:@25844.4]
  assign RetimeWrapper_65_clock = clock; // @[:@25851.4]
  assign RetimeWrapper_65_reset = reset; // @[:@25852.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25854.4]
  assign RetimeWrapper_65_io_in = ~ x289; // @[package.scala 94:16:@25853.4]
  assign RetimeWrapper_66_clock = clock; // @[:@25860.4]
  assign RetimeWrapper_66_reset = reset; // @[:@25861.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25863.4]
  assign RetimeWrapper_66_io_in = x294_sum_1_io_result; // @[package.scala 94:16:@25862.4]
  assign RetimeWrapper_67_clock = clock; // @[:@25872.4]
  assign RetimeWrapper_67_reset = reset; // @[:@25873.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25875.4]
  assign RetimeWrapper_67_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25874.4]
  assign x299_sum_1_clock = clock; // @[:@25899.4]
  assign x299_sum_1_reset = reset; // @[:@25900.4]
  assign x299_sum_1_io_a = x293_mul_1_io_result; // @[Math.scala 151:17:@25901.4]
  assign x299_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@25902.4]
  assign x299_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25903.4]
  assign RetimeWrapper_68_clock = clock; // @[:@25909.4]
  assign RetimeWrapper_68_reset = reset; // @[:@25910.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25912.4]
  assign RetimeWrapper_68_io_in = ~ x297; // @[package.scala 94:16:@25911.4]
  assign RetimeWrapper_69_clock = clock; // @[:@25918.4]
  assign RetimeWrapper_69_reset = reset; // @[:@25919.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25921.4]
  assign RetimeWrapper_69_io_in = x299_sum_1_io_result; // @[package.scala 94:16:@25920.4]
  assign RetimeWrapper_70_clock = clock; // @[:@25930.4]
  assign RetimeWrapper_70_reset = reset; // @[:@25931.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25933.4]
  assign RetimeWrapper_70_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25932.4]
  assign x304_sum_1_clock = clock; // @[:@25957.4]
  assign x304_sum_1_reset = reset; // @[:@25958.4]
  assign x304_sum_1_io_a = x293_mul_1_io_result; // @[Math.scala 151:17:@25959.4]
  assign x304_sum_1_io_b = RetimeWrapper_59_io_out; // @[Math.scala 152:17:@25960.4]
  assign x304_sum_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@25961.4]
  assign RetimeWrapper_71_clock = clock; // @[:@25967.4]
  assign RetimeWrapper_71_reset = reset; // @[:@25968.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25970.4]
  assign RetimeWrapper_71_io_in = ~ x302; // @[package.scala 94:16:@25969.4]
  assign RetimeWrapper_72_clock = clock; // @[:@25976.4]
  assign RetimeWrapper_72_reset = reset; // @[:@25977.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25979.4]
  assign RetimeWrapper_72_io_in = x304_sum_1_io_result; // @[package.scala 94:16:@25978.4]
  assign RetimeWrapper_73_clock = clock; // @[:@25988.4]
  assign RetimeWrapper_73_reset = reset; // @[:@25989.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25991.4]
  assign RetimeWrapper_73_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25990.4]
  assign x312_x11_1_clock = clock; // @[:@26036.4]
  assign x312_x11_1_reset = reset; // @[:@26037.4]
  assign x312_x11_1_io_a = x218_lb_0_io_rPort_3_output_0; // @[Math.scala 151:17:@26038.4]
  assign x312_x11_1_io_b = _T_1498[7:0]; // @[Math.scala 152:17:@26039.4]
  assign x312_x11_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@26040.4]
  assign x313_x12_1_clock = clock; // @[:@26046.4]
  assign x313_x12_1_reset = reset; // @[:@26047.4]
  assign x313_x12_1_io_a = x218_lb_0_io_rPort_5_output_0; // @[Math.scala 151:17:@26048.4]
  assign x313_x12_1_io_b = _T_1502[7:0]; // @[Math.scala 152:17:@26049.4]
  assign x313_x12_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@26050.4]
  assign x314_x11_1_clock = clock; // @[:@26056.4]
  assign x314_x11_1_reset = reset; // @[:@26057.4]
  assign x314_x11_1_io_a = _T_1506[7:0]; // @[Math.scala 151:17:@26058.4]
  assign x314_x11_1_io_b = _T_1510[7:0]; // @[Math.scala 152:17:@26059.4]
  assign x314_x11_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@26060.4]
  assign x315_x12_1_clock = clock; // @[:@26066.4]
  assign x315_x12_1_reset = reset; // @[:@26067.4]
  assign x315_x12_1_io_a = x218_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@26068.4]
  assign x315_x12_1_io_b = _T_1514[7:0]; // @[Math.scala 152:17:@26069.4]
  assign x315_x12_1_io_flow = io_in_x206_TREADY; // @[Math.scala 153:20:@26070.4]
  assign x316_x11_1_io_a = x312_x11_1_io_result; // @[Math.scala 151:17:@26078.4]
  assign x316_x11_1_io_b = x313_x12_1_io_result; // @[Math.scala 152:17:@26079.4]
  assign x317_x12_1_io_a = x314_x11_1_io_result; // @[Math.scala 151:17:@26088.4]
  assign x317_x12_1_io_b = x315_x12_1_io_result; // @[Math.scala 152:17:@26089.4]
  assign x318_x11_1_io_a = x316_x11_1_io_result; // @[Math.scala 151:17:@26098.4]
  assign x318_x11_1_io_b = x317_x12_1_io_result; // @[Math.scala 152:17:@26099.4]
  assign RetimeWrapper_74_clock = clock; // @[:@26106.4]
  assign RetimeWrapper_74_reset = reset; // @[:@26107.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26109.4]
  assign RetimeWrapper_74_io_in = x218_lb_0_io_rPort_7_output_0; // @[package.scala 94:16:@26108.4]
  assign x319_sum_1_io_a = x318_x11_1_io_result; // @[Math.scala 151:17:@26117.4]
  assign x319_sum_1_io_b = RetimeWrapper_74_io_out; // @[Math.scala 152:17:@26118.4]
  assign RetimeWrapper_75_clock = clock; // @[:@26129.4]
  assign RetimeWrapper_75_reset = reset; // @[:@26130.4]
  assign RetimeWrapper_75_io_flow = io_in_x206_TREADY; // @[package.scala 95:18:@26132.4]
  assign RetimeWrapper_75_io_in = {4'h0,_T_1550}; // @[package.scala 94:16:@26131.4]
  assign RetimeWrapper_76_clock = clock; // @[:@26143.4]
  assign RetimeWrapper_76_reset = reset; // @[:@26144.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26146.4]
  assign RetimeWrapper_76_io_in = RetimeWrapper_75_io_out; // @[package.scala 94:16:@26145.4]
  assign RetimeWrapper_77_clock = clock; // @[:@26152.4]
  assign RetimeWrapper_77_reset = reset; // @[:@26153.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26155.4]
  assign RetimeWrapper_77_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@26154.4]
  assign RetimeWrapper_78_clock = clock; // @[:@26161.4]
  assign RetimeWrapper_78_reset = reset; // @[:@26162.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26164.4]
  assign RetimeWrapper_78_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@26163.4]
  assign RetimeWrapper_79_clock = clock; // @[:@26170.4]
  assign RetimeWrapper_79_reset = reset; // @[:@26171.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26173.4]
  assign RetimeWrapper_79_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26172.4]
endmodule
module x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1( // @[:@26191.2]
  input          clock, // @[:@26192.4]
  input          reset, // @[:@26193.4]
  output         io_in_x206_TVALID, // @[:@26194.4]
  input          io_in_x206_TREADY, // @[:@26194.4]
  output [255:0] io_in_x206_TDATA, // @[:@26194.4]
  input          io_in_x205_TVALID, // @[:@26194.4]
  output         io_in_x205_TREADY, // @[:@26194.4]
  input  [255:0] io_in_x205_TDATA, // @[:@26194.4]
  input  [7:0]   io_in_x205_TID, // @[:@26194.4]
  input  [7:0]   io_in_x205_TDEST, // @[:@26194.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@26194.4]
  input          io_sigsIn_smChildAcks_0, // @[:@26194.4]
  output         io_sigsOut_smDoneIn_0, // @[:@26194.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@26194.4]
  input          io_rr // @[:@26194.4]
);
  wire  x213_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire  x213_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire  x213_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire  x213_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire [31:0] x213_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire [31:0] x213_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire  x213_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire  x213_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire  x213_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@26204.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26292.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26292.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26292.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@26292.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@26292.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@26334.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@26334.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@26334.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@26334.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@26334.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@26342.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@26342.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@26342.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@26342.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@26342.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TVALID; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TREADY; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire [255:0] x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TDATA; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TREADY; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire [255:0] x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TDATA; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire [7:0] x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TID; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire [7:0] x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TDEST; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire [31:0] x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire [31:0] x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
  wire  _T_239; // @[package.scala 96:25:@26297.4 package.scala 96:25:@26298.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x326_outr_UnitPipe.scala 68:66:@26303.4]
  wire  _T_252; // @[package.scala 96:25:@26339.4 package.scala 96:25:@26340.4]
  wire  _T_258; // @[package.scala 96:25:@26347.4 package.scala 96:25:@26348.4]
  wire  _T_261; // @[SpatialBlocks.scala 138:93:@26350.4]
  wire  x325_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@26351.4]
  wire  _T_263; // @[SpatialBlocks.scala 157:36:@26359.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:78:@26360.4]
  wire  _T_271; // @[SpatialBlocks.scala 159:58:@26372.4]
  x213_ctrchain x213_ctrchain ( // @[SpatialBlocks.scala 37:22:@26204.4]
    .clock(x213_ctrchain_clock),
    .reset(x213_ctrchain_reset),
    .io_input_reset(x213_ctrchain_io_input_reset),
    .io_input_enable(x213_ctrchain_io_input_enable),
    .io_output_counts_1(x213_ctrchain_io_output_counts_1),
    .io_output_counts_0(x213_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x213_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x213_ctrchain_io_output_oobs_1),
    .io_output_done(x213_ctrchain_io_output_done)
  );
  x325_inr_Foreach_SAMPLER_BOX_sm x325_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 32:18:@26264.4]
    .clock(x325_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x325_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x325_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x325_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x325_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x325_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x325_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x325_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x325_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@26292.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@26334.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@26342.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1 x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 580:24:@26377.4]
    .clock(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x206_TVALID(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TVALID),
    .io_in_x206_TREADY(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TREADY),
    .io_in_x206_TDATA(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TDATA),
    .io_in_x205_TREADY(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TREADY),
    .io_in_x205_TDATA(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TDATA),
    .io_in_x205_TID(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TID),
    .io_in_x205_TDEST(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TDEST),
    .io_sigsIn_backpressure(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@26297.4 package.scala 96:25:@26298.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x205_TVALID | x325_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x326_outr_UnitPipe.scala 68:66:@26303.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@26339.4 package.scala 96:25:@26340.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@26347.4 package.scala 96:25:@26348.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 138:93:@26350.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 138:90:@26351.4]
  assign _T_263 = x325_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@26359.4]
  assign _T_264 = ~ x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@26360.4]
  assign _T_271 = x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@26372.4]
  assign io_in_x206_TVALID = x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TVALID; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 48:23:@26436.4]
  assign io_in_x206_TDATA = x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TDATA; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 48:23:@26434.4]
  assign io_in_x205_TREADY = x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TREADY; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 49:23:@26444.4]
  assign io_sigsOut_smDoneIn_0 = x325_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@26357.4]
  assign io_sigsOut_smCtrCopyDone_0 = x325_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 168:125:@26376.4]
  assign x213_ctrchain_clock = clock; // @[:@26205.4]
  assign x213_ctrchain_reset = reset; // @[:@26206.4]
  assign x213_ctrchain_io_input_reset = x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@26375.4]
  assign x213_ctrchain_io_input_enable = _T_271 & x325_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@26327.4 SpatialBlocks.scala 159:42:@26374.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@26265.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@26266.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sm_io_enable = x325_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x325_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@26354.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x326_outr_UnitPipe.scala 66:50:@26300.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@26356.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x206_TREADY | x325_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@26328.4]
  assign x325_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x326_outr_UnitPipe.scala 70:48:@26306.4]
  assign RetimeWrapper_clock = clock; // @[:@26293.4]
  assign RetimeWrapper_reset = reset; // @[:@26294.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@26296.4]
  assign RetimeWrapper_io_in = x213_ctrchain_io_output_done; // @[package.scala 94:16:@26295.4]
  assign RetimeWrapper_1_clock = clock; // @[:@26335.4]
  assign RetimeWrapper_1_reset = reset; // @[:@26336.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@26338.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@26337.4]
  assign RetimeWrapper_2_clock = clock; // @[:@26343.4]
  assign RetimeWrapper_2_reset = reset; // @[:@26344.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@26346.4]
  assign RetimeWrapper_2_io_in = x325_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@26345.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@26378.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@26379.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x206_TREADY = io_in_x206_TREADY; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 48:23:@26435.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TDATA = io_in_x205_TDATA; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 49:23:@26443.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TID = io_in_x205_TID; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 49:23:@26439.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x205_TDEST = io_in_x205_TDEST; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 49:23:@26438.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x206_TREADY | x325_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 585:22:@26462.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 585:22:@26460.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x325_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 585:22:@26458.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x213_ctrchain_io_output_counts_1; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 585:22:@26453.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x213_ctrchain_io_output_counts_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 585:22:@26452.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x213_ctrchain_io_output_oobs_0; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 585:22:@26450.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x213_ctrchain_io_output_oobs_1; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 585:22:@26451.4]
  assign x325_inr_Foreach_SAMPLER_BOX_kernelx325_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x325_inr_Foreach_SAMPLER_BOX.scala 584:18:@26446.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@26476.2]
  input          clock, // @[:@26477.4]
  input          reset, // @[:@26478.4]
  output         io_in_x206_TVALID, // @[:@26479.4]
  input          io_in_x206_TREADY, // @[:@26479.4]
  output [255:0] io_in_x206_TDATA, // @[:@26479.4]
  input          io_in_x205_TVALID, // @[:@26479.4]
  output         io_in_x205_TREADY, // @[:@26479.4]
  input  [255:0] io_in_x205_TDATA, // @[:@26479.4]
  input  [7:0]   io_in_x205_TID, // @[:@26479.4]
  input  [7:0]   io_in_x205_TDEST, // @[:@26479.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@26479.4]
  input          io_sigsIn_smChildAcks_0, // @[:@26479.4]
  output         io_sigsOut_smDoneIn_0, // @[:@26479.4]
  input          io_rr // @[:@26479.4]
);
  wire  x326_outr_UnitPipe_sm_clock; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_reset; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_io_enable; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_io_done; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_io_parentAck; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_io_childAck_0; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  x326_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26673.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26673.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26673.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@26673.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@26673.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@26681.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@26681.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@26681.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@26681.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@26681.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_clock; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_reset; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TVALID; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TREADY; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire [255:0] x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TDATA; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TVALID; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TREADY; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire [255:0] x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TDATA; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire [7:0] x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TID; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire [7:0] x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TDEST; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_rr; // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
  wire  _T_246; // @[package.scala 96:25:@26678.4 package.scala 96:25:@26679.4]
  wire  _T_252; // @[package.scala 96:25:@26686.4 package.scala 96:25:@26687.4]
  wire  _T_255; // @[SpatialBlocks.scala 138:93:@26689.4]
  x326_outr_UnitPipe_sm x326_outr_UnitPipe_sm ( // @[sm_x326_outr_UnitPipe.scala 32:18:@26621.4]
    .clock(x326_outr_UnitPipe_sm_clock),
    .reset(x326_outr_UnitPipe_sm_reset),
    .io_enable(x326_outr_UnitPipe_sm_io_enable),
    .io_done(x326_outr_UnitPipe_sm_io_done),
    .io_parentAck(x326_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x326_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x326_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x326_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x326_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@26673.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@26681.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1 x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1 ( // @[sm_x326_outr_UnitPipe.scala 75:24:@26711.4]
    .clock(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_clock),
    .reset(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_reset),
    .io_in_x206_TVALID(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TVALID),
    .io_in_x206_TREADY(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TREADY),
    .io_in_x206_TDATA(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TDATA),
    .io_in_x205_TVALID(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TVALID),
    .io_in_x205_TREADY(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TREADY),
    .io_in_x205_TDATA(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TDATA),
    .io_in_x205_TID(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TID),
    .io_in_x205_TDEST(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TDEST),
    .io_sigsIn_smEnableOuts_0(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@26678.4 package.scala 96:25:@26679.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@26686.4 package.scala 96:25:@26687.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 138:93:@26689.4]
  assign io_in_x206_TVALID = x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TVALID; // @[sm_x326_outr_UnitPipe.scala 48:23:@26768.4]
  assign io_in_x206_TDATA = x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TDATA; // @[sm_x326_outr_UnitPipe.scala 48:23:@26766.4]
  assign io_in_x205_TREADY = x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TREADY; // @[sm_x326_outr_UnitPipe.scala 49:23:@26776.4]
  assign io_sigsOut_smDoneIn_0 = x326_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@26696.4]
  assign x326_outr_UnitPipe_sm_clock = clock; // @[:@26622.4]
  assign x326_outr_UnitPipe_sm_reset = reset; // @[:@26623.4]
  assign x326_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 140:18:@26693.4]
  assign x326_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@26695.4]
  assign x326_outr_UnitPipe_sm_io_doneIn_0 = x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@26665.4]
  assign x326_outr_UnitPipe_sm_io_ctrCopyDone_0 = x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@26710.4]
  assign RetimeWrapper_clock = clock; // @[:@26674.4]
  assign RetimeWrapper_reset = reset; // @[:@26675.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@26677.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@26676.4]
  assign RetimeWrapper_1_clock = clock; // @[:@26682.4]
  assign RetimeWrapper_1_reset = reset; // @[:@26683.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@26685.4]
  assign RetimeWrapper_1_io_in = x326_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@26684.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_clock = clock; // @[:@26712.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_reset = reset; // @[:@26713.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x206_TREADY = io_in_x206_TREADY; // @[sm_x326_outr_UnitPipe.scala 48:23:@26767.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TVALID = io_in_x205_TVALID; // @[sm_x326_outr_UnitPipe.scala 49:23:@26777.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TDATA = io_in_x205_TDATA; // @[sm_x326_outr_UnitPipe.scala 49:23:@26775.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TID = io_in_x205_TID; // @[sm_x326_outr_UnitPipe.scala 49:23:@26771.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_in_x205_TDEST = io_in_x205_TDEST; // @[sm_x326_outr_UnitPipe.scala 49:23:@26770.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x326_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x326_outr_UnitPipe.scala 80:22:@26786.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x326_outr_UnitPipe_sm_io_childAck_0; // @[sm_x326_outr_UnitPipe.scala 80:22:@26784.4]
  assign x326_outr_UnitPipe_kernelx326_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x326_outr_UnitPipe.scala 79:18:@26778.4]
endmodule
module AccelUnit( // @[:@26806.2]
  input          clock, // @[:@26807.4]
  input          reset, // @[:@26808.4]
  input          io_enable, // @[:@26809.4]
  output         io_done, // @[:@26809.4]
  input          io_reset, // @[:@26809.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@26809.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@26809.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@26809.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@26809.4]
  output         io_memStreams_loads_0_data_ready, // @[:@26809.4]
  input          io_memStreams_loads_0_data_valid, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@26809.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@26809.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@26809.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@26809.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@26809.4]
  input          io_memStreams_stores_0_data_ready, // @[:@26809.4]
  output         io_memStreams_stores_0_data_valid, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@26809.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@26809.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@26809.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@26809.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@26809.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@26809.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@26809.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@26809.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@26809.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@26809.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@26809.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@26809.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@26809.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@26809.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@26809.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@26809.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@26809.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@26809.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@26809.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@26809.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@26809.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@26809.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@26809.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@26809.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@26809.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@26809.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@26809.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@26809.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@26809.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@26809.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@26809.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@26809.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@26809.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@26809.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@26809.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@26809.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@26809.4]
  output         io_heap_0_req_valid, // @[:@26809.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@26809.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@26809.4]
  input          io_heap_0_resp_valid, // @[:@26809.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@26809.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@26809.4]
  input  [63:0]  io_argIns_0, // @[:@26809.4]
  input  [63:0]  io_argIns_1, // @[:@26809.4]
  input          io_argOuts_0_port_ready, // @[:@26809.4]
  output         io_argOuts_0_port_valid, // @[:@26809.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@26809.4]
  input  [63:0]  io_argOuts_0_echo // @[:@26809.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@26972.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@26972.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@26972.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@26972.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26990.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26990.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26990.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@26990.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@26990.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@26999.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@26999.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@26999.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@26999.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@26999.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@26999.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@27038.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27070.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27070.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27070.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@27070.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@27070.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_in_x206_TVALID; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_in_x206_TREADY; // @[sm_RootController.scala 73:24:@27132.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x206_TDATA; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_in_x205_TVALID; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_in_x205_TREADY; // @[sm_RootController.scala 73:24:@27132.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x205_TDATA; // @[sm_RootController.scala 73:24:@27132.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x205_TID; // @[sm_RootController.scala 73:24:@27132.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x205_TDEST; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@27132.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@27132.4]
  wire  _T_599; // @[package.scala 96:25:@26995.4 package.scala 96:25:@26996.4]
  wire  _T_664; // @[Main.scala 41:50:@27066.4]
  wire  _T_665; // @[Main.scala 41:59:@27067.4]
  wire  _T_677; // @[package.scala 100:49:@27087.4]
  reg  _T_680; // @[package.scala 48:56:@27088.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@26972.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@26990.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@26999.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@27038.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@27070.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@27132.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x206_TVALID(RootController_kernelRootController_concrete1_io_in_x206_TVALID),
    .io_in_x206_TREADY(RootController_kernelRootController_concrete1_io_in_x206_TREADY),
    .io_in_x206_TDATA(RootController_kernelRootController_concrete1_io_in_x206_TDATA),
    .io_in_x205_TVALID(RootController_kernelRootController_concrete1_io_in_x205_TVALID),
    .io_in_x205_TREADY(RootController_kernelRootController_concrete1_io_in_x205_TREADY),
    .io_in_x205_TDATA(RootController_kernelRootController_concrete1_io_in_x205_TDATA),
    .io_in_x205_TID(RootController_kernelRootController_concrete1_io_in_x205_TID),
    .io_in_x205_TDEST(RootController_kernelRootController_concrete1_io_in_x205_TDEST),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@26995.4 package.scala 96:25:@26996.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@27066.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@27067.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@27087.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@27086.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x205_TREADY; // @[sm_RootController.scala 49:23:@27197.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x206_TVALID; // @[sm_RootController.scala 48:23:@27189.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x206_TDATA; // @[sm_RootController.scala 48:23:@27187.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 48:23:@27186.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 48:23:@27185.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 48:23:@27184.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 48:23:@27183.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 48:23:@27182.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 48:23:@27181.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@26973.4]
  assign SingleCounter_reset = reset; // @[:@26974.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@26988.4]
  assign RetimeWrapper_clock = clock; // @[:@26991.4]
  assign RetimeWrapper_reset = reset; // @[:@26992.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@26994.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@26993.4]
  assign SRFF_clock = clock; // @[:@27000.4]
  assign SRFF_reset = reset; // @[:@27001.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@27226.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@27084.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@27085.4]
  assign RootController_sm_clock = clock; // @[:@27039.4]
  assign RootController_sm_reset = reset; // @[:@27040.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@27083.4 SpatialBlocks.scala 140:18:@27117.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@27111.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@27091.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@27108.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27071.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27072.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@27074.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@27073.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@27133.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@27134.4]
  assign RootController_kernelRootController_concrete1_io_in_x206_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 48:23:@27188.4]
  assign RootController_kernelRootController_concrete1_io_in_x205_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 49:23:@27198.4]
  assign RootController_kernelRootController_concrete1_io_in_x205_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 49:23:@27196.4]
  assign RootController_kernelRootController_concrete1_io_in_x205_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 49:23:@27192.4]
  assign RootController_kernelRootController_concrete1_io_in_x205_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 49:23:@27191.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 78:22:@27207.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 78:22:@27205.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 77:18:@27199.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@27228.2]
  input         clock, // @[:@27229.4]
  input         reset, // @[:@27230.4]
  input  [31:0] io_raddr, // @[:@27231.4]
  input         io_wen, // @[:@27231.4]
  input  [31:0] io_waddr, // @[:@27231.4]
  input  [63:0] io_wdata, // @[:@27231.4]
  output [63:0] io_rdata // @[:@27231.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@27233.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@27233.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@27233.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@27233.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@27233.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@27233.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@27233.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@27233.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@27233.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@27233.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@27233.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@27233.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@27234.4]
  assign accel_reset = reset; // @[:@27235.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
