// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x244_TREADY(dontcare), // @[:@1298.4]
    .io_in_x244_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x244_TID(8'h0),
    .io_in_x244_TDEST(8'h0),
    .io_in_x245_TVALID(valid_down), // @[:@1298.4]
    .io_in_x245_TDATA({O_0_0_0,O_1_0_0}), // @[:@1298.4]
    .io_in_x245_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x252_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh22); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh22); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 284:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x401_outr_UnitPipe_sm( // @[:@2390.2]
  input   clock, // @[:@2391.4]
  input   reset, // @[:@2392.4]
  input   io_enable, // @[:@2393.4]
  output  io_done, // @[:@2393.4]
  input   io_parentAck, // @[:@2393.4]
  input   io_doneIn_0, // @[:@2393.4]
  output  io_enableOut_0, // @[:@2393.4]
  output  io_childAck_0, // @[:@2393.4]
  input   io_ctrCopyDone_0 // @[:@2393.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2396.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2399.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2416.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2533.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2431.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2432.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2433.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2434.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2435.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2438.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2440.4]
  wire  _T_126; // @[package.scala 96:25:@2452.4 package.scala 96:25:@2453.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2455.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2456.4]
  wire  _T_138; // @[package.scala 96:25:@2466.4 package.scala 96:25:@2467.4]
  wire  _T_156; // @[package.scala 96:25:@2484.4 package.scala 96:25:@2485.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2487.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2488.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2502.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2504.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2506.4]
  reg  _T_186; // @[package.scala 48:56:@2512.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2514.4]
  reg  _T_200; // @[package.scala 48:56:@2530.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2396.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2399.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2416.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2447.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2461.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2479.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2516.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2533.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2431.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2432.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2433.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2434.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2435.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2438.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2440.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2452.4 package.scala 96:25:@2453.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2455.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2456.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2466.4 package.scala 96:25:@2467.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2484.4 package.scala 96:25:@2485.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2487.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2488.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2502.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2504.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2506.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2514.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2540.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2510.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2501.4]
  assign active_0_clock = clock; // @[:@2397.4]
  assign active_0_reset = reset; // @[:@2398.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2442.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2446.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2404.4]
  assign done_0_clock = clock; // @[:@2400.4]
  assign done_0_reset = reset; // @[:@2401.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2492.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2414.4 Controllers.scala 170:32:@2499.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2405.4]
  assign iterDone_0_clock = clock; // @[:@2417.4]
  assign iterDone_0_reset = reset; // @[:@2418.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2460.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2428.4 Controllers.scala 168:36:@2476.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2419.4]
  assign RetimeWrapper_clock = clock; // @[:@2448.4]
  assign RetimeWrapper_reset = reset; // @[:@2449.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2451.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2450.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2462.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2463.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2465.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2464.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2480.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2481.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2483.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2482.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2517.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2518.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2520.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2519.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2534.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2535.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2537.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2536.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2661.2]
  input         clock, // @[:@2662.4]
  input         reset, // @[:@2663.4]
  input         io_input_reset, // @[:@2664.4]
  input         io_input_enable, // @[:@2664.4]
  output [31:0] io_output_count_0, // @[:@2664.4]
  output        io_output_oobs_0, // @[:@2664.4]
  output        io_output_done, // @[:@2664.4]
  output        io_output_saturated // @[:@2664.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@2677.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@2677.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@2677.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@2693.4]
  wire  _T_36; // @[Counter.scala 264:45:@2696.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@2721.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@2722.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@2723.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@2724.4]
  wire  _T_57; // @[Counter.scala 293:18:@2726.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@2734.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@2737.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@2738.4]
  wire  _T_75; // @[Counter.scala 322:102:@2742.4]
  wire  _T_77; // @[Counter.scala 322:130:@2743.4]
  FF bases_0 ( // @[Counter.scala 261:53:@2677.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@2693.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@2696.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@2721.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2722.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2723.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@2724.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh780); // @[Counter.scala 293:18:@2726.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@2734.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@2737.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@2738.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 322:102:@2742.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh780); // @[Counter.scala 322:130:@2743.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@2741.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@2745.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@2747.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh780); // @[Counter.scala 340:25:@2750.4]
  assign bases_0_clock = clock; // @[:@2678.4]
  assign bases_0_reset = reset; // @[:@2679.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:12:@2740.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@2719.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@2720.4]
  assign SRFF_clock = clock; // @[:@2694.4]
  assign SRFF_reset = reset; // @[:@2695.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@2698.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@2700.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@2701.4]
endmodule
module SingleCounter_2( // @[:@2790.2]
  input         clock, // @[:@2791.4]
  input         reset, // @[:@2792.4]
  input         io_setup_saturate, // @[:@2793.4]
  input         io_input_reset, // @[:@2793.4]
  input         io_input_enable, // @[:@2793.4]
  output [12:0] io_output_count_0, // @[:@2793.4]
  output        io_output_oobs_0, // @[:@2793.4]
  output        io_output_done // @[:@2793.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@2806.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@2806.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@2806.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@2822.4]
  wire  _T_36; // @[Counter.scala 264:45:@2825.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@2850.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@2851.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@2852.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@2853.4]
  wire  _T_57; // @[Counter.scala 293:18:@2855.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@2863.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@2865.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@2866.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@2867.4]
  wire  _T_75; // @[Counter.scala 322:102:@2871.4]
  wire  _T_77; // @[Counter.scala 322:130:@2872.4]
  FF bases_0 ( // @[Counter.scala 261:53:@2806.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@2822.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@2825.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@2850.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 291:33:@2851.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 291:33:@2852.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@2853.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh400); // @[Counter.scala 293:18:@2855.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@2863.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 299:85:@2865.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@2866.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@2867.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 322:102:@2871.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh400); // @[Counter.scala 322:130:@2872.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@2870.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@2874.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@2876.4]
  assign bases_0_clock = clock; // @[:@2807.4]
  assign bases_0_reset = reset; // @[:@2808.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:12:@2869.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@2848.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@2849.4]
  assign SRFF_clock = clock; // @[:@2823.4]
  assign SRFF_reset = reset; // @[:@2824.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@2827.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@2829.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@2830.4]
endmodule
module x252_ctrchain( // @[:@2881.2]
  input         clock, // @[:@2882.4]
  input         reset, // @[:@2883.4]
  input         io_input_reset, // @[:@2884.4]
  input         io_input_enable, // @[:@2884.4]
  output [31:0] io_output_counts_1, // @[:@2884.4]
  output [31:0] io_output_counts_0, // @[:@2884.4]
  output        io_output_oobs_0, // @[:@2884.4]
  output        io_output_oobs_1, // @[:@2884.4]
  output        io_output_done // @[:@2884.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@2886.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@2889.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@2889.4]
  wire  isDone; // @[Counter.scala 541:51:@2906.4]
  reg  wasDone; // @[Counter.scala 542:24:@2907.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@2915.4]
  wire  _T_66; // @[Counter.scala 546:80:@2916.4]
  reg  doneLatch; // @[Counter.scala 550:26:@2921.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@2922.4]
  wire  _T_74; // @[Counter.scala 551:19:@2923.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@2886.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@2889.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@2906.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@2915.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@2916.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@2922.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@2923.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@2928.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@2925.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@2927.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@2930.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@2918.4]
  assign ctrs_0_clock = clock; // @[:@2887.4]
  assign ctrs_0_reset = reset; // @[:@2888.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@2895.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@2902.4]
  assign ctrs_1_clock = clock; // @[:@2890.4]
  assign ctrs_1_reset = reset; // @[:@2891.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@2905.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@2899.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@2900.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2970.2]
  input   clock, // @[:@2971.4]
  input   reset, // @[:@2972.4]
  input   io_flow, // @[:@2973.4]
  input   io_in, // @[:@2973.4]
  output  io_out // @[:@2973.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(34)) sr ( // @[RetimeShiftRegister.scala 15:20:@2975.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2988.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2987.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2986.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2985.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2984.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2982.4]
endmodule
module RetimeWrapper_16( // @[:@3098.2]
  input   clock, // @[:@3099.4]
  input   reset, // @[:@3100.4]
  input   io_flow, // @[:@3101.4]
  input   io_in, // @[:@3101.4]
  output  io_out // @[:@3101.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(33)) sr ( // @[RetimeShiftRegister.scala 15:20:@3103.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3116.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3115.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3114.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3113.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3112.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3110.4]
endmodule
module x400_inr_Foreach_SAMPLER_BOX_sm( // @[:@3118.2]
  input   clock, // @[:@3119.4]
  input   reset, // @[:@3120.4]
  input   io_enable, // @[:@3121.4]
  output  io_done, // @[:@3121.4]
  output  io_doneLatch, // @[:@3121.4]
  input   io_ctrDone, // @[:@3121.4]
  output  io_datapathEn, // @[:@3121.4]
  output  io_ctrInc, // @[:@3121.4]
  output  io_ctrRst, // @[:@3121.4]
  input   io_parentAck, // @[:@3121.4]
  input   io_backpressure, // @[:@3121.4]
  input   io_break // @[:@3121.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3123.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3123.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3126.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3126.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3218.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3131.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3132.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3133.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3134.4]
  wire  _T_100; // @[package.scala 100:49:@3151.4]
  reg  _T_103; // @[package.scala 48:56:@3152.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3165.4 package.scala 96:25:@3166.4]
  wire  _T_110; // @[package.scala 100:49:@3167.4]
  reg  _T_113; // @[package.scala 48:56:@3168.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3170.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3175.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3176.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3179.4]
  wire  _T_124; // @[package.scala 96:25:@3187.4 package.scala 96:25:@3188.4]
  wire  _T_126; // @[package.scala 100:49:@3189.4]
  reg  _T_129; // @[package.scala 48:56:@3190.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3212.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3214.4]
  reg  _T_153; // @[package.scala 48:56:@3215.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3223.4 package.scala 96:25:@3224.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3225.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3226.4]
  SRFF active ( // @[Controllers.scala 261:22:@3123.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3126.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3160.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3182.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3194.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3202.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3218.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3131.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3132.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3133.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3134.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3151.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3165.4 package.scala 96:25:@3166.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3167.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3170.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3175.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3176.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3179.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3187.4 package.scala 96:25:@3188.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3189.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3214.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3223.4 package.scala 96:25:@3224.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3225.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3226.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3193.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3228.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3178.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3181.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3173.4]
  assign active_clock = clock; // @[:@3124.4]
  assign active_reset = reset; // @[:@3125.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3136.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3140.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3141.4]
  assign done_clock = clock; // @[:@3127.4]
  assign done_reset = reset; // @[:@3128.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3156.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3149.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3150.4]
  assign RetimeWrapper_clock = clock; // @[:@3161.4]
  assign RetimeWrapper_reset = reset; // @[:@3162.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3164.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3163.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3183.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3184.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3186.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3185.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3195.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3196.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3198.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3197.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3203.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3204.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3206.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3205.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3219.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3220.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3222.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3221.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3335.2]
  input  [31:0] io_a, // @[:@3338.4]
  output [31:0] io_b // @[:@3338.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3351.4]
endmodule
module _( // @[:@3353.2]
  input  [31:0] io_b, // @[:@3356.4]
  output [31:0] io_result // @[:@3356.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3361.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3361.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3361.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3374.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3369.4]
endmodule
module SRAM( // @[:@3433.2]
  input        clock, // @[:@3434.4]
  input  [7:0] io_raddr, // @[:@3436.4]
  input        io_wen, // @[:@3436.4]
  input  [7:0] io_waddr, // @[:@3436.4]
  input  [7:0] io_wdata, // @[:@3436.4]
  output [7:0] io_rdata, // @[:@3436.4]
  input        io_backpressure // @[:@3436.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 143:23:@3438.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 143:23:@3438.4]
  wire [7:0] SRAMVerilogSim_waddr; // @[SRAM.scala 143:23:@3438.4]
  wire [7:0] SRAMVerilogSim_raddr; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 143:23:@3438.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(256), .AWIDTH(8)) SRAMVerilogSim ( // @[SRAM.scala 143:23:@3438.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 153:16:@3458.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 148:20:@3452.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 149:27:@3453.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 146:18:@3450.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 151:22:@3455.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 150:22:@3454.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 147:20:@3451.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 145:20:@3449.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 144:18:@3448.4]
endmodule
module RetimeWrapper_20( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_flow, // @[:@3475.4]
  input  [8:0] io_in, // @[:@3475.4]
  output [8:0] io_out // @[:@3475.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3477.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3490.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3489.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@3488.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3487.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3486.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3484.4]
endmodule
module Mem1D_4( // @[:@3492.2]
  input        clock, // @[:@3493.4]
  input        reset, // @[:@3494.4]
  input  [8:0] io_r_ofs_0, // @[:@3495.4]
  input        io_r_backpressure, // @[:@3495.4]
  input  [8:0] io_w_ofs_0, // @[:@3495.4]
  input  [7:0] io_w_data_0, // @[:@3495.4]
  input        io_w_en_0, // @[:@3495.4]
  output [7:0] io_output // @[:@3495.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_raddr; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_waddr; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_wdata; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3502.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3502.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3502.4]
  wire  wInBound; // @[MemPrimitives.scala 554:32:@3497.4]
  wire [8:0] _T_126; // @[package.scala 96:25:@3507.4 package.scala 96:25:@3508.4]
  SRAM SRAM ( // @[MemPrimitives.scala 567:21:@3499.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_20 RetimeWrapper ( // @[package.scala 93:22:@3502.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h100; // @[MemPrimitives.scala 554:32:@3497.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@3507.4 package.scala 96:25:@3508.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 574:17:@3515.4]
  assign SRAM_clock = clock; // @[:@3500.4]
  assign SRAM_io_raddr = _T_126[7:0]; // @[MemPrimitives.scala 568:37:@3509.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 571:22:@3512.4]
  assign SRAM_io_waddr = io_w_ofs_0[7:0]; // @[MemPrimitives.scala 570:22:@3510.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 572:22:@3513.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 573:30:@3514.4]
  assign RetimeWrapper_clock = clock; // @[:@3503.4]
  assign RetimeWrapper_reset = reset; // @[:@3504.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3506.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3505.4]
endmodule
module StickySelects( // @[:@5017.2]
  input   clock, // @[:@5018.4]
  input   reset, // @[:@5019.4]
  input   io_ins_0, // @[:@5020.4]
  input   io_ins_1, // @[:@5020.4]
  input   io_ins_2, // @[:@5020.4]
  input   io_ins_3, // @[:@5020.4]
  input   io_ins_4, // @[:@5020.4]
  input   io_ins_5, // @[:@5020.4]
  output  io_outs_0, // @[:@5020.4]
  output  io_outs_1, // @[:@5020.4]
  output  io_outs_2, // @[:@5020.4]
  output  io_outs_3, // @[:@5020.4]
  output  io_outs_4, // @[:@5020.4]
  output  io_outs_5 // @[:@5020.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@5022.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@5023.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@5024.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@5025.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@5026.4]
  wire  _T_25; // @[StickySelects.scala 24:52:@5027.4]
  wire  _T_26; // @[StickySelects.scala 24:21:@5028.4]
  reg  _T_29; // @[StickySelects.scala 21:22:@5030.4]
  reg [31:0] _RAND_1;
  wire  _T_30; // @[StickySelects.scala 22:54:@5031.4]
  wire  _T_31; // @[StickySelects.scala 22:54:@5032.4]
  wire  _T_32; // @[StickySelects.scala 22:54:@5033.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@5034.4]
  wire  _T_35; // @[StickySelects.scala 24:52:@5035.4]
  wire  _T_36; // @[StickySelects.scala 24:21:@5036.4]
  reg  _T_39; // @[StickySelects.scala 21:22:@5038.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[StickySelects.scala 22:54:@5039.4]
  wire  _T_41; // @[StickySelects.scala 22:54:@5040.4]
  wire  _T_42; // @[StickySelects.scala 22:54:@5041.4]
  wire  _T_43; // @[StickySelects.scala 22:54:@5042.4]
  wire  _T_45; // @[StickySelects.scala 24:52:@5043.4]
  wire  _T_46; // @[StickySelects.scala 24:21:@5044.4]
  reg  _T_49; // @[StickySelects.scala 21:22:@5046.4]
  reg [31:0] _RAND_3;
  wire  _T_51; // @[StickySelects.scala 22:54:@5048.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@5049.4]
  wire  _T_53; // @[StickySelects.scala 22:54:@5050.4]
  wire  _T_55; // @[StickySelects.scala 24:52:@5051.4]
  wire  _T_56; // @[StickySelects.scala 24:21:@5052.4]
  reg  _T_59; // @[StickySelects.scala 21:22:@5054.4]
  reg [31:0] _RAND_4;
  wire  _T_62; // @[StickySelects.scala 22:54:@5057.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@5058.4]
  wire  _T_65; // @[StickySelects.scala 24:52:@5059.4]
  wire  _T_66; // @[StickySelects.scala 24:21:@5060.4]
  reg  _T_69; // @[StickySelects.scala 21:22:@5062.4]
  reg [31:0] _RAND_5;
  wire  _T_73; // @[StickySelects.scala 22:54:@5066.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@5067.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@5068.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@5023.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@5024.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@5025.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@5026.4]
  assign _T_25 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@5027.4]
  assign _T_26 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 24:21:@5028.4]
  assign _T_30 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@5031.4]
  assign _T_31 = _T_30 | io_ins_3; // @[StickySelects.scala 22:54:@5032.4]
  assign _T_32 = _T_31 | io_ins_4; // @[StickySelects.scala 22:54:@5033.4]
  assign _T_33 = _T_32 | io_ins_5; // @[StickySelects.scala 22:54:@5034.4]
  assign _T_35 = io_ins_1 | _T_29; // @[StickySelects.scala 24:52:@5035.4]
  assign _T_36 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 24:21:@5036.4]
  assign _T_40 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@5039.4]
  assign _T_41 = _T_40 | io_ins_3; // @[StickySelects.scala 22:54:@5040.4]
  assign _T_42 = _T_41 | io_ins_4; // @[StickySelects.scala 22:54:@5041.4]
  assign _T_43 = _T_42 | io_ins_5; // @[StickySelects.scala 22:54:@5042.4]
  assign _T_45 = io_ins_2 | _T_39; // @[StickySelects.scala 24:52:@5043.4]
  assign _T_46 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 24:21:@5044.4]
  assign _T_51 = _T_40 | io_ins_2; // @[StickySelects.scala 22:54:@5048.4]
  assign _T_52 = _T_51 | io_ins_4; // @[StickySelects.scala 22:54:@5049.4]
  assign _T_53 = _T_52 | io_ins_5; // @[StickySelects.scala 22:54:@5050.4]
  assign _T_55 = io_ins_3 | _T_49; // @[StickySelects.scala 24:52:@5051.4]
  assign _T_56 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 24:21:@5052.4]
  assign _T_62 = _T_51 | io_ins_3; // @[StickySelects.scala 22:54:@5057.4]
  assign _T_63 = _T_62 | io_ins_5; // @[StickySelects.scala 22:54:@5058.4]
  assign _T_65 = io_ins_4 | _T_59; // @[StickySelects.scala 24:52:@5059.4]
  assign _T_66 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 24:21:@5060.4]
  assign _T_73 = _T_62 | io_ins_4; // @[StickySelects.scala 22:54:@5066.4]
  assign _T_75 = io_ins_5 | _T_69; // @[StickySelects.scala 24:52:@5067.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@5068.4]
  assign io_outs_0 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 28:52:@5070.4]
  assign io_outs_1 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 28:52:@5071.4]
  assign io_outs_2 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 28:52:@5072.4]
  assign io_outs_3 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 28:52:@5073.4]
  assign io_outs_4 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 28:52:@5074.4]
  assign io_outs_5 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@5075.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_49 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_59 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_69 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_23) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_25;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_33) begin
        _T_29 <= 1'h0;
      end else begin
        _T_29 <= _T_35;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_43) begin
        _T_39 <= 1'h0;
      end else begin
        _T_39 <= _T_45;
      end
    end
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_53) begin
        _T_49 <= 1'h0;
      end else begin
        _T_49 <= _T_55;
      end
    end
    if (reset) begin
      _T_59 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_59 <= 1'h0;
      end else begin
        _T_59 <= _T_65;
      end
    end
    if (reset) begin
      _T_69 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_69 <= 1'h0;
      end else begin
        _T_69 <= _T_75;
      end
    end
  end
endmodule
module RetimeWrapper_36( // @[:@5989.2]
  input   clock, // @[:@5990.4]
  input   reset, // @[:@5991.4]
  input   io_flow, // @[:@5992.4]
  input   io_in, // @[:@5992.4]
  output  io_out // @[:@5992.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5994.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5994.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5994.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5994.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5994.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5994.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5994.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6007.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6006.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6005.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6004.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6003.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6001.4]
endmodule
module x257_lb_0( // @[:@9049.2]
  input        clock, // @[:@9050.4]
  input        reset, // @[:@9051.4]
  input  [2:0] io_rPort_11_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_11_ofs_0, // @[:@9052.4]
  input        io_rPort_11_en_0, // @[:@9052.4]
  input        io_rPort_11_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_11_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_10_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_10_ofs_0, // @[:@9052.4]
  input        io_rPort_10_en_0, // @[:@9052.4]
  input        io_rPort_10_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_10_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_9_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_9_ofs_0, // @[:@9052.4]
  input        io_rPort_9_en_0, // @[:@9052.4]
  input        io_rPort_9_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_9_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_8_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_8_ofs_0, // @[:@9052.4]
  input        io_rPort_8_en_0, // @[:@9052.4]
  input        io_rPort_8_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_8_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_7_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_7_ofs_0, // @[:@9052.4]
  input        io_rPort_7_en_0, // @[:@9052.4]
  input        io_rPort_7_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_7_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_6_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_6_ofs_0, // @[:@9052.4]
  input        io_rPort_6_en_0, // @[:@9052.4]
  input        io_rPort_6_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_6_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_5_ofs_0, // @[:@9052.4]
  input        io_rPort_5_en_0, // @[:@9052.4]
  input        io_rPort_5_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_5_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_4_ofs_0, // @[:@9052.4]
  input        io_rPort_4_en_0, // @[:@9052.4]
  input        io_rPort_4_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_4_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_3_ofs_0, // @[:@9052.4]
  input        io_rPort_3_en_0, // @[:@9052.4]
  input        io_rPort_3_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_3_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_2_ofs_0, // @[:@9052.4]
  input        io_rPort_2_en_0, // @[:@9052.4]
  input        io_rPort_2_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_2_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_1_ofs_0, // @[:@9052.4]
  input        io_rPort_1_en_0, // @[:@9052.4]
  input        io_rPort_1_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_1_output_0, // @[:@9052.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@9052.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@9052.4]
  input  [8:0] io_rPort_0_ofs_0, // @[:@9052.4]
  input        io_rPort_0_en_0, // @[:@9052.4]
  input        io_rPort_0_backpressure, // @[:@9052.4]
  output [7:0] io_rPort_0_output_0, // @[:@9052.4]
  input  [2:0] io_wPort_1_banks_1, // @[:@9052.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@9052.4]
  input  [8:0] io_wPort_1_ofs_0, // @[:@9052.4]
  input  [7:0] io_wPort_1_data_0, // @[:@9052.4]
  input        io_wPort_1_en_0, // @[:@9052.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@9052.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@9052.4]
  input  [8:0] io_wPort_0_ofs_0, // @[:@9052.4]
  input  [7:0] io_wPort_0_data_0, // @[:@9052.4]
  input        io_wPort_0_en_0 // @[:@9052.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@9143.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@9143.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9143.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9143.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9143.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@9143.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@9143.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@9143.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@9159.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@9159.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9159.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9159.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9159.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@9159.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@9159.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@9159.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@9175.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@9175.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9175.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9175.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9175.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@9175.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@9175.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@9175.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@9191.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@9191.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9191.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9191.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9191.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@9191.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@9191.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@9191.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@9207.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@9207.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9207.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9207.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9207.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@9207.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@9207.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@9207.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@9223.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@9223.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9223.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9223.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9223.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@9223.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@9223.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@9223.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@9239.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@9239.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9239.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9239.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9239.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@9239.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@9239.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@9239.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@9255.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@9255.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9255.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9255.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9255.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@9255.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@9255.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@9255.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@9271.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@9271.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9271.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9271.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9271.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@9271.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@9271.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@9271.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@9287.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@9287.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9287.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9287.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9287.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@9287.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@9287.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@9287.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@9303.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@9303.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9303.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9303.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9303.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@9303.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@9303.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@9303.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@9319.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@9319.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9319.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9319.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9319.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@9319.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@9319.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@9319.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@9335.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@9335.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9335.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9335.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9335.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@9335.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@9335.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@9335.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@9351.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@9351.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9351.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9351.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9351.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@9351.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@9351.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@9351.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@9367.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@9367.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9367.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9367.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9367.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@9367.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@9367.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@9367.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@9383.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@9383.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9383.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9383.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9383.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@9383.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@9383.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@9383.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@9615.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@9677.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@9739.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@9801.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@9863.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@9925.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@9987.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@10049.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@10111.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@10173.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@10235.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@10297.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@10359.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@10421.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@10483.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@10545.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10608.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10608.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10608.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10608.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10608.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10616.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10616.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10616.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10616.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10616.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10624.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10624.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10624.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10624.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10624.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10632.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10632.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10632.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10632.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10632.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10640.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10640.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10640.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10640.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10640.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10648.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10648.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10648.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10648.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10648.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10656.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10656.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10656.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10656.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10656.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@10664.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@10664.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@10664.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@10664.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@10664.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@10704.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@10704.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@10704.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@10704.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@10704.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@10712.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@10712.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@10712.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@10712.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@10712.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@10720.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@10720.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@10720.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@10720.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@10720.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@10728.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@10728.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@10728.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@10728.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@10728.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@10736.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@10736.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@10736.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@10736.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@10736.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@10744.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@10744.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@10744.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@10744.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@10744.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@10752.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@10752.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@10752.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@10752.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@10752.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@10760.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@10760.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@10760.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@10760.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@10760.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@10800.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@10800.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@10800.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@10800.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@10800.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@10808.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@10808.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@10808.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@10808.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@10808.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@10816.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@10816.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@10816.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@10816.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@10816.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@10824.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@10824.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@10824.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@10824.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@10824.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@10832.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@10832.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@10832.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@10832.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@10832.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@10840.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@10840.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@10840.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@10840.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@10840.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@10848.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@10848.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@10848.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@10848.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@10848.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@10856.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@10856.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@10856.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@10856.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@10856.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@10896.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@10896.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@10896.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@10896.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@10896.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@10904.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@10904.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@10904.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@10904.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@10904.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@10912.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@10912.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@10912.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@10912.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@10912.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@10920.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@10920.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@10920.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@10920.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@10920.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@10928.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@10928.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@10928.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@10928.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@10928.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@10936.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@10936.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@10936.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@10936.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@10936.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@10944.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@10944.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@10944.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@10944.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@10944.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@10952.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@10952.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@10952.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@10952.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@10952.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@10992.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@10992.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@10992.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@10992.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@10992.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@11000.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@11000.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@11000.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@11000.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@11000.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@11008.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@11008.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@11008.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@11008.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@11008.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@11016.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@11016.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@11016.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@11016.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@11016.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@11024.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@11024.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@11024.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@11024.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@11024.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@11032.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@11032.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@11032.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@11032.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@11032.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@11040.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@11040.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@11040.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@11040.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@11040.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@11048.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@11048.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@11048.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@11048.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@11048.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@11088.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@11088.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@11088.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@11088.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@11088.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@11096.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@11096.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@11096.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@11096.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@11096.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@11104.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@11104.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@11104.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@11104.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@11104.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@11112.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@11112.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@11112.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@11112.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@11112.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@11120.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@11120.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@11120.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@11120.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@11120.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@11128.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@11128.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@11128.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@11128.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@11128.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@11136.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@11136.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@11136.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@11136.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@11136.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@11144.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@11144.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@11144.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@11144.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@11144.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@11184.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@11184.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@11184.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@11184.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@11184.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@11200.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@11200.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@11200.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@11200.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@11200.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@11208.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@11208.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@11208.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@11208.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@11208.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@11216.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@11216.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@11216.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@11216.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@11216.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@11224.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@11224.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@11224.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@11224.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@11224.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@11232.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@11232.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@11232.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@11232.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@11232.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@11240.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@11240.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@11240.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@11240.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@11240.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@11280.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@11280.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@11280.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@11280.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@11280.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@11288.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@11288.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@11288.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@11288.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@11288.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@11296.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@11296.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@11296.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@11296.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@11296.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@11312.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@11312.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@11312.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@11312.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@11312.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@11320.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@11320.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@11320.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@11320.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@11320.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@11328.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@11328.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@11328.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@11328.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@11328.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@11336.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@11336.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@11336.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@11336.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@11336.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@11376.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@11376.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@11376.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@11376.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@11376.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@11384.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@11384.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@11384.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@11384.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@11384.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@11392.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@11392.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@11392.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@11392.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@11392.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@11400.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@11400.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@11400.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@11400.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@11400.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@11408.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@11408.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@11408.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@11408.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@11408.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@11416.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@11416.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@11416.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@11416.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@11416.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@11424.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@11424.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@11424.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@11424.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@11424.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@11432.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@11432.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@11432.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@11432.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@11432.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@11472.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@11472.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@11472.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@11472.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@11472.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@11480.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@11480.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@11480.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@11480.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@11480.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@11488.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@11488.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@11488.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@11488.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@11488.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@11496.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@11496.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@11496.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@11496.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@11496.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@11504.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@11504.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@11504.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@11504.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@11504.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@11512.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@11512.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@11512.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@11512.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@11512.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@11520.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@11520.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@11520.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@11520.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@11520.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@11528.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@11528.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@11528.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@11528.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@11528.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@11568.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@11568.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@11568.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@11568.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@11568.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@11576.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@11576.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@11576.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@11576.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@11576.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@11584.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@11584.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@11584.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@11584.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@11584.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@11592.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@11592.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@11592.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@11592.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@11592.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@11600.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@11600.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@11600.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@11600.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@11600.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@11608.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@11608.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@11608.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@11608.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@11608.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@11616.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@11616.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@11616.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@11616.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@11616.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@11624.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@11624.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@11624.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@11624.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@11624.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@11664.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@11664.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@11664.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@11664.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@11664.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@11672.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@11672.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@11672.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@11672.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@11672.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@11680.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@11680.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@11680.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@11680.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@11680.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@11688.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@11688.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@11688.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@11688.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@11688.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@11696.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@11696.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@11696.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@11696.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@11696.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@11704.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@11704.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@11704.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@11704.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@11704.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@11712.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@11712.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@11712.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@11712.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@11712.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@11720.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@11720.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@11720.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@11720.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@11720.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@9399.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@9400.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@9401.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@9402.4]
  wire [17:0] _T_450; // @[Cat.scala 30:58:@9404.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@9411.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@9412.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@9413.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@9414.4]
  wire [17:0] _T_461; // @[Cat.scala 30:58:@9416.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@9424.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@9425.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@9426.4]
  wire [17:0] _T_472; // @[Cat.scala 30:58:@9428.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@9436.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@9437.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@9438.4]
  wire [17:0] _T_483; // @[Cat.scala 30:58:@9440.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@9447.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@9449.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@9450.4]
  wire [17:0] _T_494; // @[Cat.scala 30:58:@9452.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@9459.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@9461.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@9462.4]
  wire [17:0] _T_505; // @[Cat.scala 30:58:@9464.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@9473.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@9474.4]
  wire [17:0] _T_516; // @[Cat.scala 30:58:@9476.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@9485.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@9486.4]
  wire [17:0] _T_527; // @[Cat.scala 30:58:@9488.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@9495.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@9497.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@9498.4]
  wire [17:0] _T_538; // @[Cat.scala 30:58:@9500.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@9507.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@9509.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@9510.4]
  wire [17:0] _T_549; // @[Cat.scala 30:58:@9512.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@9521.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@9522.4]
  wire [17:0] _T_560; // @[Cat.scala 30:58:@9524.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@9533.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@9534.4]
  wire [17:0] _T_571; // @[Cat.scala 30:58:@9536.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@9543.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@9545.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@9546.4]
  wire [17:0] _T_582; // @[Cat.scala 30:58:@9548.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@9555.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@9557.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@9558.4]
  wire [17:0] _T_593; // @[Cat.scala 30:58:@9560.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@9569.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@9570.4]
  wire [17:0] _T_604; // @[Cat.scala 30:58:@9572.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@9581.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@9582.4]
  wire [17:0] _T_615; // @[Cat.scala 30:58:@9584.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@9591.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@9592.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@9593.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@9595.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@9596.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@9597.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@9599.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@9600.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@9601.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@9603.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@9604.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@9605.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@9607.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@9608.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@9609.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@9611.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@9612.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@9613.4]
  wire  _T_655; // @[MemPrimitives.scala 123:41:@9624.4]
  wire  _T_656; // @[MemPrimitives.scala 123:41:@9625.4]
  wire  _T_657; // @[MemPrimitives.scala 123:41:@9626.4]
  wire  _T_658; // @[MemPrimitives.scala 123:41:@9627.4]
  wire  _T_659; // @[MemPrimitives.scala 123:41:@9628.4]
  wire  _T_660; // @[MemPrimitives.scala 123:41:@9629.4]
  wire [10:0] _T_662; // @[Cat.scala 30:58:@9631.4]
  wire [10:0] _T_664; // @[Cat.scala 30:58:@9633.4]
  wire [10:0] _T_666; // @[Cat.scala 30:58:@9635.4]
  wire [10:0] _T_668; // @[Cat.scala 30:58:@9637.4]
  wire [10:0] _T_670; // @[Cat.scala 30:58:@9639.4]
  wire [10:0] _T_672; // @[Cat.scala 30:58:@9641.4]
  wire [10:0] _T_673; // @[Mux.scala 31:69:@9642.4]
  wire [10:0] _T_674; // @[Mux.scala 31:69:@9643.4]
  wire [10:0] _T_675; // @[Mux.scala 31:69:@9644.4]
  wire [10:0] _T_676; // @[Mux.scala 31:69:@9645.4]
  wire [10:0] _T_677; // @[Mux.scala 31:69:@9646.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@9653.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@9654.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@9655.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@9657.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@9658.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@9659.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@9661.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@9662.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@9663.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@9665.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@9666.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@9667.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@9669.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@9670.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@9671.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@9673.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@9674.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@9675.4]
  wire  _T_717; // @[MemPrimitives.scala 123:41:@9686.4]
  wire  _T_718; // @[MemPrimitives.scala 123:41:@9687.4]
  wire  _T_719; // @[MemPrimitives.scala 123:41:@9688.4]
  wire  _T_720; // @[MemPrimitives.scala 123:41:@9689.4]
  wire  _T_721; // @[MemPrimitives.scala 123:41:@9690.4]
  wire  _T_722; // @[MemPrimitives.scala 123:41:@9691.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@9693.4]
  wire [10:0] _T_726; // @[Cat.scala 30:58:@9695.4]
  wire [10:0] _T_728; // @[Cat.scala 30:58:@9697.4]
  wire [10:0] _T_730; // @[Cat.scala 30:58:@9699.4]
  wire [10:0] _T_732; // @[Cat.scala 30:58:@9701.4]
  wire [10:0] _T_734; // @[Cat.scala 30:58:@9703.4]
  wire [10:0] _T_735; // @[Mux.scala 31:69:@9704.4]
  wire [10:0] _T_736; // @[Mux.scala 31:69:@9705.4]
  wire [10:0] _T_737; // @[Mux.scala 31:69:@9706.4]
  wire [10:0] _T_738; // @[Mux.scala 31:69:@9707.4]
  wire [10:0] _T_739; // @[Mux.scala 31:69:@9708.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@9716.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@9717.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@9720.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@9721.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@9724.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@9725.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@9728.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@9729.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@9732.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@9733.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@9736.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@9737.4]
  wire  _T_779; // @[MemPrimitives.scala 123:41:@9748.4]
  wire  _T_780; // @[MemPrimitives.scala 123:41:@9749.4]
  wire  _T_781; // @[MemPrimitives.scala 123:41:@9750.4]
  wire  _T_782; // @[MemPrimitives.scala 123:41:@9751.4]
  wire  _T_783; // @[MemPrimitives.scala 123:41:@9752.4]
  wire  _T_784; // @[MemPrimitives.scala 123:41:@9753.4]
  wire [10:0] _T_786; // @[Cat.scala 30:58:@9755.4]
  wire [10:0] _T_788; // @[Cat.scala 30:58:@9757.4]
  wire [10:0] _T_790; // @[Cat.scala 30:58:@9759.4]
  wire [10:0] _T_792; // @[Cat.scala 30:58:@9761.4]
  wire [10:0] _T_794; // @[Cat.scala 30:58:@9763.4]
  wire [10:0] _T_796; // @[Cat.scala 30:58:@9765.4]
  wire [10:0] _T_797; // @[Mux.scala 31:69:@9766.4]
  wire [10:0] _T_798; // @[Mux.scala 31:69:@9767.4]
  wire [10:0] _T_799; // @[Mux.scala 31:69:@9768.4]
  wire [10:0] _T_800; // @[Mux.scala 31:69:@9769.4]
  wire [10:0] _T_801; // @[Mux.scala 31:69:@9770.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@9778.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@9779.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@9782.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@9783.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@9786.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@9787.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@9790.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@9791.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@9794.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@9795.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@9798.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@9799.4]
  wire  _T_841; // @[MemPrimitives.scala 123:41:@9810.4]
  wire  _T_842; // @[MemPrimitives.scala 123:41:@9811.4]
  wire  _T_843; // @[MemPrimitives.scala 123:41:@9812.4]
  wire  _T_844; // @[MemPrimitives.scala 123:41:@9813.4]
  wire  _T_845; // @[MemPrimitives.scala 123:41:@9814.4]
  wire  _T_846; // @[MemPrimitives.scala 123:41:@9815.4]
  wire [10:0] _T_848; // @[Cat.scala 30:58:@9817.4]
  wire [10:0] _T_850; // @[Cat.scala 30:58:@9819.4]
  wire [10:0] _T_852; // @[Cat.scala 30:58:@9821.4]
  wire [10:0] _T_854; // @[Cat.scala 30:58:@9823.4]
  wire [10:0] _T_856; // @[Cat.scala 30:58:@9825.4]
  wire [10:0] _T_858; // @[Cat.scala 30:58:@9827.4]
  wire [10:0] _T_859; // @[Mux.scala 31:69:@9828.4]
  wire [10:0] _T_860; // @[Mux.scala 31:69:@9829.4]
  wire [10:0] _T_861; // @[Mux.scala 31:69:@9830.4]
  wire [10:0] _T_862; // @[Mux.scala 31:69:@9831.4]
  wire [10:0] _T_863; // @[Mux.scala 31:69:@9832.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@9839.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@9841.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@9843.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@9845.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@9847.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@9849.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@9851.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@9853.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@9855.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@9857.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@9859.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@9861.4]
  wire  _T_903; // @[MemPrimitives.scala 123:41:@9872.4]
  wire  _T_904; // @[MemPrimitives.scala 123:41:@9873.4]
  wire  _T_905; // @[MemPrimitives.scala 123:41:@9874.4]
  wire  _T_906; // @[MemPrimitives.scala 123:41:@9875.4]
  wire  _T_907; // @[MemPrimitives.scala 123:41:@9876.4]
  wire  _T_908; // @[MemPrimitives.scala 123:41:@9877.4]
  wire [10:0] _T_910; // @[Cat.scala 30:58:@9879.4]
  wire [10:0] _T_912; // @[Cat.scala 30:58:@9881.4]
  wire [10:0] _T_914; // @[Cat.scala 30:58:@9883.4]
  wire [10:0] _T_916; // @[Cat.scala 30:58:@9885.4]
  wire [10:0] _T_918; // @[Cat.scala 30:58:@9887.4]
  wire [10:0] _T_920; // @[Cat.scala 30:58:@9889.4]
  wire [10:0] _T_921; // @[Mux.scala 31:69:@9890.4]
  wire [10:0] _T_922; // @[Mux.scala 31:69:@9891.4]
  wire [10:0] _T_923; // @[Mux.scala 31:69:@9892.4]
  wire [10:0] _T_924; // @[Mux.scala 31:69:@9893.4]
  wire [10:0] _T_925; // @[Mux.scala 31:69:@9894.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@9901.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@9903.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@9905.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@9907.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@9909.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@9911.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@9913.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@9915.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@9917.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@9919.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@9921.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@9923.4]
  wire  _T_965; // @[MemPrimitives.scala 123:41:@9934.4]
  wire  _T_966; // @[MemPrimitives.scala 123:41:@9935.4]
  wire  _T_967; // @[MemPrimitives.scala 123:41:@9936.4]
  wire  _T_968; // @[MemPrimitives.scala 123:41:@9937.4]
  wire  _T_969; // @[MemPrimitives.scala 123:41:@9938.4]
  wire  _T_970; // @[MemPrimitives.scala 123:41:@9939.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@9941.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@9943.4]
  wire [10:0] _T_976; // @[Cat.scala 30:58:@9945.4]
  wire [10:0] _T_978; // @[Cat.scala 30:58:@9947.4]
  wire [10:0] _T_980; // @[Cat.scala 30:58:@9949.4]
  wire [10:0] _T_982; // @[Cat.scala 30:58:@9951.4]
  wire [10:0] _T_983; // @[Mux.scala 31:69:@9952.4]
  wire [10:0] _T_984; // @[Mux.scala 31:69:@9953.4]
  wire [10:0] _T_985; // @[Mux.scala 31:69:@9954.4]
  wire [10:0] _T_986; // @[Mux.scala 31:69:@9955.4]
  wire [10:0] _T_987; // @[Mux.scala 31:69:@9956.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@9965.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@9969.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@9973.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@9977.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@9981.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@9985.4]
  wire  _T_1027; // @[MemPrimitives.scala 123:41:@9996.4]
  wire  _T_1028; // @[MemPrimitives.scala 123:41:@9997.4]
  wire  _T_1029; // @[MemPrimitives.scala 123:41:@9998.4]
  wire  _T_1030; // @[MemPrimitives.scala 123:41:@9999.4]
  wire  _T_1031; // @[MemPrimitives.scala 123:41:@10000.4]
  wire  _T_1032; // @[MemPrimitives.scala 123:41:@10001.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@10003.4]
  wire [10:0] _T_1036; // @[Cat.scala 30:58:@10005.4]
  wire [10:0] _T_1038; // @[Cat.scala 30:58:@10007.4]
  wire [10:0] _T_1040; // @[Cat.scala 30:58:@10009.4]
  wire [10:0] _T_1042; // @[Cat.scala 30:58:@10011.4]
  wire [10:0] _T_1044; // @[Cat.scala 30:58:@10013.4]
  wire [10:0] _T_1045; // @[Mux.scala 31:69:@10014.4]
  wire [10:0] _T_1046; // @[Mux.scala 31:69:@10015.4]
  wire [10:0] _T_1047; // @[Mux.scala 31:69:@10016.4]
  wire [10:0] _T_1048; // @[Mux.scala 31:69:@10017.4]
  wire [10:0] _T_1049; // @[Mux.scala 31:69:@10018.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@10027.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@10031.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@10035.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@10039.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@10043.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@10047.4]
  wire  _T_1089; // @[MemPrimitives.scala 123:41:@10058.4]
  wire  _T_1090; // @[MemPrimitives.scala 123:41:@10059.4]
  wire  _T_1091; // @[MemPrimitives.scala 123:41:@10060.4]
  wire  _T_1092; // @[MemPrimitives.scala 123:41:@10061.4]
  wire  _T_1093; // @[MemPrimitives.scala 123:41:@10062.4]
  wire  _T_1094; // @[MemPrimitives.scala 123:41:@10063.4]
  wire [10:0] _T_1096; // @[Cat.scala 30:58:@10065.4]
  wire [10:0] _T_1098; // @[Cat.scala 30:58:@10067.4]
  wire [10:0] _T_1100; // @[Cat.scala 30:58:@10069.4]
  wire [10:0] _T_1102; // @[Cat.scala 30:58:@10071.4]
  wire [10:0] _T_1104; // @[Cat.scala 30:58:@10073.4]
  wire [10:0] _T_1106; // @[Cat.scala 30:58:@10075.4]
  wire [10:0] _T_1107; // @[Mux.scala 31:69:@10076.4]
  wire [10:0] _T_1108; // @[Mux.scala 31:69:@10077.4]
  wire [10:0] _T_1109; // @[Mux.scala 31:69:@10078.4]
  wire [10:0] _T_1110; // @[Mux.scala 31:69:@10079.4]
  wire [10:0] _T_1111; // @[Mux.scala 31:69:@10080.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@10087.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@10089.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@10091.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@10093.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@10095.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@10097.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@10099.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@10101.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@10103.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@10105.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@10107.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@10109.4]
  wire  _T_1151; // @[MemPrimitives.scala 123:41:@10120.4]
  wire  _T_1152; // @[MemPrimitives.scala 123:41:@10121.4]
  wire  _T_1153; // @[MemPrimitives.scala 123:41:@10122.4]
  wire  _T_1154; // @[MemPrimitives.scala 123:41:@10123.4]
  wire  _T_1155; // @[MemPrimitives.scala 123:41:@10124.4]
  wire  _T_1156; // @[MemPrimitives.scala 123:41:@10125.4]
  wire [10:0] _T_1158; // @[Cat.scala 30:58:@10127.4]
  wire [10:0] _T_1160; // @[Cat.scala 30:58:@10129.4]
  wire [10:0] _T_1162; // @[Cat.scala 30:58:@10131.4]
  wire [10:0] _T_1164; // @[Cat.scala 30:58:@10133.4]
  wire [10:0] _T_1166; // @[Cat.scala 30:58:@10135.4]
  wire [10:0] _T_1168; // @[Cat.scala 30:58:@10137.4]
  wire [10:0] _T_1169; // @[Mux.scala 31:69:@10138.4]
  wire [10:0] _T_1170; // @[Mux.scala 31:69:@10139.4]
  wire [10:0] _T_1171; // @[Mux.scala 31:69:@10140.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@10141.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@10142.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@10149.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@10151.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@10153.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@10155.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@10157.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@10159.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@10161.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@10163.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@10165.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@10167.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@10169.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@10171.4]
  wire  _T_1213; // @[MemPrimitives.scala 123:41:@10182.4]
  wire  _T_1214; // @[MemPrimitives.scala 123:41:@10183.4]
  wire  _T_1215; // @[MemPrimitives.scala 123:41:@10184.4]
  wire  _T_1216; // @[MemPrimitives.scala 123:41:@10185.4]
  wire  _T_1217; // @[MemPrimitives.scala 123:41:@10186.4]
  wire  _T_1218; // @[MemPrimitives.scala 123:41:@10187.4]
  wire [10:0] _T_1220; // @[Cat.scala 30:58:@10189.4]
  wire [10:0] _T_1222; // @[Cat.scala 30:58:@10191.4]
  wire [10:0] _T_1224; // @[Cat.scala 30:58:@10193.4]
  wire [10:0] _T_1226; // @[Cat.scala 30:58:@10195.4]
  wire [10:0] _T_1228; // @[Cat.scala 30:58:@10197.4]
  wire [10:0] _T_1230; // @[Cat.scala 30:58:@10199.4]
  wire [10:0] _T_1231; // @[Mux.scala 31:69:@10200.4]
  wire [10:0] _T_1232; // @[Mux.scala 31:69:@10201.4]
  wire [10:0] _T_1233; // @[Mux.scala 31:69:@10202.4]
  wire [10:0] _T_1234; // @[Mux.scala 31:69:@10203.4]
  wire [10:0] _T_1235; // @[Mux.scala 31:69:@10204.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@10213.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@10217.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@10221.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@10225.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@10229.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@10233.4]
  wire  _T_1275; // @[MemPrimitives.scala 123:41:@10244.4]
  wire  _T_1276; // @[MemPrimitives.scala 123:41:@10245.4]
  wire  _T_1277; // @[MemPrimitives.scala 123:41:@10246.4]
  wire  _T_1278; // @[MemPrimitives.scala 123:41:@10247.4]
  wire  _T_1279; // @[MemPrimitives.scala 123:41:@10248.4]
  wire  _T_1280; // @[MemPrimitives.scala 123:41:@10249.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@10251.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@10253.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@10255.4]
  wire [10:0] _T_1288; // @[Cat.scala 30:58:@10257.4]
  wire [10:0] _T_1290; // @[Cat.scala 30:58:@10259.4]
  wire [10:0] _T_1292; // @[Cat.scala 30:58:@10261.4]
  wire [10:0] _T_1293; // @[Mux.scala 31:69:@10262.4]
  wire [10:0] _T_1294; // @[Mux.scala 31:69:@10263.4]
  wire [10:0] _T_1295; // @[Mux.scala 31:69:@10264.4]
  wire [10:0] _T_1296; // @[Mux.scala 31:69:@10265.4]
  wire [10:0] _T_1297; // @[Mux.scala 31:69:@10266.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@10275.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@10279.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@10283.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@10287.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@10291.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@10295.4]
  wire  _T_1337; // @[MemPrimitives.scala 123:41:@10306.4]
  wire  _T_1338; // @[MemPrimitives.scala 123:41:@10307.4]
  wire  _T_1339; // @[MemPrimitives.scala 123:41:@10308.4]
  wire  _T_1340; // @[MemPrimitives.scala 123:41:@10309.4]
  wire  _T_1341; // @[MemPrimitives.scala 123:41:@10310.4]
  wire  _T_1342; // @[MemPrimitives.scala 123:41:@10311.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@10313.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@10315.4]
  wire [10:0] _T_1348; // @[Cat.scala 30:58:@10317.4]
  wire [10:0] _T_1350; // @[Cat.scala 30:58:@10319.4]
  wire [10:0] _T_1352; // @[Cat.scala 30:58:@10321.4]
  wire [10:0] _T_1354; // @[Cat.scala 30:58:@10323.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@10324.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@10325.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@10326.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@10327.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@10328.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@10335.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@10337.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@10339.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@10341.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@10343.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@10345.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@10347.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@10349.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@10351.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@10353.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@10355.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@10357.4]
  wire  _T_1399; // @[MemPrimitives.scala 123:41:@10368.4]
  wire  _T_1400; // @[MemPrimitives.scala 123:41:@10369.4]
  wire  _T_1401; // @[MemPrimitives.scala 123:41:@10370.4]
  wire  _T_1402; // @[MemPrimitives.scala 123:41:@10371.4]
  wire  _T_1403; // @[MemPrimitives.scala 123:41:@10372.4]
  wire  _T_1404; // @[MemPrimitives.scala 123:41:@10373.4]
  wire [10:0] _T_1406; // @[Cat.scala 30:58:@10375.4]
  wire [10:0] _T_1408; // @[Cat.scala 30:58:@10377.4]
  wire [10:0] _T_1410; // @[Cat.scala 30:58:@10379.4]
  wire [10:0] _T_1412; // @[Cat.scala 30:58:@10381.4]
  wire [10:0] _T_1414; // @[Cat.scala 30:58:@10383.4]
  wire [10:0] _T_1416; // @[Cat.scala 30:58:@10385.4]
  wire [10:0] _T_1417; // @[Mux.scala 31:69:@10386.4]
  wire [10:0] _T_1418; // @[Mux.scala 31:69:@10387.4]
  wire [10:0] _T_1419; // @[Mux.scala 31:69:@10388.4]
  wire [10:0] _T_1420; // @[Mux.scala 31:69:@10389.4]
  wire [10:0] _T_1421; // @[Mux.scala 31:69:@10390.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@10397.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@10399.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@10401.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@10403.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@10405.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@10407.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@10409.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@10411.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@10413.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@10415.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@10417.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@10419.4]
  wire  _T_1461; // @[MemPrimitives.scala 123:41:@10430.4]
  wire  _T_1462; // @[MemPrimitives.scala 123:41:@10431.4]
  wire  _T_1463; // @[MemPrimitives.scala 123:41:@10432.4]
  wire  _T_1464; // @[MemPrimitives.scala 123:41:@10433.4]
  wire  _T_1465; // @[MemPrimitives.scala 123:41:@10434.4]
  wire  _T_1466; // @[MemPrimitives.scala 123:41:@10435.4]
  wire [10:0] _T_1468; // @[Cat.scala 30:58:@10437.4]
  wire [10:0] _T_1470; // @[Cat.scala 30:58:@10439.4]
  wire [10:0] _T_1472; // @[Cat.scala 30:58:@10441.4]
  wire [10:0] _T_1474; // @[Cat.scala 30:58:@10443.4]
  wire [10:0] _T_1476; // @[Cat.scala 30:58:@10445.4]
  wire [10:0] _T_1478; // @[Cat.scala 30:58:@10447.4]
  wire [10:0] _T_1479; // @[Mux.scala 31:69:@10448.4]
  wire [10:0] _T_1480; // @[Mux.scala 31:69:@10449.4]
  wire [10:0] _T_1481; // @[Mux.scala 31:69:@10450.4]
  wire [10:0] _T_1482; // @[Mux.scala 31:69:@10451.4]
  wire [10:0] _T_1483; // @[Mux.scala 31:69:@10452.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@10461.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@10465.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@10469.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@10473.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@10477.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@10481.4]
  wire  _T_1523; // @[MemPrimitives.scala 123:41:@10492.4]
  wire  _T_1524; // @[MemPrimitives.scala 123:41:@10493.4]
  wire  _T_1525; // @[MemPrimitives.scala 123:41:@10494.4]
  wire  _T_1526; // @[MemPrimitives.scala 123:41:@10495.4]
  wire  _T_1527; // @[MemPrimitives.scala 123:41:@10496.4]
  wire  _T_1528; // @[MemPrimitives.scala 123:41:@10497.4]
  wire [10:0] _T_1530; // @[Cat.scala 30:58:@10499.4]
  wire [10:0] _T_1532; // @[Cat.scala 30:58:@10501.4]
  wire [10:0] _T_1534; // @[Cat.scala 30:58:@10503.4]
  wire [10:0] _T_1536; // @[Cat.scala 30:58:@10505.4]
  wire [10:0] _T_1538; // @[Cat.scala 30:58:@10507.4]
  wire [10:0] _T_1540; // @[Cat.scala 30:58:@10509.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@10510.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@10511.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@10512.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@10513.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@10514.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@10523.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@10527.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@10531.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@10535.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@10539.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@10543.4]
  wire  _T_1585; // @[MemPrimitives.scala 123:41:@10554.4]
  wire  _T_1586; // @[MemPrimitives.scala 123:41:@10555.4]
  wire  _T_1587; // @[MemPrimitives.scala 123:41:@10556.4]
  wire  _T_1588; // @[MemPrimitives.scala 123:41:@10557.4]
  wire  _T_1589; // @[MemPrimitives.scala 123:41:@10558.4]
  wire  _T_1590; // @[MemPrimitives.scala 123:41:@10559.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@10561.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@10563.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@10565.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@10567.4]
  wire [10:0] _T_1600; // @[Cat.scala 30:58:@10569.4]
  wire [10:0] _T_1602; // @[Cat.scala 30:58:@10571.4]
  wire [10:0] _T_1603; // @[Mux.scala 31:69:@10572.4]
  wire [10:0] _T_1604; // @[Mux.scala 31:69:@10573.4]
  wire [10:0] _T_1605; // @[Mux.scala 31:69:@10574.4]
  wire [10:0] _T_1606; // @[Mux.scala 31:69:@10575.4]
  wire [10:0] _T_1607; // @[Mux.scala 31:69:@10576.4]
  wire  _T_1671; // @[package.scala 96:25:@10661.4 package.scala 96:25:@10662.4]
  wire [7:0] _T_1675; // @[Mux.scala 31:69:@10671.4]
  wire  _T_1668; // @[package.scala 96:25:@10653.4 package.scala 96:25:@10654.4]
  wire [7:0] _T_1676; // @[Mux.scala 31:69:@10672.4]
  wire  _T_1665; // @[package.scala 96:25:@10645.4 package.scala 96:25:@10646.4]
  wire [7:0] _T_1677; // @[Mux.scala 31:69:@10673.4]
  wire  _T_1662; // @[package.scala 96:25:@10637.4 package.scala 96:25:@10638.4]
  wire [7:0] _T_1678; // @[Mux.scala 31:69:@10674.4]
  wire  _T_1659; // @[package.scala 96:25:@10629.4 package.scala 96:25:@10630.4]
  wire [7:0] _T_1679; // @[Mux.scala 31:69:@10675.4]
  wire  _T_1656; // @[package.scala 96:25:@10621.4 package.scala 96:25:@10622.4]
  wire [7:0] _T_1680; // @[Mux.scala 31:69:@10676.4]
  wire  _T_1653; // @[package.scala 96:25:@10613.4 package.scala 96:25:@10614.4]
  wire  _T_1742; // @[package.scala 96:25:@10757.4 package.scala 96:25:@10758.4]
  wire [7:0] _T_1746; // @[Mux.scala 31:69:@10767.4]
  wire  _T_1739; // @[package.scala 96:25:@10749.4 package.scala 96:25:@10750.4]
  wire [7:0] _T_1747; // @[Mux.scala 31:69:@10768.4]
  wire  _T_1736; // @[package.scala 96:25:@10741.4 package.scala 96:25:@10742.4]
  wire [7:0] _T_1748; // @[Mux.scala 31:69:@10769.4]
  wire  _T_1733; // @[package.scala 96:25:@10733.4 package.scala 96:25:@10734.4]
  wire [7:0] _T_1749; // @[Mux.scala 31:69:@10770.4]
  wire  _T_1730; // @[package.scala 96:25:@10725.4 package.scala 96:25:@10726.4]
  wire [7:0] _T_1750; // @[Mux.scala 31:69:@10771.4]
  wire  _T_1727; // @[package.scala 96:25:@10717.4 package.scala 96:25:@10718.4]
  wire [7:0] _T_1751; // @[Mux.scala 31:69:@10772.4]
  wire  _T_1724; // @[package.scala 96:25:@10709.4 package.scala 96:25:@10710.4]
  wire  _T_1813; // @[package.scala 96:25:@10853.4 package.scala 96:25:@10854.4]
  wire [7:0] _T_1817; // @[Mux.scala 31:69:@10863.4]
  wire  _T_1810; // @[package.scala 96:25:@10845.4 package.scala 96:25:@10846.4]
  wire [7:0] _T_1818; // @[Mux.scala 31:69:@10864.4]
  wire  _T_1807; // @[package.scala 96:25:@10837.4 package.scala 96:25:@10838.4]
  wire [7:0] _T_1819; // @[Mux.scala 31:69:@10865.4]
  wire  _T_1804; // @[package.scala 96:25:@10829.4 package.scala 96:25:@10830.4]
  wire [7:0] _T_1820; // @[Mux.scala 31:69:@10866.4]
  wire  _T_1801; // @[package.scala 96:25:@10821.4 package.scala 96:25:@10822.4]
  wire [7:0] _T_1821; // @[Mux.scala 31:69:@10867.4]
  wire  _T_1798; // @[package.scala 96:25:@10813.4 package.scala 96:25:@10814.4]
  wire [7:0] _T_1822; // @[Mux.scala 31:69:@10868.4]
  wire  _T_1795; // @[package.scala 96:25:@10805.4 package.scala 96:25:@10806.4]
  wire  _T_1884; // @[package.scala 96:25:@10949.4 package.scala 96:25:@10950.4]
  wire [7:0] _T_1888; // @[Mux.scala 31:69:@10959.4]
  wire  _T_1881; // @[package.scala 96:25:@10941.4 package.scala 96:25:@10942.4]
  wire [7:0] _T_1889; // @[Mux.scala 31:69:@10960.4]
  wire  _T_1878; // @[package.scala 96:25:@10933.4 package.scala 96:25:@10934.4]
  wire [7:0] _T_1890; // @[Mux.scala 31:69:@10961.4]
  wire  _T_1875; // @[package.scala 96:25:@10925.4 package.scala 96:25:@10926.4]
  wire [7:0] _T_1891; // @[Mux.scala 31:69:@10962.4]
  wire  _T_1872; // @[package.scala 96:25:@10917.4 package.scala 96:25:@10918.4]
  wire [7:0] _T_1892; // @[Mux.scala 31:69:@10963.4]
  wire  _T_1869; // @[package.scala 96:25:@10909.4 package.scala 96:25:@10910.4]
  wire [7:0] _T_1893; // @[Mux.scala 31:69:@10964.4]
  wire  _T_1866; // @[package.scala 96:25:@10901.4 package.scala 96:25:@10902.4]
  wire  _T_1955; // @[package.scala 96:25:@11045.4 package.scala 96:25:@11046.4]
  wire [7:0] _T_1959; // @[Mux.scala 31:69:@11055.4]
  wire  _T_1952; // @[package.scala 96:25:@11037.4 package.scala 96:25:@11038.4]
  wire [7:0] _T_1960; // @[Mux.scala 31:69:@11056.4]
  wire  _T_1949; // @[package.scala 96:25:@11029.4 package.scala 96:25:@11030.4]
  wire [7:0] _T_1961; // @[Mux.scala 31:69:@11057.4]
  wire  _T_1946; // @[package.scala 96:25:@11021.4 package.scala 96:25:@11022.4]
  wire [7:0] _T_1962; // @[Mux.scala 31:69:@11058.4]
  wire  _T_1943; // @[package.scala 96:25:@11013.4 package.scala 96:25:@11014.4]
  wire [7:0] _T_1963; // @[Mux.scala 31:69:@11059.4]
  wire  _T_1940; // @[package.scala 96:25:@11005.4 package.scala 96:25:@11006.4]
  wire [7:0] _T_1964; // @[Mux.scala 31:69:@11060.4]
  wire  _T_1937; // @[package.scala 96:25:@10997.4 package.scala 96:25:@10998.4]
  wire  _T_2026; // @[package.scala 96:25:@11141.4 package.scala 96:25:@11142.4]
  wire [7:0] _T_2030; // @[Mux.scala 31:69:@11151.4]
  wire  _T_2023; // @[package.scala 96:25:@11133.4 package.scala 96:25:@11134.4]
  wire [7:0] _T_2031; // @[Mux.scala 31:69:@11152.4]
  wire  _T_2020; // @[package.scala 96:25:@11125.4 package.scala 96:25:@11126.4]
  wire [7:0] _T_2032; // @[Mux.scala 31:69:@11153.4]
  wire  _T_2017; // @[package.scala 96:25:@11117.4 package.scala 96:25:@11118.4]
  wire [7:0] _T_2033; // @[Mux.scala 31:69:@11154.4]
  wire  _T_2014; // @[package.scala 96:25:@11109.4 package.scala 96:25:@11110.4]
  wire [7:0] _T_2034; // @[Mux.scala 31:69:@11155.4]
  wire  _T_2011; // @[package.scala 96:25:@11101.4 package.scala 96:25:@11102.4]
  wire [7:0] _T_2035; // @[Mux.scala 31:69:@11156.4]
  wire  _T_2008; // @[package.scala 96:25:@11093.4 package.scala 96:25:@11094.4]
  wire  _T_2097; // @[package.scala 96:25:@11237.4 package.scala 96:25:@11238.4]
  wire [7:0] _T_2101; // @[Mux.scala 31:69:@11247.4]
  wire  _T_2094; // @[package.scala 96:25:@11229.4 package.scala 96:25:@11230.4]
  wire [7:0] _T_2102; // @[Mux.scala 31:69:@11248.4]
  wire  _T_2091; // @[package.scala 96:25:@11221.4 package.scala 96:25:@11222.4]
  wire [7:0] _T_2103; // @[Mux.scala 31:69:@11249.4]
  wire  _T_2088; // @[package.scala 96:25:@11213.4 package.scala 96:25:@11214.4]
  wire [7:0] _T_2104; // @[Mux.scala 31:69:@11250.4]
  wire  _T_2085; // @[package.scala 96:25:@11205.4 package.scala 96:25:@11206.4]
  wire [7:0] _T_2105; // @[Mux.scala 31:69:@11251.4]
  wire  _T_2082; // @[package.scala 96:25:@11197.4 package.scala 96:25:@11198.4]
  wire [7:0] _T_2106; // @[Mux.scala 31:69:@11252.4]
  wire  _T_2079; // @[package.scala 96:25:@11189.4 package.scala 96:25:@11190.4]
  wire  _T_2168; // @[package.scala 96:25:@11333.4 package.scala 96:25:@11334.4]
  wire [7:0] _T_2172; // @[Mux.scala 31:69:@11343.4]
  wire  _T_2165; // @[package.scala 96:25:@11325.4 package.scala 96:25:@11326.4]
  wire [7:0] _T_2173; // @[Mux.scala 31:69:@11344.4]
  wire  _T_2162; // @[package.scala 96:25:@11317.4 package.scala 96:25:@11318.4]
  wire [7:0] _T_2174; // @[Mux.scala 31:69:@11345.4]
  wire  _T_2159; // @[package.scala 96:25:@11309.4 package.scala 96:25:@11310.4]
  wire [7:0] _T_2175; // @[Mux.scala 31:69:@11346.4]
  wire  _T_2156; // @[package.scala 96:25:@11301.4 package.scala 96:25:@11302.4]
  wire [7:0] _T_2176; // @[Mux.scala 31:69:@11347.4]
  wire  _T_2153; // @[package.scala 96:25:@11293.4 package.scala 96:25:@11294.4]
  wire [7:0] _T_2177; // @[Mux.scala 31:69:@11348.4]
  wire  _T_2150; // @[package.scala 96:25:@11285.4 package.scala 96:25:@11286.4]
  wire  _T_2239; // @[package.scala 96:25:@11429.4 package.scala 96:25:@11430.4]
  wire [7:0] _T_2243; // @[Mux.scala 31:69:@11439.4]
  wire  _T_2236; // @[package.scala 96:25:@11421.4 package.scala 96:25:@11422.4]
  wire [7:0] _T_2244; // @[Mux.scala 31:69:@11440.4]
  wire  _T_2233; // @[package.scala 96:25:@11413.4 package.scala 96:25:@11414.4]
  wire [7:0] _T_2245; // @[Mux.scala 31:69:@11441.4]
  wire  _T_2230; // @[package.scala 96:25:@11405.4 package.scala 96:25:@11406.4]
  wire [7:0] _T_2246; // @[Mux.scala 31:69:@11442.4]
  wire  _T_2227; // @[package.scala 96:25:@11397.4 package.scala 96:25:@11398.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@11443.4]
  wire  _T_2224; // @[package.scala 96:25:@11389.4 package.scala 96:25:@11390.4]
  wire [7:0] _T_2248; // @[Mux.scala 31:69:@11444.4]
  wire  _T_2221; // @[package.scala 96:25:@11381.4 package.scala 96:25:@11382.4]
  wire  _T_2310; // @[package.scala 96:25:@11525.4 package.scala 96:25:@11526.4]
  wire [7:0] _T_2314; // @[Mux.scala 31:69:@11535.4]
  wire  _T_2307; // @[package.scala 96:25:@11517.4 package.scala 96:25:@11518.4]
  wire [7:0] _T_2315; // @[Mux.scala 31:69:@11536.4]
  wire  _T_2304; // @[package.scala 96:25:@11509.4 package.scala 96:25:@11510.4]
  wire [7:0] _T_2316; // @[Mux.scala 31:69:@11537.4]
  wire  _T_2301; // @[package.scala 96:25:@11501.4 package.scala 96:25:@11502.4]
  wire [7:0] _T_2317; // @[Mux.scala 31:69:@11538.4]
  wire  _T_2298; // @[package.scala 96:25:@11493.4 package.scala 96:25:@11494.4]
  wire [7:0] _T_2318; // @[Mux.scala 31:69:@11539.4]
  wire  _T_2295; // @[package.scala 96:25:@11485.4 package.scala 96:25:@11486.4]
  wire [7:0] _T_2319; // @[Mux.scala 31:69:@11540.4]
  wire  _T_2292; // @[package.scala 96:25:@11477.4 package.scala 96:25:@11478.4]
  wire  _T_2381; // @[package.scala 96:25:@11621.4 package.scala 96:25:@11622.4]
  wire [7:0] _T_2385; // @[Mux.scala 31:69:@11631.4]
  wire  _T_2378; // @[package.scala 96:25:@11613.4 package.scala 96:25:@11614.4]
  wire [7:0] _T_2386; // @[Mux.scala 31:69:@11632.4]
  wire  _T_2375; // @[package.scala 96:25:@11605.4 package.scala 96:25:@11606.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@11633.4]
  wire  _T_2372; // @[package.scala 96:25:@11597.4 package.scala 96:25:@11598.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@11634.4]
  wire  _T_2369; // @[package.scala 96:25:@11589.4 package.scala 96:25:@11590.4]
  wire [7:0] _T_2389; // @[Mux.scala 31:69:@11635.4]
  wire  _T_2366; // @[package.scala 96:25:@11581.4 package.scala 96:25:@11582.4]
  wire [7:0] _T_2390; // @[Mux.scala 31:69:@11636.4]
  wire  _T_2363; // @[package.scala 96:25:@11573.4 package.scala 96:25:@11574.4]
  wire  _T_2452; // @[package.scala 96:25:@11717.4 package.scala 96:25:@11718.4]
  wire [7:0] _T_2456; // @[Mux.scala 31:69:@11727.4]
  wire  _T_2449; // @[package.scala 96:25:@11709.4 package.scala 96:25:@11710.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@11728.4]
  wire  _T_2446; // @[package.scala 96:25:@11701.4 package.scala 96:25:@11702.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@11729.4]
  wire  _T_2443; // @[package.scala 96:25:@11693.4 package.scala 96:25:@11694.4]
  wire [7:0] _T_2459; // @[Mux.scala 31:69:@11730.4]
  wire  _T_2440; // @[package.scala 96:25:@11685.4 package.scala 96:25:@11686.4]
  wire [7:0] _T_2460; // @[Mux.scala 31:69:@11731.4]
  wire  _T_2437; // @[package.scala 96:25:@11677.4 package.scala 96:25:@11678.4]
  wire [7:0] _T_2461; // @[Mux.scala 31:69:@11732.4]
  wire  _T_2434; // @[package.scala 96:25:@11669.4 package.scala 96:25:@11670.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@9143.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@9159.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@9175.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@9191.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@9207.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@9223.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@9239.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@9255.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@9271.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@9287.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@9303.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@9319.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@9335.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@9351.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@9367.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@9383.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@9615.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@9677.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@9739.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@9801.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@9863.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@9925.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@9987.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@10049.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@10111.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@10173.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects StickySelects_10 ( // @[MemPrimitives.scala 121:29:@10235.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects StickySelects_11 ( // @[MemPrimitives.scala 121:29:@10297.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@10359.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@10421.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects StickySelects_14 ( // @[MemPrimitives.scala 121:29:@10483.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects StickySelects_15 ( // @[MemPrimitives.scala 121:29:@10545.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_36 RetimeWrapper ( // @[package.scala 93:22:@10608.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_1 ( // @[package.scala 93:22:@10616.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_2 ( // @[package.scala 93:22:@10624.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_3 ( // @[package.scala 93:22:@10632.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_4 ( // @[package.scala 93:22:@10640.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_5 ( // @[package.scala 93:22:@10648.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_6 ( // @[package.scala 93:22:@10656.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_7 ( // @[package.scala 93:22:@10664.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_8 ( // @[package.scala 93:22:@10704.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_9 ( // @[package.scala 93:22:@10712.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_10 ( // @[package.scala 93:22:@10720.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_11 ( // @[package.scala 93:22:@10728.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_12 ( // @[package.scala 93:22:@10736.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_13 ( // @[package.scala 93:22:@10744.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_14 ( // @[package.scala 93:22:@10752.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_15 ( // @[package.scala 93:22:@10760.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_16 ( // @[package.scala 93:22:@10800.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_17 ( // @[package.scala 93:22:@10808.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_18 ( // @[package.scala 93:22:@10816.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_19 ( // @[package.scala 93:22:@10824.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_20 ( // @[package.scala 93:22:@10832.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_21 ( // @[package.scala 93:22:@10840.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_22 ( // @[package.scala 93:22:@10848.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_23 ( // @[package.scala 93:22:@10856.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_24 ( // @[package.scala 93:22:@10896.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_25 ( // @[package.scala 93:22:@10904.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_26 ( // @[package.scala 93:22:@10912.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_27 ( // @[package.scala 93:22:@10920.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_28 ( // @[package.scala 93:22:@10928.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_29 ( // @[package.scala 93:22:@10936.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_30 ( // @[package.scala 93:22:@10944.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_31 ( // @[package.scala 93:22:@10952.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_32 ( // @[package.scala 93:22:@10992.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_33 ( // @[package.scala 93:22:@11000.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_34 ( // @[package.scala 93:22:@11008.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_35 ( // @[package.scala 93:22:@11016.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_36 ( // @[package.scala 93:22:@11024.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_37 ( // @[package.scala 93:22:@11032.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_38 ( // @[package.scala 93:22:@11040.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_39 ( // @[package.scala 93:22:@11048.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_40 ( // @[package.scala 93:22:@11088.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_41 ( // @[package.scala 93:22:@11096.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_42 ( // @[package.scala 93:22:@11104.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_43 ( // @[package.scala 93:22:@11112.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_44 ( // @[package.scala 93:22:@11120.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_45 ( // @[package.scala 93:22:@11128.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_46 ( // @[package.scala 93:22:@11136.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_47 ( // @[package.scala 93:22:@11144.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_48 ( // @[package.scala 93:22:@11184.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_49 ( // @[package.scala 93:22:@11192.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_50 ( // @[package.scala 93:22:@11200.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_51 ( // @[package.scala 93:22:@11208.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_52 ( // @[package.scala 93:22:@11216.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_53 ( // @[package.scala 93:22:@11224.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_54 ( // @[package.scala 93:22:@11232.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_55 ( // @[package.scala 93:22:@11240.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_56 ( // @[package.scala 93:22:@11280.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_57 ( // @[package.scala 93:22:@11288.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_58 ( // @[package.scala 93:22:@11296.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_59 ( // @[package.scala 93:22:@11304.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_60 ( // @[package.scala 93:22:@11312.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_61 ( // @[package.scala 93:22:@11320.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_62 ( // @[package.scala 93:22:@11328.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_63 ( // @[package.scala 93:22:@11336.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_64 ( // @[package.scala 93:22:@11376.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_65 ( // @[package.scala 93:22:@11384.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_66 ( // @[package.scala 93:22:@11392.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_67 ( // @[package.scala 93:22:@11400.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_68 ( // @[package.scala 93:22:@11408.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_69 ( // @[package.scala 93:22:@11416.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_70 ( // @[package.scala 93:22:@11424.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_71 ( // @[package.scala 93:22:@11432.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_72 ( // @[package.scala 93:22:@11472.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_73 ( // @[package.scala 93:22:@11480.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_74 ( // @[package.scala 93:22:@11488.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_75 ( // @[package.scala 93:22:@11496.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_76 ( // @[package.scala 93:22:@11504.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_77 ( // @[package.scala 93:22:@11512.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_78 ( // @[package.scala 93:22:@11520.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_79 ( // @[package.scala 93:22:@11528.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_80 ( // @[package.scala 93:22:@11568.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_81 ( // @[package.scala 93:22:@11576.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_82 ( // @[package.scala 93:22:@11584.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_83 ( // @[package.scala 93:22:@11592.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_84 ( // @[package.scala 93:22:@11600.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_85 ( // @[package.scala 93:22:@11608.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_86 ( // @[package.scala 93:22:@11616.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_87 ( // @[package.scala 93:22:@11624.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_88 ( // @[package.scala 93:22:@11664.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_89 ( // @[package.scala 93:22:@11672.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_90 ( // @[package.scala 93:22:@11680.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_91 ( // @[package.scala 93:22:@11688.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_92 ( // @[package.scala 93:22:@11696.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_93 ( // @[package.scala 93:22:@11704.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_94 ( // @[package.scala 93:22:@11712.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_95 ( // @[package.scala 93:22:@11720.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9399.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@9400.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@9401.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@9402.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9404.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9411.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@9412.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@9413.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@9414.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9416.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@9424.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@9425.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@9426.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9428.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@9436.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@9437.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@9438.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9440.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9447.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@9449.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@9450.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9452.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9459.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@9461.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@9462.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9464.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@9473.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@9474.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9476.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@9485.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@9486.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9488.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9495.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@9497.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@9498.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9500.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9507.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@9509.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@9510.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9512.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@9521.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@9522.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9524.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@9533.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@9534.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9536.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9543.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@9545.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@9546.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9548.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9555.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@9557.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@9558.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9560.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@9569.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@9570.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9572.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@9581.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@9582.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9584.4]
  assign _T_620 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9591.4]
  assign _T_622 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9592.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@9593.4]
  assign _T_626 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9595.4]
  assign _T_628 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9596.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@9597.4]
  assign _T_632 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9599.4]
  assign _T_634 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9600.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@9601.4]
  assign _T_638 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9603.4]
  assign _T_640 = io_rPort_5_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9604.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@9605.4]
  assign _T_644 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9607.4]
  assign _T_646 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9608.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@9609.4]
  assign _T_650 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9611.4]
  assign _T_652 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9612.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@9613.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@9624.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@9625.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@9626.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@9627.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@9628.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@9629.4]
  assign _T_662 = {_T_655,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9631.4]
  assign _T_664 = {_T_656,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9633.4]
  assign _T_666 = {_T_657,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9635.4]
  assign _T_668 = {_T_658,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9637.4]
  assign _T_670 = {_T_659,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9639.4]
  assign _T_672 = {_T_660,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9641.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@9642.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@9643.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@9644.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@9645.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@9646.4]
  assign _T_682 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9653.4]
  assign _T_684 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9654.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@9655.4]
  assign _T_688 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9657.4]
  assign _T_690 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9658.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@9659.4]
  assign _T_694 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9661.4]
  assign _T_696 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9662.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@9663.4]
  assign _T_700 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9665.4]
  assign _T_702 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9666.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@9667.4]
  assign _T_706 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9669.4]
  assign _T_708 = io_rPort_10_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9670.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@9671.4]
  assign _T_712 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9673.4]
  assign _T_714 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9674.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@9675.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@9686.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@9687.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@9688.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@9689.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@9690.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@9691.4]
  assign _T_724 = {_T_717,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9693.4]
  assign _T_726 = {_T_718,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9695.4]
  assign _T_728 = {_T_719,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9697.4]
  assign _T_730 = {_T_720,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9699.4]
  assign _T_732 = {_T_721,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9701.4]
  assign _T_734 = {_T_722,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9703.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@9704.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@9705.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@9706.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@9707.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@9708.4]
  assign _T_746 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9716.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@9717.4]
  assign _T_752 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9720.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@9721.4]
  assign _T_758 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9724.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@9725.4]
  assign _T_764 = io_rPort_5_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9728.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@9729.4]
  assign _T_770 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9732.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@9733.4]
  assign _T_776 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9736.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@9737.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@9748.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@9749.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@9750.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@9751.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@9752.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@9753.4]
  assign _T_786 = {_T_779,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9755.4]
  assign _T_788 = {_T_780,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9757.4]
  assign _T_790 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9759.4]
  assign _T_792 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9761.4]
  assign _T_794 = {_T_783,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9763.4]
  assign _T_796 = {_T_784,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9765.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@9766.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@9767.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@9768.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@9769.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@9770.4]
  assign _T_808 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9778.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@9779.4]
  assign _T_814 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9782.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@9783.4]
  assign _T_820 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9786.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@9787.4]
  assign _T_826 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9790.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@9791.4]
  assign _T_832 = io_rPort_10_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9794.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@9795.4]
  assign _T_838 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9798.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@9799.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@9810.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@9811.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@9812.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@9813.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@9814.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@9815.4]
  assign _T_848 = {_T_841,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9817.4]
  assign _T_850 = {_T_842,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9819.4]
  assign _T_852 = {_T_843,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9821.4]
  assign _T_854 = {_T_844,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9823.4]
  assign _T_856 = {_T_845,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9825.4]
  assign _T_858 = {_T_846,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9827.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@9828.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@9829.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@9830.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@9831.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@9832.4]
  assign _T_868 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9839.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@9841.4]
  assign _T_874 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9843.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@9845.4]
  assign _T_880 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9847.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@9849.4]
  assign _T_886 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9851.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@9853.4]
  assign _T_892 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9855.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@9857.4]
  assign _T_898 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9859.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@9861.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@9872.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@9873.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@9874.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@9875.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@9876.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@9877.4]
  assign _T_910 = {_T_903,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9879.4]
  assign _T_912 = {_T_904,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9881.4]
  assign _T_914 = {_T_905,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9883.4]
  assign _T_916 = {_T_906,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9885.4]
  assign _T_918 = {_T_907,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9887.4]
  assign _T_920 = {_T_908,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9889.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@9890.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@9891.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@9892.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@9893.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@9894.4]
  assign _T_930 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9901.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@9903.4]
  assign _T_936 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9905.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@9907.4]
  assign _T_942 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9909.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@9911.4]
  assign _T_948 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9913.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@9915.4]
  assign _T_954 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9917.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@9919.4]
  assign _T_960 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9921.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@9923.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@9934.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@9935.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@9936.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@9937.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@9938.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@9939.4]
  assign _T_972 = {_T_965,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9941.4]
  assign _T_974 = {_T_966,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9943.4]
  assign _T_976 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9945.4]
  assign _T_978 = {_T_968,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9947.4]
  assign _T_980 = {_T_969,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9949.4]
  assign _T_982 = {_T_970,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9951.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@9952.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@9953.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@9954.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@9955.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@9956.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@9965.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@9969.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@9973.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@9977.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@9981.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@9985.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@9996.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@9997.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@9998.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@9999.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@10000.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@10001.4]
  assign _T_1034 = {_T_1027,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10003.4]
  assign _T_1036 = {_T_1028,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10005.4]
  assign _T_1038 = {_T_1029,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10007.4]
  assign _T_1040 = {_T_1030,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10009.4]
  assign _T_1042 = {_T_1031,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10011.4]
  assign _T_1044 = {_T_1032,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10013.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@10014.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@10015.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@10016.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@10017.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@10018.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@10027.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@10031.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@10035.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@10039.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@10043.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@10047.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@10058.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@10059.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@10060.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@10061.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@10062.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@10063.4]
  assign _T_1096 = {_T_1089,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10065.4]
  assign _T_1098 = {_T_1090,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10067.4]
  assign _T_1100 = {_T_1091,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10069.4]
  assign _T_1102 = {_T_1092,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10071.4]
  assign _T_1104 = {_T_1093,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10073.4]
  assign _T_1106 = {_T_1094,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10075.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@10076.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@10077.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@10078.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@10079.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@10080.4]
  assign _T_1116 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10087.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@10089.4]
  assign _T_1122 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10091.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@10093.4]
  assign _T_1128 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10095.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@10097.4]
  assign _T_1134 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10099.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@10101.4]
  assign _T_1140 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10103.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@10105.4]
  assign _T_1146 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10107.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@10109.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@10120.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@10121.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@10122.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@10123.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@10124.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@10125.4]
  assign _T_1158 = {_T_1151,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10127.4]
  assign _T_1160 = {_T_1152,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10129.4]
  assign _T_1162 = {_T_1153,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10131.4]
  assign _T_1164 = {_T_1154,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10133.4]
  assign _T_1166 = {_T_1155,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10135.4]
  assign _T_1168 = {_T_1156,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10137.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@10138.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@10139.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@10140.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@10141.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@10142.4]
  assign _T_1178 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10149.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@10151.4]
  assign _T_1184 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10153.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@10155.4]
  assign _T_1190 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10157.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@10159.4]
  assign _T_1196 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10161.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@10163.4]
  assign _T_1202 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10165.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@10167.4]
  assign _T_1208 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10169.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@10171.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@10182.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@10183.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@10184.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@10185.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@10186.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@10187.4]
  assign _T_1220 = {_T_1213,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10189.4]
  assign _T_1222 = {_T_1214,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10191.4]
  assign _T_1224 = {_T_1215,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10193.4]
  assign _T_1226 = {_T_1216,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10195.4]
  assign _T_1228 = {_T_1217,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10197.4]
  assign _T_1230 = {_T_1218,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10199.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@10200.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@10201.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@10202.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@10203.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@10204.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@10213.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@10217.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@10221.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@10225.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@10229.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@10233.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@10244.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@10245.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@10246.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@10247.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@10248.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@10249.4]
  assign _T_1282 = {_T_1275,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10251.4]
  assign _T_1284 = {_T_1276,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10253.4]
  assign _T_1286 = {_T_1277,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10255.4]
  assign _T_1288 = {_T_1278,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10257.4]
  assign _T_1290 = {_T_1279,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10259.4]
  assign _T_1292 = {_T_1280,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10261.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@10262.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@10263.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@10264.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@10265.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@10266.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@10275.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@10279.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@10283.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@10287.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@10291.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@10295.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@10306.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@10307.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@10308.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@10309.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@10310.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@10311.4]
  assign _T_1344 = {_T_1337,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10313.4]
  assign _T_1346 = {_T_1338,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10315.4]
  assign _T_1348 = {_T_1339,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10317.4]
  assign _T_1350 = {_T_1340,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10319.4]
  assign _T_1352 = {_T_1341,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10321.4]
  assign _T_1354 = {_T_1342,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10323.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@10324.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@10325.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@10326.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@10327.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@10328.4]
  assign _T_1364 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10335.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@10337.4]
  assign _T_1370 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10339.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@10341.4]
  assign _T_1376 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10343.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@10345.4]
  assign _T_1382 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10347.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@10349.4]
  assign _T_1388 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10351.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@10353.4]
  assign _T_1394 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10355.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@10357.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@10368.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@10369.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@10370.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@10371.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@10372.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@10373.4]
  assign _T_1406 = {_T_1399,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10375.4]
  assign _T_1408 = {_T_1400,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10377.4]
  assign _T_1410 = {_T_1401,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10379.4]
  assign _T_1412 = {_T_1402,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10381.4]
  assign _T_1414 = {_T_1403,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10383.4]
  assign _T_1416 = {_T_1404,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10385.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@10386.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@10387.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@10388.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@10389.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@10390.4]
  assign _T_1426 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10397.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@10399.4]
  assign _T_1432 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10401.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@10403.4]
  assign _T_1438 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10405.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@10407.4]
  assign _T_1444 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10409.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@10411.4]
  assign _T_1450 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10413.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@10415.4]
  assign _T_1456 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10417.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@10419.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@10430.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@10431.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@10432.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@10433.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@10434.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@10435.4]
  assign _T_1468 = {_T_1461,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10437.4]
  assign _T_1470 = {_T_1462,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10439.4]
  assign _T_1472 = {_T_1463,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10441.4]
  assign _T_1474 = {_T_1464,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10443.4]
  assign _T_1476 = {_T_1465,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10445.4]
  assign _T_1478 = {_T_1466,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10447.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@10448.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@10449.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@10450.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@10451.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@10452.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@10461.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@10465.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@10469.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@10473.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@10477.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@10481.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@10492.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@10493.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@10494.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@10495.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@10496.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@10497.4]
  assign _T_1530 = {_T_1523,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10499.4]
  assign _T_1532 = {_T_1524,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10501.4]
  assign _T_1534 = {_T_1525,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10503.4]
  assign _T_1536 = {_T_1526,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10505.4]
  assign _T_1538 = {_T_1527,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10507.4]
  assign _T_1540 = {_T_1528,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10509.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@10510.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@10511.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@10512.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@10513.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@10514.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@10523.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@10527.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@10531.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@10535.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@10539.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@10543.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@10554.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@10555.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@10556.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@10557.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@10558.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@10559.4]
  assign _T_1592 = {_T_1585,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10561.4]
  assign _T_1594 = {_T_1586,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10563.4]
  assign _T_1596 = {_T_1587,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10565.4]
  assign _T_1598 = {_T_1588,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10567.4]
  assign _T_1600 = {_T_1589,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10569.4]
  assign _T_1602 = {_T_1590,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10571.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@10572.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@10573.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@10574.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@10575.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@10576.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@10661.4 package.scala 96:25:@10662.4]
  assign _T_1675 = _T_1671 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10671.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10653.4 package.scala 96:25:@10654.4]
  assign _T_1676 = _T_1668 ? Mem1D_10_io_output : _T_1675; // @[Mux.scala 31:69:@10672.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10645.4 package.scala 96:25:@10646.4]
  assign _T_1677 = _T_1665 ? Mem1D_8_io_output : _T_1676; // @[Mux.scala 31:69:@10673.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@10637.4 package.scala 96:25:@10638.4]
  assign _T_1678 = _T_1662 ? Mem1D_6_io_output : _T_1677; // @[Mux.scala 31:69:@10674.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@10629.4 package.scala 96:25:@10630.4]
  assign _T_1679 = _T_1659 ? Mem1D_4_io_output : _T_1678; // @[Mux.scala 31:69:@10675.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@10621.4 package.scala 96:25:@10622.4]
  assign _T_1680 = _T_1656 ? Mem1D_2_io_output : _T_1679; // @[Mux.scala 31:69:@10676.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@10613.4 package.scala 96:25:@10614.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@10757.4 package.scala 96:25:@10758.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10767.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@10749.4 package.scala 96:25:@10750.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@10768.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@10741.4 package.scala 96:25:@10742.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@10769.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@10733.4 package.scala 96:25:@10734.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@10770.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@10725.4 package.scala 96:25:@10726.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@10771.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@10717.4 package.scala 96:25:@10718.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@10772.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@10709.4 package.scala 96:25:@10710.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@10853.4 package.scala 96:25:@10854.4]
  assign _T_1817 = _T_1813 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10863.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@10845.4 package.scala 96:25:@10846.4]
  assign _T_1818 = _T_1810 ? Mem1D_10_io_output : _T_1817; // @[Mux.scala 31:69:@10864.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@10837.4 package.scala 96:25:@10838.4]
  assign _T_1819 = _T_1807 ? Mem1D_8_io_output : _T_1818; // @[Mux.scala 31:69:@10865.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@10829.4 package.scala 96:25:@10830.4]
  assign _T_1820 = _T_1804 ? Mem1D_6_io_output : _T_1819; // @[Mux.scala 31:69:@10866.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@10821.4 package.scala 96:25:@10822.4]
  assign _T_1821 = _T_1801 ? Mem1D_4_io_output : _T_1820; // @[Mux.scala 31:69:@10867.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@10813.4 package.scala 96:25:@10814.4]
  assign _T_1822 = _T_1798 ? Mem1D_2_io_output : _T_1821; // @[Mux.scala 31:69:@10868.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@10805.4 package.scala 96:25:@10806.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@10949.4 package.scala 96:25:@10950.4]
  assign _T_1888 = _T_1884 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10959.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@10941.4 package.scala 96:25:@10942.4]
  assign _T_1889 = _T_1881 ? Mem1D_11_io_output : _T_1888; // @[Mux.scala 31:69:@10960.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@10933.4 package.scala 96:25:@10934.4]
  assign _T_1890 = _T_1878 ? Mem1D_9_io_output : _T_1889; // @[Mux.scala 31:69:@10961.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@10925.4 package.scala 96:25:@10926.4]
  assign _T_1891 = _T_1875 ? Mem1D_7_io_output : _T_1890; // @[Mux.scala 31:69:@10962.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@10917.4 package.scala 96:25:@10918.4]
  assign _T_1892 = _T_1872 ? Mem1D_5_io_output : _T_1891; // @[Mux.scala 31:69:@10963.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@10909.4 package.scala 96:25:@10910.4]
  assign _T_1893 = _T_1869 ? Mem1D_3_io_output : _T_1892; // @[Mux.scala 31:69:@10964.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@10901.4 package.scala 96:25:@10902.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@11045.4 package.scala 96:25:@11046.4]
  assign _T_1959 = _T_1955 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11055.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@11037.4 package.scala 96:25:@11038.4]
  assign _T_1960 = _T_1952 ? Mem1D_10_io_output : _T_1959; // @[Mux.scala 31:69:@11056.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@11029.4 package.scala 96:25:@11030.4]
  assign _T_1961 = _T_1949 ? Mem1D_8_io_output : _T_1960; // @[Mux.scala 31:69:@11057.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@11021.4 package.scala 96:25:@11022.4]
  assign _T_1962 = _T_1946 ? Mem1D_6_io_output : _T_1961; // @[Mux.scala 31:69:@11058.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@11013.4 package.scala 96:25:@11014.4]
  assign _T_1963 = _T_1943 ? Mem1D_4_io_output : _T_1962; // @[Mux.scala 31:69:@11059.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@11005.4 package.scala 96:25:@11006.4]
  assign _T_1964 = _T_1940 ? Mem1D_2_io_output : _T_1963; // @[Mux.scala 31:69:@11060.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@10997.4 package.scala 96:25:@10998.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@11141.4 package.scala 96:25:@11142.4]
  assign _T_2030 = _T_2026 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11151.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@11133.4 package.scala 96:25:@11134.4]
  assign _T_2031 = _T_2023 ? Mem1D_10_io_output : _T_2030; // @[Mux.scala 31:69:@11152.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@11125.4 package.scala 96:25:@11126.4]
  assign _T_2032 = _T_2020 ? Mem1D_8_io_output : _T_2031; // @[Mux.scala 31:69:@11153.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@11117.4 package.scala 96:25:@11118.4]
  assign _T_2033 = _T_2017 ? Mem1D_6_io_output : _T_2032; // @[Mux.scala 31:69:@11154.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@11109.4 package.scala 96:25:@11110.4]
  assign _T_2034 = _T_2014 ? Mem1D_4_io_output : _T_2033; // @[Mux.scala 31:69:@11155.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@11101.4 package.scala 96:25:@11102.4]
  assign _T_2035 = _T_2011 ? Mem1D_2_io_output : _T_2034; // @[Mux.scala 31:69:@11156.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@11093.4 package.scala 96:25:@11094.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@11237.4 package.scala 96:25:@11238.4]
  assign _T_2101 = _T_2097 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11247.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@11229.4 package.scala 96:25:@11230.4]
  assign _T_2102 = _T_2094 ? Mem1D_11_io_output : _T_2101; // @[Mux.scala 31:69:@11248.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@11221.4 package.scala 96:25:@11222.4]
  assign _T_2103 = _T_2091 ? Mem1D_9_io_output : _T_2102; // @[Mux.scala 31:69:@11249.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@11213.4 package.scala 96:25:@11214.4]
  assign _T_2104 = _T_2088 ? Mem1D_7_io_output : _T_2103; // @[Mux.scala 31:69:@11250.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@11205.4 package.scala 96:25:@11206.4]
  assign _T_2105 = _T_2085 ? Mem1D_5_io_output : _T_2104; // @[Mux.scala 31:69:@11251.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@11197.4 package.scala 96:25:@11198.4]
  assign _T_2106 = _T_2082 ? Mem1D_3_io_output : _T_2105; // @[Mux.scala 31:69:@11252.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@11189.4 package.scala 96:25:@11190.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@11333.4 package.scala 96:25:@11334.4]
  assign _T_2172 = _T_2168 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11343.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@11325.4 package.scala 96:25:@11326.4]
  assign _T_2173 = _T_2165 ? Mem1D_10_io_output : _T_2172; // @[Mux.scala 31:69:@11344.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@11317.4 package.scala 96:25:@11318.4]
  assign _T_2174 = _T_2162 ? Mem1D_8_io_output : _T_2173; // @[Mux.scala 31:69:@11345.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@11309.4 package.scala 96:25:@11310.4]
  assign _T_2175 = _T_2159 ? Mem1D_6_io_output : _T_2174; // @[Mux.scala 31:69:@11346.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@11301.4 package.scala 96:25:@11302.4]
  assign _T_2176 = _T_2156 ? Mem1D_4_io_output : _T_2175; // @[Mux.scala 31:69:@11347.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@11293.4 package.scala 96:25:@11294.4]
  assign _T_2177 = _T_2153 ? Mem1D_2_io_output : _T_2176; // @[Mux.scala 31:69:@11348.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@11285.4 package.scala 96:25:@11286.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@11429.4 package.scala 96:25:@11430.4]
  assign _T_2243 = _T_2239 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11439.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@11421.4 package.scala 96:25:@11422.4]
  assign _T_2244 = _T_2236 ? Mem1D_10_io_output : _T_2243; // @[Mux.scala 31:69:@11440.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@11413.4 package.scala 96:25:@11414.4]
  assign _T_2245 = _T_2233 ? Mem1D_8_io_output : _T_2244; // @[Mux.scala 31:69:@11441.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@11405.4 package.scala 96:25:@11406.4]
  assign _T_2246 = _T_2230 ? Mem1D_6_io_output : _T_2245; // @[Mux.scala 31:69:@11442.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@11397.4 package.scala 96:25:@11398.4]
  assign _T_2247 = _T_2227 ? Mem1D_4_io_output : _T_2246; // @[Mux.scala 31:69:@11443.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@11389.4 package.scala 96:25:@11390.4]
  assign _T_2248 = _T_2224 ? Mem1D_2_io_output : _T_2247; // @[Mux.scala 31:69:@11444.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@11381.4 package.scala 96:25:@11382.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@11525.4 package.scala 96:25:@11526.4]
  assign _T_2314 = _T_2310 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11535.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@11517.4 package.scala 96:25:@11518.4]
  assign _T_2315 = _T_2307 ? Mem1D_11_io_output : _T_2314; // @[Mux.scala 31:69:@11536.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@11509.4 package.scala 96:25:@11510.4]
  assign _T_2316 = _T_2304 ? Mem1D_9_io_output : _T_2315; // @[Mux.scala 31:69:@11537.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@11501.4 package.scala 96:25:@11502.4]
  assign _T_2317 = _T_2301 ? Mem1D_7_io_output : _T_2316; // @[Mux.scala 31:69:@11538.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@11493.4 package.scala 96:25:@11494.4]
  assign _T_2318 = _T_2298 ? Mem1D_5_io_output : _T_2317; // @[Mux.scala 31:69:@11539.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@11485.4 package.scala 96:25:@11486.4]
  assign _T_2319 = _T_2295 ? Mem1D_3_io_output : _T_2318; // @[Mux.scala 31:69:@11540.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@11477.4 package.scala 96:25:@11478.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@11621.4 package.scala 96:25:@11622.4]
  assign _T_2385 = _T_2381 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11631.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@11613.4 package.scala 96:25:@11614.4]
  assign _T_2386 = _T_2378 ? Mem1D_11_io_output : _T_2385; // @[Mux.scala 31:69:@11632.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@11605.4 package.scala 96:25:@11606.4]
  assign _T_2387 = _T_2375 ? Mem1D_9_io_output : _T_2386; // @[Mux.scala 31:69:@11633.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@11597.4 package.scala 96:25:@11598.4]
  assign _T_2388 = _T_2372 ? Mem1D_7_io_output : _T_2387; // @[Mux.scala 31:69:@11634.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@11589.4 package.scala 96:25:@11590.4]
  assign _T_2389 = _T_2369 ? Mem1D_5_io_output : _T_2388; // @[Mux.scala 31:69:@11635.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@11581.4 package.scala 96:25:@11582.4]
  assign _T_2390 = _T_2366 ? Mem1D_3_io_output : _T_2389; // @[Mux.scala 31:69:@11636.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@11573.4 package.scala 96:25:@11574.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@11717.4 package.scala 96:25:@11718.4]
  assign _T_2456 = _T_2452 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11727.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@11709.4 package.scala 96:25:@11710.4]
  assign _T_2457 = _T_2449 ? Mem1D_11_io_output : _T_2456; // @[Mux.scala 31:69:@11728.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@11701.4 package.scala 96:25:@11702.4]
  assign _T_2458 = _T_2446 ? Mem1D_9_io_output : _T_2457; // @[Mux.scala 31:69:@11729.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@11693.4 package.scala 96:25:@11694.4]
  assign _T_2459 = _T_2443 ? Mem1D_7_io_output : _T_2458; // @[Mux.scala 31:69:@11730.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@11685.4 package.scala 96:25:@11686.4]
  assign _T_2460 = _T_2440 ? Mem1D_5_io_output : _T_2459; // @[Mux.scala 31:69:@11731.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@11677.4 package.scala 96:25:@11678.4]
  assign _T_2461 = _T_2437 ? Mem1D_3_io_output : _T_2460; // @[Mux.scala 31:69:@11732.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@11669.4 package.scala 96:25:@11670.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_1_io_output : _T_2461; // @[MemPrimitives.scala 148:13:@11734.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_1_io_output : _T_2390; // @[MemPrimitives.scala 148:13:@11638.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_1_io_output : _T_2319; // @[MemPrimitives.scala 148:13:@11542.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_io_output : _T_2248; // @[MemPrimitives.scala 148:13:@11446.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_io_output : _T_2177; // @[MemPrimitives.scala 148:13:@11350.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_1_io_output : _T_2106; // @[MemPrimitives.scala 148:13:@11254.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_io_output : _T_2035; // @[MemPrimitives.scala 148:13:@11158.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_io_output : _T_1964; // @[MemPrimitives.scala 148:13:@11062.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_1_io_output : _T_1893; // @[MemPrimitives.scala 148:13:@10966.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_io_output : _T_1822; // @[MemPrimitives.scala 148:13:@10870.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 148:13:@10774.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_io_output : _T_1680; // @[MemPrimitives.scala 148:13:@10678.4]
  assign Mem1D_clock = clock; // @[:@9144.4]
  assign Mem1D_reset = reset; // @[:@9145.4]
  assign Mem1D_io_r_ofs_0 = _T_677[8:0]; // @[MemPrimitives.scala 127:28:@9650.4]
  assign Mem1D_io_r_backpressure = _T_677[9]; // @[MemPrimitives.scala 128:32:@9651.4]
  assign Mem1D_io_w_ofs_0 = _T_450[8:0]; // @[MemPrimitives.scala 94:28:@9408.4]
  assign Mem1D_io_w_data_0 = _T_450[16:9]; // @[MemPrimitives.scala 95:29:@9409.4]
  assign Mem1D_io_w_en_0 = _T_450[17]; // @[MemPrimitives.scala 96:27:@9410.4]
  assign Mem1D_1_clock = clock; // @[:@9160.4]
  assign Mem1D_1_reset = reset; // @[:@9161.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[8:0]; // @[MemPrimitives.scala 127:28:@9712.4]
  assign Mem1D_1_io_r_backpressure = _T_739[9]; // @[MemPrimitives.scala 128:32:@9713.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[8:0]; // @[MemPrimitives.scala 94:28:@9420.4]
  assign Mem1D_1_io_w_data_0 = _T_461[16:9]; // @[MemPrimitives.scala 95:29:@9421.4]
  assign Mem1D_1_io_w_en_0 = _T_461[17]; // @[MemPrimitives.scala 96:27:@9422.4]
  assign Mem1D_2_clock = clock; // @[:@9176.4]
  assign Mem1D_2_reset = reset; // @[:@9177.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[8:0]; // @[MemPrimitives.scala 127:28:@9774.4]
  assign Mem1D_2_io_r_backpressure = _T_801[9]; // @[MemPrimitives.scala 128:32:@9775.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[8:0]; // @[MemPrimitives.scala 94:28:@9432.4]
  assign Mem1D_2_io_w_data_0 = _T_472[16:9]; // @[MemPrimitives.scala 95:29:@9433.4]
  assign Mem1D_2_io_w_en_0 = _T_472[17]; // @[MemPrimitives.scala 96:27:@9434.4]
  assign Mem1D_3_clock = clock; // @[:@9192.4]
  assign Mem1D_3_reset = reset; // @[:@9193.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[8:0]; // @[MemPrimitives.scala 127:28:@9836.4]
  assign Mem1D_3_io_r_backpressure = _T_863[9]; // @[MemPrimitives.scala 128:32:@9837.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[8:0]; // @[MemPrimitives.scala 94:28:@9444.4]
  assign Mem1D_3_io_w_data_0 = _T_483[16:9]; // @[MemPrimitives.scala 95:29:@9445.4]
  assign Mem1D_3_io_w_en_0 = _T_483[17]; // @[MemPrimitives.scala 96:27:@9446.4]
  assign Mem1D_4_clock = clock; // @[:@9208.4]
  assign Mem1D_4_reset = reset; // @[:@9209.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[8:0]; // @[MemPrimitives.scala 127:28:@9898.4]
  assign Mem1D_4_io_r_backpressure = _T_925[9]; // @[MemPrimitives.scala 128:32:@9899.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[8:0]; // @[MemPrimitives.scala 94:28:@9456.4]
  assign Mem1D_4_io_w_data_0 = _T_494[16:9]; // @[MemPrimitives.scala 95:29:@9457.4]
  assign Mem1D_4_io_w_en_0 = _T_494[17]; // @[MemPrimitives.scala 96:27:@9458.4]
  assign Mem1D_5_clock = clock; // @[:@9224.4]
  assign Mem1D_5_reset = reset; // @[:@9225.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[8:0]; // @[MemPrimitives.scala 127:28:@9960.4]
  assign Mem1D_5_io_r_backpressure = _T_987[9]; // @[MemPrimitives.scala 128:32:@9961.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[8:0]; // @[MemPrimitives.scala 94:28:@9468.4]
  assign Mem1D_5_io_w_data_0 = _T_505[16:9]; // @[MemPrimitives.scala 95:29:@9469.4]
  assign Mem1D_5_io_w_en_0 = _T_505[17]; // @[MemPrimitives.scala 96:27:@9470.4]
  assign Mem1D_6_clock = clock; // @[:@9240.4]
  assign Mem1D_6_reset = reset; // @[:@9241.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[8:0]; // @[MemPrimitives.scala 127:28:@10022.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[9]; // @[MemPrimitives.scala 128:32:@10023.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[8:0]; // @[MemPrimitives.scala 94:28:@9480.4]
  assign Mem1D_6_io_w_data_0 = _T_516[16:9]; // @[MemPrimitives.scala 95:29:@9481.4]
  assign Mem1D_6_io_w_en_0 = _T_516[17]; // @[MemPrimitives.scala 96:27:@9482.4]
  assign Mem1D_7_clock = clock; // @[:@9256.4]
  assign Mem1D_7_reset = reset; // @[:@9257.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[8:0]; // @[MemPrimitives.scala 127:28:@10084.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[9]; // @[MemPrimitives.scala 128:32:@10085.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[8:0]; // @[MemPrimitives.scala 94:28:@9492.4]
  assign Mem1D_7_io_w_data_0 = _T_527[16:9]; // @[MemPrimitives.scala 95:29:@9493.4]
  assign Mem1D_7_io_w_en_0 = _T_527[17]; // @[MemPrimitives.scala 96:27:@9494.4]
  assign Mem1D_8_clock = clock; // @[:@9272.4]
  assign Mem1D_8_reset = reset; // @[:@9273.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[8:0]; // @[MemPrimitives.scala 127:28:@10146.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[9]; // @[MemPrimitives.scala 128:32:@10147.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[8:0]; // @[MemPrimitives.scala 94:28:@9504.4]
  assign Mem1D_8_io_w_data_0 = _T_538[16:9]; // @[MemPrimitives.scala 95:29:@9505.4]
  assign Mem1D_8_io_w_en_0 = _T_538[17]; // @[MemPrimitives.scala 96:27:@9506.4]
  assign Mem1D_9_clock = clock; // @[:@9288.4]
  assign Mem1D_9_reset = reset; // @[:@9289.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[8:0]; // @[MemPrimitives.scala 127:28:@10208.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[9]; // @[MemPrimitives.scala 128:32:@10209.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[8:0]; // @[MemPrimitives.scala 94:28:@9516.4]
  assign Mem1D_9_io_w_data_0 = _T_549[16:9]; // @[MemPrimitives.scala 95:29:@9517.4]
  assign Mem1D_9_io_w_en_0 = _T_549[17]; // @[MemPrimitives.scala 96:27:@9518.4]
  assign Mem1D_10_clock = clock; // @[:@9304.4]
  assign Mem1D_10_reset = reset; // @[:@9305.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[8:0]; // @[MemPrimitives.scala 127:28:@10270.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[9]; // @[MemPrimitives.scala 128:32:@10271.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[8:0]; // @[MemPrimitives.scala 94:28:@9528.4]
  assign Mem1D_10_io_w_data_0 = _T_560[16:9]; // @[MemPrimitives.scala 95:29:@9529.4]
  assign Mem1D_10_io_w_en_0 = _T_560[17]; // @[MemPrimitives.scala 96:27:@9530.4]
  assign Mem1D_11_clock = clock; // @[:@9320.4]
  assign Mem1D_11_reset = reset; // @[:@9321.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 127:28:@10332.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 128:32:@10333.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[8:0]; // @[MemPrimitives.scala 94:28:@9540.4]
  assign Mem1D_11_io_w_data_0 = _T_571[16:9]; // @[MemPrimitives.scala 95:29:@9541.4]
  assign Mem1D_11_io_w_en_0 = _T_571[17]; // @[MemPrimitives.scala 96:27:@9542.4]
  assign Mem1D_12_clock = clock; // @[:@9336.4]
  assign Mem1D_12_reset = reset; // @[:@9337.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[8:0]; // @[MemPrimitives.scala 127:28:@10394.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[9]; // @[MemPrimitives.scala 128:32:@10395.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[8:0]; // @[MemPrimitives.scala 94:28:@9552.4]
  assign Mem1D_12_io_w_data_0 = _T_582[16:9]; // @[MemPrimitives.scala 95:29:@9553.4]
  assign Mem1D_12_io_w_en_0 = _T_582[17]; // @[MemPrimitives.scala 96:27:@9554.4]
  assign Mem1D_13_clock = clock; // @[:@9352.4]
  assign Mem1D_13_reset = reset; // @[:@9353.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[8:0]; // @[MemPrimitives.scala 127:28:@10456.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[9]; // @[MemPrimitives.scala 128:32:@10457.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[8:0]; // @[MemPrimitives.scala 94:28:@9564.4]
  assign Mem1D_13_io_w_data_0 = _T_593[16:9]; // @[MemPrimitives.scala 95:29:@9565.4]
  assign Mem1D_13_io_w_en_0 = _T_593[17]; // @[MemPrimitives.scala 96:27:@9566.4]
  assign Mem1D_14_clock = clock; // @[:@9368.4]
  assign Mem1D_14_reset = reset; // @[:@9369.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[8:0]; // @[MemPrimitives.scala 127:28:@10518.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[9]; // @[MemPrimitives.scala 128:32:@10519.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[8:0]; // @[MemPrimitives.scala 94:28:@9576.4]
  assign Mem1D_14_io_w_data_0 = _T_604[16:9]; // @[MemPrimitives.scala 95:29:@9577.4]
  assign Mem1D_14_io_w_en_0 = _T_604[17]; // @[MemPrimitives.scala 96:27:@9578.4]
  assign Mem1D_15_clock = clock; // @[:@9384.4]
  assign Mem1D_15_reset = reset; // @[:@9385.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[8:0]; // @[MemPrimitives.scala 127:28:@10580.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[9]; // @[MemPrimitives.scala 128:32:@10581.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@9588.4]
  assign Mem1D_15_io_w_data_0 = _T_615[16:9]; // @[MemPrimitives.scala 95:29:@9589.4]
  assign Mem1D_15_io_w_en_0 = _T_615[17]; // @[MemPrimitives.scala 96:27:@9590.4]
  assign StickySelects_clock = clock; // @[:@9616.4]
  assign StickySelects_reset = reset; // @[:@9617.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_623; // @[MemPrimitives.scala 122:60:@9618.4]
  assign StickySelects_io_ins_1 = io_rPort_2_en_0 & _T_629; // @[MemPrimitives.scala 122:60:@9619.4]
  assign StickySelects_io_ins_2 = io_rPort_4_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@9620.4]
  assign StickySelects_io_ins_3 = io_rPort_5_en_0 & _T_641; // @[MemPrimitives.scala 122:60:@9621.4]
  assign StickySelects_io_ins_4 = io_rPort_7_en_0 & _T_647; // @[MemPrimitives.scala 122:60:@9622.4]
  assign StickySelects_io_ins_5 = io_rPort_8_en_0 & _T_653; // @[MemPrimitives.scala 122:60:@9623.4]
  assign StickySelects_1_clock = clock; // @[:@9678.4]
  assign StickySelects_1_reset = reset; // @[:@9679.4]
  assign StickySelects_1_io_ins_0 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 122:60:@9680.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_691; // @[MemPrimitives.scala 122:60:@9681.4]
  assign StickySelects_1_io_ins_2 = io_rPort_6_en_0 & _T_697; // @[MemPrimitives.scala 122:60:@9682.4]
  assign StickySelects_1_io_ins_3 = io_rPort_9_en_0 & _T_703; // @[MemPrimitives.scala 122:60:@9683.4]
  assign StickySelects_1_io_ins_4 = io_rPort_10_en_0 & _T_709; // @[MemPrimitives.scala 122:60:@9684.4]
  assign StickySelects_1_io_ins_5 = io_rPort_11_en_0 & _T_715; // @[MemPrimitives.scala 122:60:@9685.4]
  assign StickySelects_2_clock = clock; // @[:@9740.4]
  assign StickySelects_2_reset = reset; // @[:@9741.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_747; // @[MemPrimitives.scala 122:60:@9742.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_753; // @[MemPrimitives.scala 122:60:@9743.4]
  assign StickySelects_2_io_ins_2 = io_rPort_4_en_0 & _T_759; // @[MemPrimitives.scala 122:60:@9744.4]
  assign StickySelects_2_io_ins_3 = io_rPort_5_en_0 & _T_765; // @[MemPrimitives.scala 122:60:@9745.4]
  assign StickySelects_2_io_ins_4 = io_rPort_7_en_0 & _T_771; // @[MemPrimitives.scala 122:60:@9746.4]
  assign StickySelects_2_io_ins_5 = io_rPort_8_en_0 & _T_777; // @[MemPrimitives.scala 122:60:@9747.4]
  assign StickySelects_3_clock = clock; // @[:@9802.4]
  assign StickySelects_3_reset = reset; // @[:@9803.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_809; // @[MemPrimitives.scala 122:60:@9804.4]
  assign StickySelects_3_io_ins_1 = io_rPort_3_en_0 & _T_815; // @[MemPrimitives.scala 122:60:@9805.4]
  assign StickySelects_3_io_ins_2 = io_rPort_6_en_0 & _T_821; // @[MemPrimitives.scala 122:60:@9806.4]
  assign StickySelects_3_io_ins_3 = io_rPort_9_en_0 & _T_827; // @[MemPrimitives.scala 122:60:@9807.4]
  assign StickySelects_3_io_ins_4 = io_rPort_10_en_0 & _T_833; // @[MemPrimitives.scala 122:60:@9808.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_839; // @[MemPrimitives.scala 122:60:@9809.4]
  assign StickySelects_4_clock = clock; // @[:@9864.4]
  assign StickySelects_4_reset = reset; // @[:@9865.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_871; // @[MemPrimitives.scala 122:60:@9866.4]
  assign StickySelects_4_io_ins_1 = io_rPort_2_en_0 & _T_877; // @[MemPrimitives.scala 122:60:@9867.4]
  assign StickySelects_4_io_ins_2 = io_rPort_4_en_0 & _T_883; // @[MemPrimitives.scala 122:60:@9868.4]
  assign StickySelects_4_io_ins_3 = io_rPort_5_en_0 & _T_889; // @[MemPrimitives.scala 122:60:@9869.4]
  assign StickySelects_4_io_ins_4 = io_rPort_7_en_0 & _T_895; // @[MemPrimitives.scala 122:60:@9870.4]
  assign StickySelects_4_io_ins_5 = io_rPort_8_en_0 & _T_901; // @[MemPrimitives.scala 122:60:@9871.4]
  assign StickySelects_5_clock = clock; // @[:@9926.4]
  assign StickySelects_5_reset = reset; // @[:@9927.4]
  assign StickySelects_5_io_ins_0 = io_rPort_1_en_0 & _T_933; // @[MemPrimitives.scala 122:60:@9928.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_939; // @[MemPrimitives.scala 122:60:@9929.4]
  assign StickySelects_5_io_ins_2 = io_rPort_6_en_0 & _T_945; // @[MemPrimitives.scala 122:60:@9930.4]
  assign StickySelects_5_io_ins_3 = io_rPort_9_en_0 & _T_951; // @[MemPrimitives.scala 122:60:@9931.4]
  assign StickySelects_5_io_ins_4 = io_rPort_10_en_0 & _T_957; // @[MemPrimitives.scala 122:60:@9932.4]
  assign StickySelects_5_io_ins_5 = io_rPort_11_en_0 & _T_963; // @[MemPrimitives.scala 122:60:@9933.4]
  assign StickySelects_6_clock = clock; // @[:@9988.4]
  assign StickySelects_6_reset = reset; // @[:@9989.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_995; // @[MemPrimitives.scala 122:60:@9990.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_1001; // @[MemPrimitives.scala 122:60:@9991.4]
  assign StickySelects_6_io_ins_2 = io_rPort_4_en_0 & _T_1007; // @[MemPrimitives.scala 122:60:@9992.4]
  assign StickySelects_6_io_ins_3 = io_rPort_5_en_0 & _T_1013; // @[MemPrimitives.scala 122:60:@9993.4]
  assign StickySelects_6_io_ins_4 = io_rPort_7_en_0 & _T_1019; // @[MemPrimitives.scala 122:60:@9994.4]
  assign StickySelects_6_io_ins_5 = io_rPort_8_en_0 & _T_1025; // @[MemPrimitives.scala 122:60:@9995.4]
  assign StickySelects_7_clock = clock; // @[:@10050.4]
  assign StickySelects_7_reset = reset; // @[:@10051.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1057; // @[MemPrimitives.scala 122:60:@10052.4]
  assign StickySelects_7_io_ins_1 = io_rPort_3_en_0 & _T_1063; // @[MemPrimitives.scala 122:60:@10053.4]
  assign StickySelects_7_io_ins_2 = io_rPort_6_en_0 & _T_1069; // @[MemPrimitives.scala 122:60:@10054.4]
  assign StickySelects_7_io_ins_3 = io_rPort_9_en_0 & _T_1075; // @[MemPrimitives.scala 122:60:@10055.4]
  assign StickySelects_7_io_ins_4 = io_rPort_10_en_0 & _T_1081; // @[MemPrimitives.scala 122:60:@10056.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1087; // @[MemPrimitives.scala 122:60:@10057.4]
  assign StickySelects_8_clock = clock; // @[:@10112.4]
  assign StickySelects_8_reset = reset; // @[:@10113.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1119; // @[MemPrimitives.scala 122:60:@10114.4]
  assign StickySelects_8_io_ins_1 = io_rPort_2_en_0 & _T_1125; // @[MemPrimitives.scala 122:60:@10115.4]
  assign StickySelects_8_io_ins_2 = io_rPort_4_en_0 & _T_1131; // @[MemPrimitives.scala 122:60:@10116.4]
  assign StickySelects_8_io_ins_3 = io_rPort_5_en_0 & _T_1137; // @[MemPrimitives.scala 122:60:@10117.4]
  assign StickySelects_8_io_ins_4 = io_rPort_7_en_0 & _T_1143; // @[MemPrimitives.scala 122:60:@10118.4]
  assign StickySelects_8_io_ins_5 = io_rPort_8_en_0 & _T_1149; // @[MemPrimitives.scala 122:60:@10119.4]
  assign StickySelects_9_clock = clock; // @[:@10174.4]
  assign StickySelects_9_reset = reset; // @[:@10175.4]
  assign StickySelects_9_io_ins_0 = io_rPort_1_en_0 & _T_1181; // @[MemPrimitives.scala 122:60:@10176.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_1187; // @[MemPrimitives.scala 122:60:@10177.4]
  assign StickySelects_9_io_ins_2 = io_rPort_6_en_0 & _T_1193; // @[MemPrimitives.scala 122:60:@10178.4]
  assign StickySelects_9_io_ins_3 = io_rPort_9_en_0 & _T_1199; // @[MemPrimitives.scala 122:60:@10179.4]
  assign StickySelects_9_io_ins_4 = io_rPort_10_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@10180.4]
  assign StickySelects_9_io_ins_5 = io_rPort_11_en_0 & _T_1211; // @[MemPrimitives.scala 122:60:@10181.4]
  assign StickySelects_10_clock = clock; // @[:@10236.4]
  assign StickySelects_10_reset = reset; // @[:@10237.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1243; // @[MemPrimitives.scala 122:60:@10238.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_1249; // @[MemPrimitives.scala 122:60:@10239.4]
  assign StickySelects_10_io_ins_2 = io_rPort_4_en_0 & _T_1255; // @[MemPrimitives.scala 122:60:@10240.4]
  assign StickySelects_10_io_ins_3 = io_rPort_5_en_0 & _T_1261; // @[MemPrimitives.scala 122:60:@10241.4]
  assign StickySelects_10_io_ins_4 = io_rPort_7_en_0 & _T_1267; // @[MemPrimitives.scala 122:60:@10242.4]
  assign StickySelects_10_io_ins_5 = io_rPort_8_en_0 & _T_1273; // @[MemPrimitives.scala 122:60:@10243.4]
  assign StickySelects_11_clock = clock; // @[:@10298.4]
  assign StickySelects_11_reset = reset; // @[:@10299.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1305; // @[MemPrimitives.scala 122:60:@10300.4]
  assign StickySelects_11_io_ins_1 = io_rPort_3_en_0 & _T_1311; // @[MemPrimitives.scala 122:60:@10301.4]
  assign StickySelects_11_io_ins_2 = io_rPort_6_en_0 & _T_1317; // @[MemPrimitives.scala 122:60:@10302.4]
  assign StickySelects_11_io_ins_3 = io_rPort_9_en_0 & _T_1323; // @[MemPrimitives.scala 122:60:@10303.4]
  assign StickySelects_11_io_ins_4 = io_rPort_10_en_0 & _T_1329; // @[MemPrimitives.scala 122:60:@10304.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@10305.4]
  assign StickySelects_12_clock = clock; // @[:@10360.4]
  assign StickySelects_12_reset = reset; // @[:@10361.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 122:60:@10362.4]
  assign StickySelects_12_io_ins_1 = io_rPort_2_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@10363.4]
  assign StickySelects_12_io_ins_2 = io_rPort_4_en_0 & _T_1379; // @[MemPrimitives.scala 122:60:@10364.4]
  assign StickySelects_12_io_ins_3 = io_rPort_5_en_0 & _T_1385; // @[MemPrimitives.scala 122:60:@10365.4]
  assign StickySelects_12_io_ins_4 = io_rPort_7_en_0 & _T_1391; // @[MemPrimitives.scala 122:60:@10366.4]
  assign StickySelects_12_io_ins_5 = io_rPort_8_en_0 & _T_1397; // @[MemPrimitives.scala 122:60:@10367.4]
  assign StickySelects_13_clock = clock; // @[:@10422.4]
  assign StickySelects_13_reset = reset; // @[:@10423.4]
  assign StickySelects_13_io_ins_0 = io_rPort_1_en_0 & _T_1429; // @[MemPrimitives.scala 122:60:@10424.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_1435; // @[MemPrimitives.scala 122:60:@10425.4]
  assign StickySelects_13_io_ins_2 = io_rPort_6_en_0 & _T_1441; // @[MemPrimitives.scala 122:60:@10426.4]
  assign StickySelects_13_io_ins_3 = io_rPort_9_en_0 & _T_1447; // @[MemPrimitives.scala 122:60:@10427.4]
  assign StickySelects_13_io_ins_4 = io_rPort_10_en_0 & _T_1453; // @[MemPrimitives.scala 122:60:@10428.4]
  assign StickySelects_13_io_ins_5 = io_rPort_11_en_0 & _T_1459; // @[MemPrimitives.scala 122:60:@10429.4]
  assign StickySelects_14_clock = clock; // @[:@10484.4]
  assign StickySelects_14_reset = reset; // @[:@10485.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_1491; // @[MemPrimitives.scala 122:60:@10486.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_1497; // @[MemPrimitives.scala 122:60:@10487.4]
  assign StickySelects_14_io_ins_2 = io_rPort_4_en_0 & _T_1503; // @[MemPrimitives.scala 122:60:@10488.4]
  assign StickySelects_14_io_ins_3 = io_rPort_5_en_0 & _T_1509; // @[MemPrimitives.scala 122:60:@10489.4]
  assign StickySelects_14_io_ins_4 = io_rPort_7_en_0 & _T_1515; // @[MemPrimitives.scala 122:60:@10490.4]
  assign StickySelects_14_io_ins_5 = io_rPort_8_en_0 & _T_1521; // @[MemPrimitives.scala 122:60:@10491.4]
  assign StickySelects_15_clock = clock; // @[:@10546.4]
  assign StickySelects_15_reset = reset; // @[:@10547.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_1553; // @[MemPrimitives.scala 122:60:@10548.4]
  assign StickySelects_15_io_ins_1 = io_rPort_3_en_0 & _T_1559; // @[MemPrimitives.scala 122:60:@10549.4]
  assign StickySelects_15_io_ins_2 = io_rPort_6_en_0 & _T_1565; // @[MemPrimitives.scala 122:60:@10550.4]
  assign StickySelects_15_io_ins_3 = io_rPort_9_en_0 & _T_1571; // @[MemPrimitives.scala 122:60:@10551.4]
  assign StickySelects_15_io_ins_4 = io_rPort_10_en_0 & _T_1577; // @[MemPrimitives.scala 122:60:@10552.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_1583; // @[MemPrimitives.scala 122:60:@10553.4]
  assign RetimeWrapper_clock = clock; // @[:@10609.4]
  assign RetimeWrapper_reset = reset; // @[:@10610.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10612.4]
  assign RetimeWrapper_io_in = _T_623 & io_rPort_0_en_0; // @[package.scala 94:16:@10611.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10617.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10618.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10620.4]
  assign RetimeWrapper_1_io_in = _T_747 & io_rPort_0_en_0; // @[package.scala 94:16:@10619.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10625.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10626.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10628.4]
  assign RetimeWrapper_2_io_in = _T_871 & io_rPort_0_en_0; // @[package.scala 94:16:@10627.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10633.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10634.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10636.4]
  assign RetimeWrapper_3_io_in = _T_995 & io_rPort_0_en_0; // @[package.scala 94:16:@10635.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10641.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10642.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10644.4]
  assign RetimeWrapper_4_io_in = _T_1119 & io_rPort_0_en_0; // @[package.scala 94:16:@10643.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10649.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10650.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10652.4]
  assign RetimeWrapper_5_io_in = _T_1243 & io_rPort_0_en_0; // @[package.scala 94:16:@10651.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10657.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10658.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10660.4]
  assign RetimeWrapper_6_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@10659.4]
  assign RetimeWrapper_7_clock = clock; // @[:@10665.4]
  assign RetimeWrapper_7_reset = reset; // @[:@10666.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10668.4]
  assign RetimeWrapper_7_io_in = _T_1491 & io_rPort_0_en_0; // @[package.scala 94:16:@10667.4]
  assign RetimeWrapper_8_clock = clock; // @[:@10705.4]
  assign RetimeWrapper_8_reset = reset; // @[:@10706.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10708.4]
  assign RetimeWrapper_8_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@10707.4]
  assign RetimeWrapper_9_clock = clock; // @[:@10713.4]
  assign RetimeWrapper_9_reset = reset; // @[:@10714.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10716.4]
  assign RetimeWrapper_9_io_in = _T_809 & io_rPort_1_en_0; // @[package.scala 94:16:@10715.4]
  assign RetimeWrapper_10_clock = clock; // @[:@10721.4]
  assign RetimeWrapper_10_reset = reset; // @[:@10722.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10724.4]
  assign RetimeWrapper_10_io_in = _T_933 & io_rPort_1_en_0; // @[package.scala 94:16:@10723.4]
  assign RetimeWrapper_11_clock = clock; // @[:@10729.4]
  assign RetimeWrapper_11_reset = reset; // @[:@10730.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10732.4]
  assign RetimeWrapper_11_io_in = _T_1057 & io_rPort_1_en_0; // @[package.scala 94:16:@10731.4]
  assign RetimeWrapper_12_clock = clock; // @[:@10737.4]
  assign RetimeWrapper_12_reset = reset; // @[:@10738.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10740.4]
  assign RetimeWrapper_12_io_in = _T_1181 & io_rPort_1_en_0; // @[package.scala 94:16:@10739.4]
  assign RetimeWrapper_13_clock = clock; // @[:@10745.4]
  assign RetimeWrapper_13_reset = reset; // @[:@10746.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10748.4]
  assign RetimeWrapper_13_io_in = _T_1305 & io_rPort_1_en_0; // @[package.scala 94:16:@10747.4]
  assign RetimeWrapper_14_clock = clock; // @[:@10753.4]
  assign RetimeWrapper_14_reset = reset; // @[:@10754.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10756.4]
  assign RetimeWrapper_14_io_in = _T_1429 & io_rPort_1_en_0; // @[package.scala 94:16:@10755.4]
  assign RetimeWrapper_15_clock = clock; // @[:@10761.4]
  assign RetimeWrapper_15_reset = reset; // @[:@10762.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10764.4]
  assign RetimeWrapper_15_io_in = _T_1553 & io_rPort_1_en_0; // @[package.scala 94:16:@10763.4]
  assign RetimeWrapper_16_clock = clock; // @[:@10801.4]
  assign RetimeWrapper_16_reset = reset; // @[:@10802.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10804.4]
  assign RetimeWrapper_16_io_in = _T_629 & io_rPort_2_en_0; // @[package.scala 94:16:@10803.4]
  assign RetimeWrapper_17_clock = clock; // @[:@10809.4]
  assign RetimeWrapper_17_reset = reset; // @[:@10810.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10812.4]
  assign RetimeWrapper_17_io_in = _T_753 & io_rPort_2_en_0; // @[package.scala 94:16:@10811.4]
  assign RetimeWrapper_18_clock = clock; // @[:@10817.4]
  assign RetimeWrapper_18_reset = reset; // @[:@10818.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10820.4]
  assign RetimeWrapper_18_io_in = _T_877 & io_rPort_2_en_0; // @[package.scala 94:16:@10819.4]
  assign RetimeWrapper_19_clock = clock; // @[:@10825.4]
  assign RetimeWrapper_19_reset = reset; // @[:@10826.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10828.4]
  assign RetimeWrapper_19_io_in = _T_1001 & io_rPort_2_en_0; // @[package.scala 94:16:@10827.4]
  assign RetimeWrapper_20_clock = clock; // @[:@10833.4]
  assign RetimeWrapper_20_reset = reset; // @[:@10834.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10836.4]
  assign RetimeWrapper_20_io_in = _T_1125 & io_rPort_2_en_0; // @[package.scala 94:16:@10835.4]
  assign RetimeWrapper_21_clock = clock; // @[:@10841.4]
  assign RetimeWrapper_21_reset = reset; // @[:@10842.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10844.4]
  assign RetimeWrapper_21_io_in = _T_1249 & io_rPort_2_en_0; // @[package.scala 94:16:@10843.4]
  assign RetimeWrapper_22_clock = clock; // @[:@10849.4]
  assign RetimeWrapper_22_reset = reset; // @[:@10850.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10852.4]
  assign RetimeWrapper_22_io_in = _T_1373 & io_rPort_2_en_0; // @[package.scala 94:16:@10851.4]
  assign RetimeWrapper_23_clock = clock; // @[:@10857.4]
  assign RetimeWrapper_23_reset = reset; // @[:@10858.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10860.4]
  assign RetimeWrapper_23_io_in = _T_1497 & io_rPort_2_en_0; // @[package.scala 94:16:@10859.4]
  assign RetimeWrapper_24_clock = clock; // @[:@10897.4]
  assign RetimeWrapper_24_reset = reset; // @[:@10898.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10900.4]
  assign RetimeWrapper_24_io_in = _T_691 & io_rPort_3_en_0; // @[package.scala 94:16:@10899.4]
  assign RetimeWrapper_25_clock = clock; // @[:@10905.4]
  assign RetimeWrapper_25_reset = reset; // @[:@10906.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10908.4]
  assign RetimeWrapper_25_io_in = _T_815 & io_rPort_3_en_0; // @[package.scala 94:16:@10907.4]
  assign RetimeWrapper_26_clock = clock; // @[:@10913.4]
  assign RetimeWrapper_26_reset = reset; // @[:@10914.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10916.4]
  assign RetimeWrapper_26_io_in = _T_939 & io_rPort_3_en_0; // @[package.scala 94:16:@10915.4]
  assign RetimeWrapper_27_clock = clock; // @[:@10921.4]
  assign RetimeWrapper_27_reset = reset; // @[:@10922.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10924.4]
  assign RetimeWrapper_27_io_in = _T_1063 & io_rPort_3_en_0; // @[package.scala 94:16:@10923.4]
  assign RetimeWrapper_28_clock = clock; // @[:@10929.4]
  assign RetimeWrapper_28_reset = reset; // @[:@10930.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10932.4]
  assign RetimeWrapper_28_io_in = _T_1187 & io_rPort_3_en_0; // @[package.scala 94:16:@10931.4]
  assign RetimeWrapper_29_clock = clock; // @[:@10937.4]
  assign RetimeWrapper_29_reset = reset; // @[:@10938.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10940.4]
  assign RetimeWrapper_29_io_in = _T_1311 & io_rPort_3_en_0; // @[package.scala 94:16:@10939.4]
  assign RetimeWrapper_30_clock = clock; // @[:@10945.4]
  assign RetimeWrapper_30_reset = reset; // @[:@10946.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10948.4]
  assign RetimeWrapper_30_io_in = _T_1435 & io_rPort_3_en_0; // @[package.scala 94:16:@10947.4]
  assign RetimeWrapper_31_clock = clock; // @[:@10953.4]
  assign RetimeWrapper_31_reset = reset; // @[:@10954.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10956.4]
  assign RetimeWrapper_31_io_in = _T_1559 & io_rPort_3_en_0; // @[package.scala 94:16:@10955.4]
  assign RetimeWrapper_32_clock = clock; // @[:@10993.4]
  assign RetimeWrapper_32_reset = reset; // @[:@10994.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10996.4]
  assign RetimeWrapper_32_io_in = _T_635 & io_rPort_4_en_0; // @[package.scala 94:16:@10995.4]
  assign RetimeWrapper_33_clock = clock; // @[:@11001.4]
  assign RetimeWrapper_33_reset = reset; // @[:@11002.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11004.4]
  assign RetimeWrapper_33_io_in = _T_759 & io_rPort_4_en_0; // @[package.scala 94:16:@11003.4]
  assign RetimeWrapper_34_clock = clock; // @[:@11009.4]
  assign RetimeWrapper_34_reset = reset; // @[:@11010.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11012.4]
  assign RetimeWrapper_34_io_in = _T_883 & io_rPort_4_en_0; // @[package.scala 94:16:@11011.4]
  assign RetimeWrapper_35_clock = clock; // @[:@11017.4]
  assign RetimeWrapper_35_reset = reset; // @[:@11018.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11020.4]
  assign RetimeWrapper_35_io_in = _T_1007 & io_rPort_4_en_0; // @[package.scala 94:16:@11019.4]
  assign RetimeWrapper_36_clock = clock; // @[:@11025.4]
  assign RetimeWrapper_36_reset = reset; // @[:@11026.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11028.4]
  assign RetimeWrapper_36_io_in = _T_1131 & io_rPort_4_en_0; // @[package.scala 94:16:@11027.4]
  assign RetimeWrapper_37_clock = clock; // @[:@11033.4]
  assign RetimeWrapper_37_reset = reset; // @[:@11034.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11036.4]
  assign RetimeWrapper_37_io_in = _T_1255 & io_rPort_4_en_0; // @[package.scala 94:16:@11035.4]
  assign RetimeWrapper_38_clock = clock; // @[:@11041.4]
  assign RetimeWrapper_38_reset = reset; // @[:@11042.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11044.4]
  assign RetimeWrapper_38_io_in = _T_1379 & io_rPort_4_en_0; // @[package.scala 94:16:@11043.4]
  assign RetimeWrapper_39_clock = clock; // @[:@11049.4]
  assign RetimeWrapper_39_reset = reset; // @[:@11050.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@11052.4]
  assign RetimeWrapper_39_io_in = _T_1503 & io_rPort_4_en_0; // @[package.scala 94:16:@11051.4]
  assign RetimeWrapper_40_clock = clock; // @[:@11089.4]
  assign RetimeWrapper_40_reset = reset; // @[:@11090.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11092.4]
  assign RetimeWrapper_40_io_in = _T_641 & io_rPort_5_en_0; // @[package.scala 94:16:@11091.4]
  assign RetimeWrapper_41_clock = clock; // @[:@11097.4]
  assign RetimeWrapper_41_reset = reset; // @[:@11098.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11100.4]
  assign RetimeWrapper_41_io_in = _T_765 & io_rPort_5_en_0; // @[package.scala 94:16:@11099.4]
  assign RetimeWrapper_42_clock = clock; // @[:@11105.4]
  assign RetimeWrapper_42_reset = reset; // @[:@11106.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11108.4]
  assign RetimeWrapper_42_io_in = _T_889 & io_rPort_5_en_0; // @[package.scala 94:16:@11107.4]
  assign RetimeWrapper_43_clock = clock; // @[:@11113.4]
  assign RetimeWrapper_43_reset = reset; // @[:@11114.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11116.4]
  assign RetimeWrapper_43_io_in = _T_1013 & io_rPort_5_en_0; // @[package.scala 94:16:@11115.4]
  assign RetimeWrapper_44_clock = clock; // @[:@11121.4]
  assign RetimeWrapper_44_reset = reset; // @[:@11122.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11124.4]
  assign RetimeWrapper_44_io_in = _T_1137 & io_rPort_5_en_0; // @[package.scala 94:16:@11123.4]
  assign RetimeWrapper_45_clock = clock; // @[:@11129.4]
  assign RetimeWrapper_45_reset = reset; // @[:@11130.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11132.4]
  assign RetimeWrapper_45_io_in = _T_1261 & io_rPort_5_en_0; // @[package.scala 94:16:@11131.4]
  assign RetimeWrapper_46_clock = clock; // @[:@11137.4]
  assign RetimeWrapper_46_reset = reset; // @[:@11138.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11140.4]
  assign RetimeWrapper_46_io_in = _T_1385 & io_rPort_5_en_0; // @[package.scala 94:16:@11139.4]
  assign RetimeWrapper_47_clock = clock; // @[:@11145.4]
  assign RetimeWrapper_47_reset = reset; // @[:@11146.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11148.4]
  assign RetimeWrapper_47_io_in = _T_1509 & io_rPort_5_en_0; // @[package.scala 94:16:@11147.4]
  assign RetimeWrapper_48_clock = clock; // @[:@11185.4]
  assign RetimeWrapper_48_reset = reset; // @[:@11186.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11188.4]
  assign RetimeWrapper_48_io_in = _T_697 & io_rPort_6_en_0; // @[package.scala 94:16:@11187.4]
  assign RetimeWrapper_49_clock = clock; // @[:@11193.4]
  assign RetimeWrapper_49_reset = reset; // @[:@11194.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11196.4]
  assign RetimeWrapper_49_io_in = _T_821 & io_rPort_6_en_0; // @[package.scala 94:16:@11195.4]
  assign RetimeWrapper_50_clock = clock; // @[:@11201.4]
  assign RetimeWrapper_50_reset = reset; // @[:@11202.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11204.4]
  assign RetimeWrapper_50_io_in = _T_945 & io_rPort_6_en_0; // @[package.scala 94:16:@11203.4]
  assign RetimeWrapper_51_clock = clock; // @[:@11209.4]
  assign RetimeWrapper_51_reset = reset; // @[:@11210.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11212.4]
  assign RetimeWrapper_51_io_in = _T_1069 & io_rPort_6_en_0; // @[package.scala 94:16:@11211.4]
  assign RetimeWrapper_52_clock = clock; // @[:@11217.4]
  assign RetimeWrapper_52_reset = reset; // @[:@11218.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11220.4]
  assign RetimeWrapper_52_io_in = _T_1193 & io_rPort_6_en_0; // @[package.scala 94:16:@11219.4]
  assign RetimeWrapper_53_clock = clock; // @[:@11225.4]
  assign RetimeWrapper_53_reset = reset; // @[:@11226.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11228.4]
  assign RetimeWrapper_53_io_in = _T_1317 & io_rPort_6_en_0; // @[package.scala 94:16:@11227.4]
  assign RetimeWrapper_54_clock = clock; // @[:@11233.4]
  assign RetimeWrapper_54_reset = reset; // @[:@11234.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11236.4]
  assign RetimeWrapper_54_io_in = _T_1441 & io_rPort_6_en_0; // @[package.scala 94:16:@11235.4]
  assign RetimeWrapper_55_clock = clock; // @[:@11241.4]
  assign RetimeWrapper_55_reset = reset; // @[:@11242.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11244.4]
  assign RetimeWrapper_55_io_in = _T_1565 & io_rPort_6_en_0; // @[package.scala 94:16:@11243.4]
  assign RetimeWrapper_56_clock = clock; // @[:@11281.4]
  assign RetimeWrapper_56_reset = reset; // @[:@11282.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11284.4]
  assign RetimeWrapper_56_io_in = _T_647 & io_rPort_7_en_0; // @[package.scala 94:16:@11283.4]
  assign RetimeWrapper_57_clock = clock; // @[:@11289.4]
  assign RetimeWrapper_57_reset = reset; // @[:@11290.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11292.4]
  assign RetimeWrapper_57_io_in = _T_771 & io_rPort_7_en_0; // @[package.scala 94:16:@11291.4]
  assign RetimeWrapper_58_clock = clock; // @[:@11297.4]
  assign RetimeWrapper_58_reset = reset; // @[:@11298.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11300.4]
  assign RetimeWrapper_58_io_in = _T_895 & io_rPort_7_en_0; // @[package.scala 94:16:@11299.4]
  assign RetimeWrapper_59_clock = clock; // @[:@11305.4]
  assign RetimeWrapper_59_reset = reset; // @[:@11306.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11308.4]
  assign RetimeWrapper_59_io_in = _T_1019 & io_rPort_7_en_0; // @[package.scala 94:16:@11307.4]
  assign RetimeWrapper_60_clock = clock; // @[:@11313.4]
  assign RetimeWrapper_60_reset = reset; // @[:@11314.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11316.4]
  assign RetimeWrapper_60_io_in = _T_1143 & io_rPort_7_en_0; // @[package.scala 94:16:@11315.4]
  assign RetimeWrapper_61_clock = clock; // @[:@11321.4]
  assign RetimeWrapper_61_reset = reset; // @[:@11322.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11324.4]
  assign RetimeWrapper_61_io_in = _T_1267 & io_rPort_7_en_0; // @[package.scala 94:16:@11323.4]
  assign RetimeWrapper_62_clock = clock; // @[:@11329.4]
  assign RetimeWrapper_62_reset = reset; // @[:@11330.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11332.4]
  assign RetimeWrapper_62_io_in = _T_1391 & io_rPort_7_en_0; // @[package.scala 94:16:@11331.4]
  assign RetimeWrapper_63_clock = clock; // @[:@11337.4]
  assign RetimeWrapper_63_reset = reset; // @[:@11338.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11340.4]
  assign RetimeWrapper_63_io_in = _T_1515 & io_rPort_7_en_0; // @[package.scala 94:16:@11339.4]
  assign RetimeWrapper_64_clock = clock; // @[:@11377.4]
  assign RetimeWrapper_64_reset = reset; // @[:@11378.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11380.4]
  assign RetimeWrapper_64_io_in = _T_653 & io_rPort_8_en_0; // @[package.scala 94:16:@11379.4]
  assign RetimeWrapper_65_clock = clock; // @[:@11385.4]
  assign RetimeWrapper_65_reset = reset; // @[:@11386.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11388.4]
  assign RetimeWrapper_65_io_in = _T_777 & io_rPort_8_en_0; // @[package.scala 94:16:@11387.4]
  assign RetimeWrapper_66_clock = clock; // @[:@11393.4]
  assign RetimeWrapper_66_reset = reset; // @[:@11394.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11396.4]
  assign RetimeWrapper_66_io_in = _T_901 & io_rPort_8_en_0; // @[package.scala 94:16:@11395.4]
  assign RetimeWrapper_67_clock = clock; // @[:@11401.4]
  assign RetimeWrapper_67_reset = reset; // @[:@11402.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11404.4]
  assign RetimeWrapper_67_io_in = _T_1025 & io_rPort_8_en_0; // @[package.scala 94:16:@11403.4]
  assign RetimeWrapper_68_clock = clock; // @[:@11409.4]
  assign RetimeWrapper_68_reset = reset; // @[:@11410.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11412.4]
  assign RetimeWrapper_68_io_in = _T_1149 & io_rPort_8_en_0; // @[package.scala 94:16:@11411.4]
  assign RetimeWrapper_69_clock = clock; // @[:@11417.4]
  assign RetimeWrapper_69_reset = reset; // @[:@11418.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11420.4]
  assign RetimeWrapper_69_io_in = _T_1273 & io_rPort_8_en_0; // @[package.scala 94:16:@11419.4]
  assign RetimeWrapper_70_clock = clock; // @[:@11425.4]
  assign RetimeWrapper_70_reset = reset; // @[:@11426.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11428.4]
  assign RetimeWrapper_70_io_in = _T_1397 & io_rPort_8_en_0; // @[package.scala 94:16:@11427.4]
  assign RetimeWrapper_71_clock = clock; // @[:@11433.4]
  assign RetimeWrapper_71_reset = reset; // @[:@11434.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11436.4]
  assign RetimeWrapper_71_io_in = _T_1521 & io_rPort_8_en_0; // @[package.scala 94:16:@11435.4]
  assign RetimeWrapper_72_clock = clock; // @[:@11473.4]
  assign RetimeWrapper_72_reset = reset; // @[:@11474.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11476.4]
  assign RetimeWrapper_72_io_in = _T_703 & io_rPort_9_en_0; // @[package.scala 94:16:@11475.4]
  assign RetimeWrapper_73_clock = clock; // @[:@11481.4]
  assign RetimeWrapper_73_reset = reset; // @[:@11482.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11484.4]
  assign RetimeWrapper_73_io_in = _T_827 & io_rPort_9_en_0; // @[package.scala 94:16:@11483.4]
  assign RetimeWrapper_74_clock = clock; // @[:@11489.4]
  assign RetimeWrapper_74_reset = reset; // @[:@11490.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11492.4]
  assign RetimeWrapper_74_io_in = _T_951 & io_rPort_9_en_0; // @[package.scala 94:16:@11491.4]
  assign RetimeWrapper_75_clock = clock; // @[:@11497.4]
  assign RetimeWrapper_75_reset = reset; // @[:@11498.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11500.4]
  assign RetimeWrapper_75_io_in = _T_1075 & io_rPort_9_en_0; // @[package.scala 94:16:@11499.4]
  assign RetimeWrapper_76_clock = clock; // @[:@11505.4]
  assign RetimeWrapper_76_reset = reset; // @[:@11506.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11508.4]
  assign RetimeWrapper_76_io_in = _T_1199 & io_rPort_9_en_0; // @[package.scala 94:16:@11507.4]
  assign RetimeWrapper_77_clock = clock; // @[:@11513.4]
  assign RetimeWrapper_77_reset = reset; // @[:@11514.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11516.4]
  assign RetimeWrapper_77_io_in = _T_1323 & io_rPort_9_en_0; // @[package.scala 94:16:@11515.4]
  assign RetimeWrapper_78_clock = clock; // @[:@11521.4]
  assign RetimeWrapper_78_reset = reset; // @[:@11522.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11524.4]
  assign RetimeWrapper_78_io_in = _T_1447 & io_rPort_9_en_0; // @[package.scala 94:16:@11523.4]
  assign RetimeWrapper_79_clock = clock; // @[:@11529.4]
  assign RetimeWrapper_79_reset = reset; // @[:@11530.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11532.4]
  assign RetimeWrapper_79_io_in = _T_1571 & io_rPort_9_en_0; // @[package.scala 94:16:@11531.4]
  assign RetimeWrapper_80_clock = clock; // @[:@11569.4]
  assign RetimeWrapper_80_reset = reset; // @[:@11570.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11572.4]
  assign RetimeWrapper_80_io_in = _T_709 & io_rPort_10_en_0; // @[package.scala 94:16:@11571.4]
  assign RetimeWrapper_81_clock = clock; // @[:@11577.4]
  assign RetimeWrapper_81_reset = reset; // @[:@11578.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11580.4]
  assign RetimeWrapper_81_io_in = _T_833 & io_rPort_10_en_0; // @[package.scala 94:16:@11579.4]
  assign RetimeWrapper_82_clock = clock; // @[:@11585.4]
  assign RetimeWrapper_82_reset = reset; // @[:@11586.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11588.4]
  assign RetimeWrapper_82_io_in = _T_957 & io_rPort_10_en_0; // @[package.scala 94:16:@11587.4]
  assign RetimeWrapper_83_clock = clock; // @[:@11593.4]
  assign RetimeWrapper_83_reset = reset; // @[:@11594.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11596.4]
  assign RetimeWrapper_83_io_in = _T_1081 & io_rPort_10_en_0; // @[package.scala 94:16:@11595.4]
  assign RetimeWrapper_84_clock = clock; // @[:@11601.4]
  assign RetimeWrapper_84_reset = reset; // @[:@11602.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11604.4]
  assign RetimeWrapper_84_io_in = _T_1205 & io_rPort_10_en_0; // @[package.scala 94:16:@11603.4]
  assign RetimeWrapper_85_clock = clock; // @[:@11609.4]
  assign RetimeWrapper_85_reset = reset; // @[:@11610.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11612.4]
  assign RetimeWrapper_85_io_in = _T_1329 & io_rPort_10_en_0; // @[package.scala 94:16:@11611.4]
  assign RetimeWrapper_86_clock = clock; // @[:@11617.4]
  assign RetimeWrapper_86_reset = reset; // @[:@11618.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11620.4]
  assign RetimeWrapper_86_io_in = _T_1453 & io_rPort_10_en_0; // @[package.scala 94:16:@11619.4]
  assign RetimeWrapper_87_clock = clock; // @[:@11625.4]
  assign RetimeWrapper_87_reset = reset; // @[:@11626.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11628.4]
  assign RetimeWrapper_87_io_in = _T_1577 & io_rPort_10_en_0; // @[package.scala 94:16:@11627.4]
  assign RetimeWrapper_88_clock = clock; // @[:@11665.4]
  assign RetimeWrapper_88_reset = reset; // @[:@11666.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11668.4]
  assign RetimeWrapper_88_io_in = _T_715 & io_rPort_11_en_0; // @[package.scala 94:16:@11667.4]
  assign RetimeWrapper_89_clock = clock; // @[:@11673.4]
  assign RetimeWrapper_89_reset = reset; // @[:@11674.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11676.4]
  assign RetimeWrapper_89_io_in = _T_839 & io_rPort_11_en_0; // @[package.scala 94:16:@11675.4]
  assign RetimeWrapper_90_clock = clock; // @[:@11681.4]
  assign RetimeWrapper_90_reset = reset; // @[:@11682.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11684.4]
  assign RetimeWrapper_90_io_in = _T_963 & io_rPort_11_en_0; // @[package.scala 94:16:@11683.4]
  assign RetimeWrapper_91_clock = clock; // @[:@11689.4]
  assign RetimeWrapper_91_reset = reset; // @[:@11690.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11692.4]
  assign RetimeWrapper_91_io_in = _T_1087 & io_rPort_11_en_0; // @[package.scala 94:16:@11691.4]
  assign RetimeWrapper_92_clock = clock; // @[:@11697.4]
  assign RetimeWrapper_92_reset = reset; // @[:@11698.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11700.4]
  assign RetimeWrapper_92_io_in = _T_1211 & io_rPort_11_en_0; // @[package.scala 94:16:@11699.4]
  assign RetimeWrapper_93_clock = clock; // @[:@11705.4]
  assign RetimeWrapper_93_reset = reset; // @[:@11706.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11708.4]
  assign RetimeWrapper_93_io_in = _T_1335 & io_rPort_11_en_0; // @[package.scala 94:16:@11707.4]
  assign RetimeWrapper_94_clock = clock; // @[:@11713.4]
  assign RetimeWrapper_94_reset = reset; // @[:@11714.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11716.4]
  assign RetimeWrapper_94_io_in = _T_1459 & io_rPort_11_en_0; // @[package.scala 94:16:@11715.4]
  assign RetimeWrapper_95_clock = clock; // @[:@11721.4]
  assign RetimeWrapper_95_reset = reset; // @[:@11722.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11724.4]
  assign RetimeWrapper_95_io_in = _T_1583 & io_rPort_11_en_0; // @[package.scala 94:16:@11723.4]
endmodule
module RetimeWrapper_132( // @[:@11748.2]
  input         clock, // @[:@11749.4]
  input         reset, // @[:@11750.4]
  input         io_flow, // @[:@11751.4]
  input  [15:0] io_in, // @[:@11751.4]
  output [15:0] io_out // @[:@11751.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11753.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11753.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11753.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11753.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11753.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11753.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11753.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11766.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11765.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@11764.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11763.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11762.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11760.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@11768.2]
  input  [31:0] io_a, // @[:@11771.4]
  output [32:0] io_b // @[:@11771.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@11781.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@11781.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@11786.4]
endmodule
module __2( // @[:@11788.2]
  input  [31:0] io_b, // @[:@11791.4]
  output [32:0] io_result // @[:@11791.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@11796.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@11796.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@11796.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@11809.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@11804.4]
endmodule
module RetimeWrapper_133( // @[:@11866.2]
  input         clock, // @[:@11867.4]
  input         reset, // @[:@11868.4]
  input         io_flow, // @[:@11869.4]
  input  [31:0] io_in, // @[:@11869.4]
  output [31:0] io_out // @[:@11869.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11871.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11871.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11871.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11871.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11871.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11871.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11871.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11884.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11883.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@11882.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11881.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11880.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11878.4]
endmodule
module fix2fixBox( // @[:@11886.2]
  input         clock, // @[:@11887.4]
  input         reset, // @[:@11888.4]
  input  [32:0] io_a, // @[:@11889.4]
  input         io_flow, // @[:@11889.4]
  output [31:0] io_b // @[:@11889.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@11902.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@11902.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@11902.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@11902.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@11902.4]
  RetimeWrapper_133 RetimeWrapper ( // @[package.scala 93:22:@11902.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@11909.4]
  assign RetimeWrapper_clock = clock; // @[:@11903.4]
  assign RetimeWrapper_reset = reset; // @[:@11904.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@11906.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@11905.4]
endmodule
module x272_sum( // @[:@11911.2]
  input         clock, // @[:@11912.4]
  input         reset, // @[:@11913.4]
  input  [31:0] io_a, // @[:@11914.4]
  input  [31:0] io_b, // @[:@11914.4]
  input         io_flow, // @[:@11914.4]
  output [31:0] io_result // @[:@11914.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@11922.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@11922.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@11929.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@11929.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@11947.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@11947.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@11947.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@11947.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@11947.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@11927.4 Math.scala 713:14:@11928.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@11934.4 Math.scala 713:14:@11935.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@11936.4]
  __2 _ ( // @[Math.scala 709:24:@11922.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@11929.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@11947.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@11927.4 Math.scala 713:14:@11928.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@11934.4 Math.scala 713:14:@11935.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@11936.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@11955.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@11925.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@11932.4]
  assign fix2fixBox_clock = clock; // @[:@11948.4]
  assign fix2fixBox_reset = reset; // @[:@11949.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@11950.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@11953.4]
endmodule
module RetimeWrapper_134( // @[:@11969.2]
  input         clock, // @[:@11970.4]
  input         reset, // @[:@11971.4]
  input         io_flow, // @[:@11972.4]
  input  [31:0] io_in, // @[:@11972.4]
  output [31:0] io_out // @[:@11972.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11974.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11974.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11974.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11974.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11974.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11974.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@11974.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11987.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11986.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@11985.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11984.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11983.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11981.4]
endmodule
module RetimeWrapper_136( // @[:@12033.2]
  input        clock, // @[:@12034.4]
  input        reset, // @[:@12035.4]
  input        io_flow, // @[:@12036.4]
  input  [7:0] io_in, // @[:@12036.4]
  output [7:0] io_out // @[:@12036.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12038.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12038.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12038.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12038.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12038.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12038.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@12038.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12051.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12050.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@12049.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12048.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12047.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12045.4]
endmodule
module RetimeWrapper_147( // @[:@12699.2]
  input         clock, // @[:@12700.4]
  input         reset, // @[:@12701.4]
  input         io_flow, // @[:@12702.4]
  input  [31:0] io_in, // @[:@12702.4]
  output [31:0] io_out // @[:@12702.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12704.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12704.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12704.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12704.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12704.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12704.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@12704.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12717.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12716.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12715.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12714.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12713.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12711.4]
endmodule
module RetimeWrapper_148( // @[:@12731.2]
  input         clock, // @[:@12732.4]
  input         reset, // @[:@12733.4]
  input         io_flow, // @[:@12734.4]
  input  [31:0] io_in, // @[:@12734.4]
  output [31:0] io_out // @[:@12734.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12736.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12736.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12736.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12736.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12736.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12736.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@12736.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12749.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12748.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12747.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12746.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12745.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12743.4]
endmodule
module fix2fixBox_3( // @[:@12751.2]
  input  [63:0] io_a, // @[:@12754.4]
  output [31:0] io_b // @[:@12754.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@12767.4]
endmodule
module x281( // @[:@12769.2]
  input         clock, // @[:@12770.4]
  input         reset, // @[:@12771.4]
  input  [31:0] io_a, // @[:@12772.4]
  input         io_flow, // @[:@12772.4]
  output [31:0] io_result // @[:@12772.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@12781.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@12781.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@12781.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@12781.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@12781.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@12789.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@12789.4]
  wire [31:0] _T_19; // @[package.scala 96:25:@12786.4 package.scala 96:25:@12787.4]
  wire [31:0] _GEN_0; // @[package.scala 94:16:@12784.4]
  RetimeWrapper_148 RetimeWrapper ( // @[package.scala 93:22:@12781.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  fix2fixBox_3 fix2fixBox ( // @[Math.scala 357:30:@12789.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_19 = RetimeWrapper_io_out; // @[package.scala 96:25:@12786.4 package.scala 96:25:@12787.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@12797.4]
  assign RetimeWrapper_clock = clock; // @[:@12782.4]
  assign RetimeWrapper_reset = reset; // @[:@12783.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@12785.4]
  assign _GEN_0 = io_a % 32'h780; // @[package.scala 94:16:@12784.4]
  assign RetimeWrapper_io_in = _GEN_0[31:0]; // @[package.scala 94:16:@12784.4]
  assign fix2fixBox_io_a = {{32'd0}, _T_19}; // @[Math.scala 358:23:@12792.4]
endmodule
module RetimeWrapper_151( // @[:@12875.2]
  input         clock, // @[:@12876.4]
  input         reset, // @[:@12877.4]
  input         io_flow, // @[:@12878.4]
  input  [31:0] io_in, // @[:@12878.4]
  output [31:0] io_out // @[:@12878.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12880.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12880.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12880.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12880.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12880.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12880.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@12880.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12893.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12892.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12891.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12890.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12889.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12887.4]
endmodule
module RetimeWrapper_154( // @[:@13128.2]
  input   clock, // @[:@13129.4]
  input   reset, // @[:@13130.4]
  input   io_flow, // @[:@13131.4]
  input   io_in, // @[:@13131.4]
  output  io_out // @[:@13131.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@13133.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@13133.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@13133.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13133.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13133.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13133.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@13133.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13146.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13145.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@13144.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13143.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13142.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13140.4]
endmodule
module RetimeWrapper_156( // @[:@13192.2]
  input   clock, // @[:@13193.4]
  input   reset, // @[:@13194.4]
  input   io_flow, // @[:@13195.4]
  input   io_in, // @[:@13195.4]
  output  io_out // @[:@13195.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@13197.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@13197.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@13197.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13197.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13197.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13197.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@13197.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13210.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13209.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@13208.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13207.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13206.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13204.4]
endmodule
module RetimeWrapper_158( // @[:@13256.2]
  input         clock, // @[:@13257.4]
  input         reset, // @[:@13258.4]
  input         io_flow, // @[:@13259.4]
  input  [31:0] io_in, // @[:@13259.4]
  output [31:0] io_out // @[:@13259.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13261.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13261.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13261.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13261.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13261.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13261.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(22)) sr ( // @[RetimeShiftRegister.scala 15:20:@13261.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13274.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13273.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@13272.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13271.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13270.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13268.4]
endmodule
module RetimeWrapper_161( // @[:@13352.2]
  input         clock, // @[:@13353.4]
  input         reset, // @[:@13354.4]
  input         io_flow, // @[:@13355.4]
  input  [31:0] io_in, // @[:@13355.4]
  output [31:0] io_out // @[:@13355.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13357.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13357.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13357.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13357.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13357.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13357.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@13357.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13370.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13369.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@13368.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13367.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13366.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13364.4]
endmodule
module RetimeWrapper_164( // @[:@13605.2]
  input   clock, // @[:@13606.4]
  input   reset, // @[:@13607.4]
  input   io_flow, // @[:@13608.4]
  input   io_in, // @[:@13608.4]
  output  io_out // @[:@13608.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@13610.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@13610.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@13610.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13610.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13610.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13610.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@13610.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13623.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13622.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@13621.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13620.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13619.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13617.4]
endmodule
module RetimeWrapper_165( // @[:@13637.2]
  input         clock, // @[:@13638.4]
  input         reset, // @[:@13639.4]
  input         io_flow, // @[:@13640.4]
  input  [31:0] io_in, // @[:@13640.4]
  output [31:0] io_out // @[:@13640.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13642.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13642.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13642.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13642.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13642.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13642.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@13642.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13655.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13654.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@13653.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13652.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13651.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13649.4]
endmodule
module RetimeWrapper_168( // @[:@13890.2]
  input         clock, // @[:@13891.4]
  input         reset, // @[:@13892.4]
  input         io_flow, // @[:@13893.4]
  input  [31:0] io_in, // @[:@13893.4]
  output [31:0] io_out // @[:@13893.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13895.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13895.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13895.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13895.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13895.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13895.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(15)) sr ( // @[RetimeShiftRegister.scala 15:20:@13895.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13908.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13907.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@13906.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13905.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13904.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13902.4]
endmodule
module RetimeWrapper_170( // @[:@14111.2]
  input         clock, // @[:@14112.4]
  input         reset, // @[:@14113.4]
  input         io_flow, // @[:@14114.4]
  input  [31:0] io_in, // @[:@14114.4]
  output [31:0] io_out // @[:@14114.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14116.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14116.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14116.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14116.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14116.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14116.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@14116.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14129.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14128.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14127.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14126.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14125.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14123.4]
endmodule
module x316_rdrow( // @[:@14908.2]
  input         clock, // @[:@14909.4]
  input         reset, // @[:@14910.4]
  input  [31:0] io_a, // @[:@14911.4]
  input  [31:0] io_b, // @[:@14911.4]
  input         io_flow, // @[:@14911.4]
  output [31:0] io_result // @[:@14911.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@14919.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@14919.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@14926.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@14926.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@14945.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@14945.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@14945.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@14945.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@14945.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@14924.4 Math.scala 713:14:@14925.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@14931.4 Math.scala 713:14:@14932.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@14933.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@14934.4]
  __2 _ ( // @[Math.scala 709:24:@14919.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@14926.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@14945.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@14924.4 Math.scala 713:14:@14925.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@14931.4 Math.scala 713:14:@14932.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@14933.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@14934.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@14953.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@14922.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@14929.4]
  assign fix2fixBox_clock = clock; // @[:@14946.4]
  assign fix2fixBox_reset = reset; // @[:@14947.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@14948.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@14951.4]
endmodule
module SimBlackBoxesfix2fixBox_40( // @[:@17617.2]
  input  [7:0] io_a, // @[:@17620.4]
  output [8:0] io_b // @[:@17620.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@17634.4]
endmodule
module __40( // @[:@17636.2]
  input  [7:0] io_b, // @[:@17639.4]
  output [8:0] io_result // @[:@17639.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@17644.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@17644.4]
  SimBlackBoxesfix2fixBox_40 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@17644.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@17657.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@17652.4]
endmodule
module fix2fixBox_22( // @[:@17733.2]
  input        clock, // @[:@17734.4]
  input        reset, // @[:@17735.4]
  input  [8:0] io_a, // @[:@17736.4]
  input        io_flow, // @[:@17736.4]
  output [7:0] io_b // @[:@17736.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17749.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17749.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17749.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@17749.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@17749.4]
  RetimeWrapper_136 RetimeWrapper ( // @[package.scala 93:22:@17749.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@17756.4]
  assign RetimeWrapper_clock = clock; // @[:@17750.4]
  assign RetimeWrapper_reset = reset; // @[:@17751.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@17753.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@17752.4]
endmodule
module x373_x11( // @[:@17758.2]
  input        clock, // @[:@17759.4]
  input        reset, // @[:@17760.4]
  input  [7:0] io_a, // @[:@17761.4]
  input  [7:0] io_b, // @[:@17761.4]
  input        io_flow, // @[:@17761.4]
  output [7:0] io_result // @[:@17761.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@17769.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@17769.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@17776.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@17776.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@17786.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@17786.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@17786.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@17786.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@17786.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@17774.4 Math.scala 713:14:@17775.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@17781.4 Math.scala 713:14:@17782.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@17783.4]
  __40 _ ( // @[Math.scala 709:24:@17769.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __40 __1 ( // @[Math.scala 709:24:@17776.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_22 fix2fixBox ( // @[Math.scala 141:30:@17786.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@17774.4 Math.scala 713:14:@17775.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@17781.4 Math.scala 713:14:@17782.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@17783.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@17794.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@17772.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@17779.4]
  assign fix2fixBox_clock = clock; // @[:@17787.4]
  assign fix2fixBox_reset = reset; // @[:@17788.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@17789.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@17792.4]
endmodule
module RetimeWrapper_224( // @[:@18409.2]
  input        clock, // @[:@18410.4]
  input        reset, // @[:@18411.4]
  input        io_flow, // @[:@18412.4]
  input  [7:0] io_in, // @[:@18412.4]
  output [7:0] io_out // @[:@18412.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18414.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18414.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18414.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18414.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18414.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18414.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@18414.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18427.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18426.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18425.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18424.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18423.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18421.4]
endmodule
module fix2fixBox_26( // @[:@18545.2]
  input  [8:0] io_a, // @[:@18548.4]
  output [7:0] io_b // @[:@18548.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@18561.4]
endmodule
module x377_x11( // @[:@18563.2]
  input  [7:0] io_a, // @[:@18566.4]
  input  [7:0] io_b, // @[:@18566.4]
  output [7:0] io_result // @[:@18566.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@18574.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@18574.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@18581.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@18581.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@18591.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@18591.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@18579.4 Math.scala 713:14:@18580.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@18586.4 Math.scala 713:14:@18587.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@18588.4]
  __40 _ ( // @[Math.scala 709:24:@18574.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __40 __1 ( // @[Math.scala 709:24:@18581.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_26 fix2fixBox ( // @[Math.scala 141:30:@18591.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@18579.4 Math.scala 713:14:@18580.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@18586.4 Math.scala 713:14:@18587.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@18588.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@18599.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@18577.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@18584.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@18594.4]
endmodule
module RetimeWrapper_226( // @[:@18753.2]
  input        clock, // @[:@18754.4]
  input        reset, // @[:@18755.4]
  input        io_flow, // @[:@18756.4]
  input  [7:0] io_in, // @[:@18756.4]
  output [7:0] io_out // @[:@18756.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18758.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18758.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18758.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18758.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18758.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18758.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@18758.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18771.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18770.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18769.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18768.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18767.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18765.4]
endmodule
module RetimeWrapper_227( // @[:@18925.2]
  input        clock, // @[:@18926.4]
  input        reset, // @[:@18927.4]
  input        io_flow, // @[:@18928.4]
  input  [7:0] io_in, // @[:@18928.4]
  output [7:0] io_out // @[:@18928.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18930.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18930.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18930.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18930.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18930.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18930.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@18930.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18943.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18942.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18941.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18940.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18939.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18937.4]
endmodule
module RetimeWrapper_244( // @[:@20757.2]
  input         clock, // @[:@20758.4]
  input         reset, // @[:@20759.4]
  input         io_flow, // @[:@20760.4]
  input  [15:0] io_in, // @[:@20760.4]
  output [15:0] io_out // @[:@20760.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20762.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20762.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20762.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20762.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20762.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20762.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@20762.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20775.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20774.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@20773.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20772.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20771.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20769.4]
endmodule
module x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@20873.2]
  input          clock, // @[:@20874.4]
  input          reset, // @[:@20875.4]
  output         io_in_x244_TREADY, // @[:@20876.4]
  input  [255:0] io_in_x244_TDATA, // @[:@20876.4]
  input  [7:0]   io_in_x244_TID, // @[:@20876.4]
  input  [7:0]   io_in_x244_TDEST, // @[:@20876.4]
  output         io_in_x245_TVALID, // @[:@20876.4]
  input          io_in_x245_TREADY, // @[:@20876.4]
  output [255:0] io_in_x245_TDATA, // @[:@20876.4]
  input          io_sigsIn_backpressure, // @[:@20876.4]
  input          io_sigsIn_datapathEn, // @[:@20876.4]
  input          io_sigsIn_break, // @[:@20876.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@20876.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@20876.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@20876.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@20876.4]
  input          io_rr // @[:@20876.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@20890.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@20890.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@20902.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@20902.4]
  wire  x257_lb_0_clock; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_reset; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_11_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_11_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_11_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_11_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_11_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_11_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_10_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_10_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_10_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_10_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_10_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_10_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_9_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_9_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_9_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_9_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_9_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_9_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_8_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_8_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_8_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_8_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_8_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_8_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_7_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_7_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_7_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_7_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_7_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_7_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_6_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_6_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_6_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_6_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_6_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_6_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_5_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_5_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_5_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_5_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_5_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_5_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_4_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_4_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_4_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_4_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_4_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_4_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_3_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_3_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_3_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_3_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_3_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_3_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_2_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_2_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_2_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_2_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_2_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_2_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_1_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_1_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_1_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_1_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_1_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_1_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_0_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_rPort_0_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_rPort_0_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_0_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_rPort_0_backpressure; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_rPort_0_output_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_wPort_1_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_wPort_1_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_wPort_1_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_wPort_1_data_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_wPort_1_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_wPort_0_banks_1; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [2:0] x257_lb_0_io_wPort_0_banks_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [8:0] x257_lb_0_io_wPort_0_ofs_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire [7:0] x257_lb_0_io_wPort_0_data_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  x257_lb_0_io_wPort_0_en_0; // @[m_x257_lb_0.scala 39:17:@20912.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@21018.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@21018.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@21018.4]
  wire [15:0] RetimeWrapper_io_in; // @[package.scala 93:22:@21018.4]
  wire [15:0] RetimeWrapper_io_out; // @[package.scala 93:22:@21018.4]
  wire  x272_sum_1_clock; // @[Math.scala 150:24:@21130.4]
  wire  x272_sum_1_reset; // @[Math.scala 150:24:@21130.4]
  wire [31:0] x272_sum_1_io_a; // @[Math.scala 150:24:@21130.4]
  wire [31:0] x272_sum_1_io_b; // @[Math.scala 150:24:@21130.4]
  wire  x272_sum_1_io_flow; // @[Math.scala 150:24:@21130.4]
  wire [31:0] x272_sum_1_io_result; // @[Math.scala 150:24:@21130.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@21140.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@21140.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@21140.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@21140.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@21140.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@21149.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@21149.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@21149.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@21149.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@21149.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@21158.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@21158.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@21158.4]
  wire [7:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@21158.4]
  wire [7:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@21158.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@21167.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@21167.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@21167.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@21167.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@21167.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@21176.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@21176.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@21176.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@21176.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@21176.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@21185.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@21185.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@21185.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@21185.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@21185.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@21196.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@21196.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@21196.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@21196.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@21196.4]
  wire  x274_rdcol_1_clock; // @[Math.scala 150:24:@21219.4]
  wire  x274_rdcol_1_reset; // @[Math.scala 150:24:@21219.4]
  wire [31:0] x274_rdcol_1_io_a; // @[Math.scala 150:24:@21219.4]
  wire [31:0] x274_rdcol_1_io_b; // @[Math.scala 150:24:@21219.4]
  wire  x274_rdcol_1_io_flow; // @[Math.scala 150:24:@21219.4]
  wire [31:0] x274_rdcol_1_io_result; // @[Math.scala 150:24:@21219.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@21251.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@21251.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@21251.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@21251.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@21251.4]
  wire  x278_sum_1_clock; // @[Math.scala 150:24:@21260.4]
  wire  x278_sum_1_reset; // @[Math.scala 150:24:@21260.4]
  wire [31:0] x278_sum_1_io_a; // @[Math.scala 150:24:@21260.4]
  wire [31:0] x278_sum_1_io_b; // @[Math.scala 150:24:@21260.4]
  wire  x278_sum_1_io_flow; // @[Math.scala 150:24:@21260.4]
  wire [31:0] x278_sum_1_io_result; // @[Math.scala 150:24:@21260.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@21270.4]
  wire [7:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@21270.4]
  wire [7:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@21279.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@21279.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@21279.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@21279.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@21279.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@21290.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@21290.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@21290.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@21290.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@21290.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@21311.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@21311.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@21311.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@21311.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@21311.4]
  wire  x281_1_clock; // @[Math.scala 366:24:@21322.4]
  wire  x281_1_reset; // @[Math.scala 366:24:@21322.4]
  wire [31:0] x281_1_io_a; // @[Math.scala 366:24:@21322.4]
  wire  x281_1_io_flow; // @[Math.scala 366:24:@21322.4]
  wire [31:0] x281_1_io_result; // @[Math.scala 366:24:@21322.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@21339.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@21339.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@21339.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@21339.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@21339.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@21355.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@21355.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@21355.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@21355.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@21355.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@21395.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@21395.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@21395.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@21395.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@21395.4]
  wire  x289_sum_1_clock; // @[Math.scala 150:24:@21404.4]
  wire  x289_sum_1_reset; // @[Math.scala 150:24:@21404.4]
  wire [31:0] x289_sum_1_io_a; // @[Math.scala 150:24:@21404.4]
  wire [31:0] x289_sum_1_io_b; // @[Math.scala 150:24:@21404.4]
  wire  x289_sum_1_io_flow; // @[Math.scala 150:24:@21404.4]
  wire [31:0] x289_sum_1_io_result; // @[Math.scala 150:24:@21404.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@21414.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@21414.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@21414.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@21414.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@21414.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@21423.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@21423.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@21423.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@21423.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@21423.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@21432.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@21432.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@21432.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@21432.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@21432.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@21450.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@21450.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@21450.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@21450.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@21450.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@21459.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@21459.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@21459.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@21459.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@21459.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@21471.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@21471.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@21471.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@21471.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@21471.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@21492.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@21492.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@21492.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@21492.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@21492.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@21516.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@21516.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@21516.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@21516.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@21516.4]
  wire  x295_sum_1_clock; // @[Math.scala 150:24:@21525.4]
  wire  x295_sum_1_reset; // @[Math.scala 150:24:@21525.4]
  wire [31:0] x295_sum_1_io_a; // @[Math.scala 150:24:@21525.4]
  wire [31:0] x295_sum_1_io_b; // @[Math.scala 150:24:@21525.4]
  wire  x295_sum_1_io_flow; // @[Math.scala 150:24:@21525.4]
  wire [31:0] x295_sum_1_io_result; // @[Math.scala 150:24:@21525.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@21535.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@21535.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@21535.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@21535.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@21535.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@21544.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@21544.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@21544.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@21544.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@21544.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@21553.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@21553.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@21553.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@21553.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@21553.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@21565.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@21565.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@21565.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@21565.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@21565.4]
  wire  x298_rdcol_1_clock; // @[Math.scala 150:24:@21588.4]
  wire  x298_rdcol_1_reset; // @[Math.scala 150:24:@21588.4]
  wire [31:0] x298_rdcol_1_io_a; // @[Math.scala 150:24:@21588.4]
  wire [31:0] x298_rdcol_1_io_b; // @[Math.scala 150:24:@21588.4]
  wire  x298_rdcol_1_io_flow; // @[Math.scala 150:24:@21588.4]
  wire [31:0] x298_rdcol_1_io_result; // @[Math.scala 150:24:@21588.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@21631.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@21631.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@21631.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@21631.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@21631.4]
  wire  x304_sum_1_clock; // @[Math.scala 150:24:@21640.4]
  wire  x304_sum_1_reset; // @[Math.scala 150:24:@21640.4]
  wire [31:0] x304_sum_1_io_a; // @[Math.scala 150:24:@21640.4]
  wire [31:0] x304_sum_1_io_b; // @[Math.scala 150:24:@21640.4]
  wire  x304_sum_1_io_flow; // @[Math.scala 150:24:@21640.4]
  wire [31:0] x304_sum_1_io_result; // @[Math.scala 150:24:@21640.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@21650.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@21650.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@21650.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@21650.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@21650.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@21659.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@21659.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@21659.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@21659.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@21659.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@21668.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@21668.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@21668.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@21668.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@21668.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@21680.4]
  wire  x307_rdcol_1_clock; // @[Math.scala 150:24:@21703.4]
  wire  x307_rdcol_1_reset; // @[Math.scala 150:24:@21703.4]
  wire [31:0] x307_rdcol_1_io_a; // @[Math.scala 150:24:@21703.4]
  wire [31:0] x307_rdcol_1_io_b; // @[Math.scala 150:24:@21703.4]
  wire  x307_rdcol_1_io_flow; // @[Math.scala 150:24:@21703.4]
  wire [31:0] x307_rdcol_1_io_result; // @[Math.scala 150:24:@21703.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@21746.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@21746.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@21746.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@21746.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@21746.4]
  wire  x313_sum_1_clock; // @[Math.scala 150:24:@21755.4]
  wire  x313_sum_1_reset; // @[Math.scala 150:24:@21755.4]
  wire [31:0] x313_sum_1_io_a; // @[Math.scala 150:24:@21755.4]
  wire [31:0] x313_sum_1_io_b; // @[Math.scala 150:24:@21755.4]
  wire  x313_sum_1_io_flow; // @[Math.scala 150:24:@21755.4]
  wire [31:0] x313_sum_1_io_result; // @[Math.scala 150:24:@21755.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@21765.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@21765.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@21765.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@21765.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@21765.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@21774.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@21774.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@21774.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@21774.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@21774.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@21795.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@21795.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@21795.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@21795.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@21795.4]
  wire  x316_rdrow_1_clock; // @[Math.scala 191:24:@21818.4]
  wire  x316_rdrow_1_reset; // @[Math.scala 191:24:@21818.4]
  wire [31:0] x316_rdrow_1_io_a; // @[Math.scala 191:24:@21818.4]
  wire [31:0] x316_rdrow_1_io_b; // @[Math.scala 191:24:@21818.4]
  wire  x316_rdrow_1_io_flow; // @[Math.scala 191:24:@21818.4]
  wire [31:0] x316_rdrow_1_io_result; // @[Math.scala 191:24:@21818.4]
  wire  x317_1_clock; // @[Math.scala 366:24:@21830.4]
  wire  x317_1_reset; // @[Math.scala 366:24:@21830.4]
  wire [31:0] x317_1_io_a; // @[Math.scala 366:24:@21830.4]
  wire  x317_1_io_flow; // @[Math.scala 366:24:@21830.4]
  wire [31:0] x317_1_io_result; // @[Math.scala 366:24:@21830.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@21880.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@21880.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@21880.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@21880.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@21880.4]
  wire  x324_sum_1_clock; // @[Math.scala 150:24:@21889.4]
  wire  x324_sum_1_reset; // @[Math.scala 150:24:@21889.4]
  wire [31:0] x324_sum_1_io_a; // @[Math.scala 150:24:@21889.4]
  wire [31:0] x324_sum_1_io_b; // @[Math.scala 150:24:@21889.4]
  wire  x324_sum_1_io_flow; // @[Math.scala 150:24:@21889.4]
  wire [31:0] x324_sum_1_io_result; // @[Math.scala 150:24:@21889.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@21899.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@21899.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@21899.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@21899.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@21899.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@21908.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@21908.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@21908.4]
  wire [31:0] RetimeWrapper_41_io_in; // @[package.scala 93:22:@21908.4]
  wire [31:0] RetimeWrapper_41_io_out; // @[package.scala 93:22:@21908.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@21920.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@21920.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@21920.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@21920.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@21920.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@21941.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@21941.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@21941.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@21941.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@21941.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@21956.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@21956.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@21956.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@21956.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@21956.4]
  wire  x329_sum_1_clock; // @[Math.scala 150:24:@21965.4]
  wire  x329_sum_1_reset; // @[Math.scala 150:24:@21965.4]
  wire [31:0] x329_sum_1_io_a; // @[Math.scala 150:24:@21965.4]
  wire [31:0] x329_sum_1_io_b; // @[Math.scala 150:24:@21965.4]
  wire  x329_sum_1_io_flow; // @[Math.scala 150:24:@21965.4]
  wire [31:0] x329_sum_1_io_result; // @[Math.scala 150:24:@21965.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@21975.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@21975.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@21975.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@21975.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@21975.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@21987.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@21987.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@21987.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@21987.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@21987.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@22014.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@22014.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@22014.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@22014.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@22014.4]
  wire  x334_sum_1_clock; // @[Math.scala 150:24:@22023.4]
  wire  x334_sum_1_reset; // @[Math.scala 150:24:@22023.4]
  wire [31:0] x334_sum_1_io_a; // @[Math.scala 150:24:@22023.4]
  wire [31:0] x334_sum_1_io_b; // @[Math.scala 150:24:@22023.4]
  wire  x334_sum_1_io_flow; // @[Math.scala 150:24:@22023.4]
  wire [31:0] x334_sum_1_io_result; // @[Math.scala 150:24:@22023.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@22033.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@22033.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@22033.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@22033.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@22033.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@22045.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@22045.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@22045.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@22045.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@22045.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@22072.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@22072.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@22072.4]
  wire [31:0] RetimeWrapper_50_io_in; // @[package.scala 93:22:@22072.4]
  wire [31:0] RetimeWrapper_50_io_out; // @[package.scala 93:22:@22072.4]
  wire  x339_sum_1_clock; // @[Math.scala 150:24:@22081.4]
  wire  x339_sum_1_reset; // @[Math.scala 150:24:@22081.4]
  wire [31:0] x339_sum_1_io_a; // @[Math.scala 150:24:@22081.4]
  wire [31:0] x339_sum_1_io_b; // @[Math.scala 150:24:@22081.4]
  wire  x339_sum_1_io_flow; // @[Math.scala 150:24:@22081.4]
  wire [31:0] x339_sum_1_io_result; // @[Math.scala 150:24:@22081.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@22091.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@22091.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@22091.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@22091.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@22091.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@22103.4]
  wire  x342_rdrow_1_clock; // @[Math.scala 191:24:@22126.4]
  wire  x342_rdrow_1_reset; // @[Math.scala 191:24:@22126.4]
  wire [31:0] x342_rdrow_1_io_a; // @[Math.scala 191:24:@22126.4]
  wire [31:0] x342_rdrow_1_io_b; // @[Math.scala 191:24:@22126.4]
  wire  x342_rdrow_1_io_flow; // @[Math.scala 191:24:@22126.4]
  wire [31:0] x342_rdrow_1_io_result; // @[Math.scala 191:24:@22126.4]
  wire  x343_1_clock; // @[Math.scala 366:24:@22138.4]
  wire  x343_1_reset; // @[Math.scala 366:24:@22138.4]
  wire [31:0] x343_1_io_a; // @[Math.scala 366:24:@22138.4]
  wire  x343_1_io_flow; // @[Math.scala 366:24:@22138.4]
  wire [31:0] x343_1_io_result; // @[Math.scala 366:24:@22138.4]
  wire  x350_sum_1_clock; // @[Math.scala 150:24:@22186.4]
  wire  x350_sum_1_reset; // @[Math.scala 150:24:@22186.4]
  wire [31:0] x350_sum_1_io_a; // @[Math.scala 150:24:@22186.4]
  wire [31:0] x350_sum_1_io_b; // @[Math.scala 150:24:@22186.4]
  wire  x350_sum_1_io_flow; // @[Math.scala 150:24:@22186.4]
  wire [31:0] x350_sum_1_io_result; // @[Math.scala 150:24:@22186.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@22196.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@22196.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@22196.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@22196.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@22196.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@22205.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@22205.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@22205.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@22205.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@22205.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@22217.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@22217.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@22217.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@22217.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@22217.4]
  wire  x355_sum_1_clock; // @[Math.scala 150:24:@22244.4]
  wire  x355_sum_1_reset; // @[Math.scala 150:24:@22244.4]
  wire [31:0] x355_sum_1_io_a; // @[Math.scala 150:24:@22244.4]
  wire [31:0] x355_sum_1_io_b; // @[Math.scala 150:24:@22244.4]
  wire  x355_sum_1_io_flow; // @[Math.scala 150:24:@22244.4]
  wire [31:0] x355_sum_1_io_result; // @[Math.scala 150:24:@22244.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@22254.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@22254.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@22254.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@22254.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@22254.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@22266.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@22266.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@22266.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@22266.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@22266.4]
  wire  x360_sum_1_clock; // @[Math.scala 150:24:@22295.4]
  wire  x360_sum_1_reset; // @[Math.scala 150:24:@22295.4]
  wire [31:0] x360_sum_1_io_a; // @[Math.scala 150:24:@22295.4]
  wire [31:0] x360_sum_1_io_b; // @[Math.scala 150:24:@22295.4]
  wire  x360_sum_1_io_flow; // @[Math.scala 150:24:@22295.4]
  wire [31:0] x360_sum_1_io_result; // @[Math.scala 150:24:@22295.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@22305.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@22305.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@22305.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@22305.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@22305.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@22317.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@22317.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@22317.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@22317.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@22317.4]
  wire  x365_sum_1_clock; // @[Math.scala 150:24:@22344.4]
  wire  x365_sum_1_reset; // @[Math.scala 150:24:@22344.4]
  wire [31:0] x365_sum_1_io_a; // @[Math.scala 150:24:@22344.4]
  wire [31:0] x365_sum_1_io_b; // @[Math.scala 150:24:@22344.4]
  wire  x365_sum_1_io_flow; // @[Math.scala 150:24:@22344.4]
  wire [31:0] x365_sum_1_io_result; // @[Math.scala 150:24:@22344.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@22354.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@22354.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@22354.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@22354.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@22354.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@22366.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@22366.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@22366.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@22366.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@22366.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@22412.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@22412.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@22412.4]
  wire [7:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@22412.4]
  wire [7:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@22412.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@22421.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@22421.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@22421.4]
  wire [7:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@22421.4]
  wire [7:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@22421.4]
  wire  x373_x11_1_clock; // @[Math.scala 150:24:@22430.4]
  wire  x373_x11_1_reset; // @[Math.scala 150:24:@22430.4]
  wire [7:0] x373_x11_1_io_a; // @[Math.scala 150:24:@22430.4]
  wire [7:0] x373_x11_1_io_b; // @[Math.scala 150:24:@22430.4]
  wire  x373_x11_1_io_flow; // @[Math.scala 150:24:@22430.4]
  wire [7:0] x373_x11_1_io_result; // @[Math.scala 150:24:@22430.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@22440.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@22440.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@22440.4]
  wire [7:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@22440.4]
  wire [7:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@22440.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@22449.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@22449.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@22449.4]
  wire [7:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@22449.4]
  wire [7:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@22449.4]
  wire  x374_x12_1_clock; // @[Math.scala 150:24:@22458.4]
  wire  x374_x12_1_reset; // @[Math.scala 150:24:@22458.4]
  wire [7:0] x374_x12_1_io_a; // @[Math.scala 150:24:@22458.4]
  wire [7:0] x374_x12_1_io_b; // @[Math.scala 150:24:@22458.4]
  wire  x374_x12_1_io_flow; // @[Math.scala 150:24:@22458.4]
  wire [7:0] x374_x12_1_io_result; // @[Math.scala 150:24:@22458.4]
  wire  x375_x11_1_clock; // @[Math.scala 150:24:@22468.4]
  wire  x375_x11_1_reset; // @[Math.scala 150:24:@22468.4]
  wire [7:0] x375_x11_1_io_a; // @[Math.scala 150:24:@22468.4]
  wire [7:0] x375_x11_1_io_b; // @[Math.scala 150:24:@22468.4]
  wire  x375_x11_1_io_flow; // @[Math.scala 150:24:@22468.4]
  wire [7:0] x375_x11_1_io_result; // @[Math.scala 150:24:@22468.4]
  wire  x376_x12_1_clock; // @[Math.scala 150:24:@22478.4]
  wire  x376_x12_1_reset; // @[Math.scala 150:24:@22478.4]
  wire [7:0] x376_x12_1_io_a; // @[Math.scala 150:24:@22478.4]
  wire [7:0] x376_x12_1_io_b; // @[Math.scala 150:24:@22478.4]
  wire  x376_x12_1_io_flow; // @[Math.scala 150:24:@22478.4]
  wire [7:0] x376_x12_1_io_result; // @[Math.scala 150:24:@22478.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@22488.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@22488.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@22488.4]
  wire [7:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@22488.4]
  wire [7:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@22488.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@22497.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@22497.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@22497.4]
  wire [7:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@22497.4]
  wire [7:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@22497.4]
  wire [7:0] x377_x11_1_io_a; // @[Math.scala 150:24:@22506.4]
  wire [7:0] x377_x11_1_io_b; // @[Math.scala 150:24:@22506.4]
  wire [7:0] x377_x11_1_io_result; // @[Math.scala 150:24:@22506.4]
  wire [7:0] x378_x12_1_io_a; // @[Math.scala 150:24:@22516.4]
  wire [7:0] x378_x12_1_io_b; // @[Math.scala 150:24:@22516.4]
  wire [7:0] x378_x12_1_io_result; // @[Math.scala 150:24:@22516.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@22526.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@22526.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@22526.4]
  wire [7:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@22526.4]
  wire [7:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@22526.4]
  wire [7:0] x379_x11_1_io_a; // @[Math.scala 150:24:@22535.4]
  wire [7:0] x379_x11_1_io_b; // @[Math.scala 150:24:@22535.4]
  wire [7:0] x379_x11_1_io_result; // @[Math.scala 150:24:@22535.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@22545.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@22545.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@22545.4]
  wire [7:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@22545.4]
  wire [7:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@22545.4]
  wire [7:0] x380_sum_1_io_a; // @[Math.scala 150:24:@22554.4]
  wire [7:0] x380_sum_1_io_b; // @[Math.scala 150:24:@22554.4]
  wire [7:0] x380_sum_1_io_result; // @[Math.scala 150:24:@22554.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@22568.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@22568.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@22568.4]
  wire [7:0] RetimeWrapper_70_io_in; // @[package.scala 93:22:@22568.4]
  wire [7:0] RetimeWrapper_70_io_out; // @[package.scala 93:22:@22568.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@22603.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@22603.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@22603.4]
  wire [7:0] RetimeWrapper_71_io_in; // @[package.scala 93:22:@22603.4]
  wire [7:0] RetimeWrapper_71_io_out; // @[package.scala 93:22:@22603.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@22612.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@22612.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@22612.4]
  wire [7:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@22612.4]
  wire [7:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@22612.4]
  wire  x387_x11_1_clock; // @[Math.scala 150:24:@22621.4]
  wire  x387_x11_1_reset; // @[Math.scala 150:24:@22621.4]
  wire [7:0] x387_x11_1_io_a; // @[Math.scala 150:24:@22621.4]
  wire [7:0] x387_x11_1_io_b; // @[Math.scala 150:24:@22621.4]
  wire  x387_x11_1_io_flow; // @[Math.scala 150:24:@22621.4]
  wire [7:0] x387_x11_1_io_result; // @[Math.scala 150:24:@22621.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@22631.4]
  wire [7:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@22631.4]
  wire [7:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@22640.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@22640.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@22640.4]
  wire [7:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@22640.4]
  wire [7:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@22640.4]
  wire  x388_x12_1_clock; // @[Math.scala 150:24:@22649.4]
  wire  x388_x12_1_reset; // @[Math.scala 150:24:@22649.4]
  wire [7:0] x388_x12_1_io_a; // @[Math.scala 150:24:@22649.4]
  wire [7:0] x388_x12_1_io_b; // @[Math.scala 150:24:@22649.4]
  wire  x388_x12_1_io_flow; // @[Math.scala 150:24:@22649.4]
  wire [7:0] x388_x12_1_io_result; // @[Math.scala 150:24:@22649.4]
  wire  x389_x11_1_clock; // @[Math.scala 150:24:@22659.4]
  wire  x389_x11_1_reset; // @[Math.scala 150:24:@22659.4]
  wire [7:0] x389_x11_1_io_a; // @[Math.scala 150:24:@22659.4]
  wire [7:0] x389_x11_1_io_b; // @[Math.scala 150:24:@22659.4]
  wire  x389_x11_1_io_flow; // @[Math.scala 150:24:@22659.4]
  wire [7:0] x389_x11_1_io_result; // @[Math.scala 150:24:@22659.4]
  wire  x390_x12_1_clock; // @[Math.scala 150:24:@22669.4]
  wire  x390_x12_1_reset; // @[Math.scala 150:24:@22669.4]
  wire [7:0] x390_x12_1_io_a; // @[Math.scala 150:24:@22669.4]
  wire [7:0] x390_x12_1_io_b; // @[Math.scala 150:24:@22669.4]
  wire  x390_x12_1_io_flow; // @[Math.scala 150:24:@22669.4]
  wire [7:0] x390_x12_1_io_result; // @[Math.scala 150:24:@22669.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@22679.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@22679.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@22679.4]
  wire [7:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@22679.4]
  wire [7:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@22679.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@22688.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@22688.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@22688.4]
  wire [7:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@22688.4]
  wire [7:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@22688.4]
  wire [7:0] x391_x11_1_io_a; // @[Math.scala 150:24:@22699.4]
  wire [7:0] x391_x11_1_io_b; // @[Math.scala 150:24:@22699.4]
  wire [7:0] x391_x11_1_io_result; // @[Math.scala 150:24:@22699.4]
  wire [7:0] x392_x12_1_io_a; // @[Math.scala 150:24:@22709.4]
  wire [7:0] x392_x12_1_io_b; // @[Math.scala 150:24:@22709.4]
  wire [7:0] x392_x12_1_io_result; // @[Math.scala 150:24:@22709.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@22719.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@22719.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@22719.4]
  wire [7:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@22719.4]
  wire [7:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@22719.4]
  wire [7:0] x393_x11_1_io_a; // @[Math.scala 150:24:@22728.4]
  wire [7:0] x393_x11_1_io_b; // @[Math.scala 150:24:@22728.4]
  wire [7:0] x393_x11_1_io_result; // @[Math.scala 150:24:@22728.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@22738.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@22738.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@22738.4]
  wire [7:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@22738.4]
  wire [7:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@22738.4]
  wire [7:0] x394_sum_1_io_a; // @[Math.scala 150:24:@22747.4]
  wire [7:0] x394_sum_1_io_b; // @[Math.scala 150:24:@22747.4]
  wire [7:0] x394_sum_1_io_result; // @[Math.scala 150:24:@22747.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@22761.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@22761.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@22761.4]
  wire [7:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@22761.4]
  wire [7:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@22761.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@22771.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@22771.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@22771.4]
  wire [7:0] RetimeWrapper_80_io_in; // @[package.scala 93:22:@22771.4]
  wire [7:0] RetimeWrapper_80_io_out; // @[package.scala 93:22:@22771.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@22780.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@22780.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@22780.4]
  wire [7:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@22780.4]
  wire [7:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@22780.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@22795.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@22795.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@22795.4]
  wire [15:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@22795.4]
  wire [15:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@22795.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@22804.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@22804.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@22804.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@22804.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@22804.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@22813.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@22813.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@22813.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@22813.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@22813.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@22822.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@22822.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@22822.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@22822.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@22822.4]
  wire  b255; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 62:18:@20910.4]
  wire  b256; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 63:18:@20911.4]
  wire  _T_206; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 68:30:@21006.4]
  wire  _T_207; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 68:37:@21007.4]
  wire  _T_211; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 70:76:@21012.4]
  wire  _T_212; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 70:62:@21013.4]
  wire  _T_214; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 70:101:@21014.4]
  wire [15:0] x476_x258_D1_0_number; // @[package.scala 96:25:@21023.4 package.scala 96:25:@21024.4]
  wire [31:0] b253_number; // @[Math.scala 712:22:@20895.4 Math.scala 713:14:@20896.4]
  wire [31:0] _T_242; // @[Math.scala 499:52:@21039.4]
  wire  x262; // @[Math.scala 499:44:@21047.4]
  wire  x263; // @[Math.scala 499:44:@21054.4]
  wire  x264; // @[Math.scala 499:44:@21061.4]
  wire [31:0] _T_289; // @[Mux.scala 19:72:@21073.4]
  wire [31:0] _T_291; // @[Mux.scala 19:72:@21074.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@21075.4]
  wire [31:0] _T_295; // @[Mux.scala 19:72:@21077.4]
  wire [31:0] x265_number; // @[Mux.scala 19:72:@21078.4]
  wire [31:0] _T_307; // @[Math.scala 406:49:@21088.4]
  wire [31:0] _T_309; // @[Math.scala 406:56:@21090.4]
  wire [31:0] _T_310; // @[Math.scala 406:56:@21091.4]
  wire [31:0] b254_number; // @[Math.scala 712:22:@20907.4 Math.scala 713:14:@20908.4]
  wire [31:0] _T_319; // @[Math.scala 406:49:@21099.4]
  wire [31:0] _T_321; // @[Math.scala 406:56:@21101.4]
  wire [31:0] _T_322; // @[Math.scala 406:56:@21102.4]
  wire  _T_327; // @[FixedPoint.scala 50:25:@21108.4]
  wire [1:0] _T_331; // @[Bitwise.scala 72:12:@21110.4]
  wire [29:0] _T_332; // @[FixedPoint.scala 18:52:@21111.4]
  wire [31:0] x269_number; // @[Cat.scala 30:58:@21112.4]
  wire [39:0] _GEN_0; // @[Math.scala 450:32:@21117.4]
  wire [39:0] _T_337; // @[Math.scala 450:32:@21117.4]
  wire  _T_341; // @[FixedPoint.scala 50:25:@21122.4]
  wire [1:0] _T_345; // @[Bitwise.scala 72:12:@21124.4]
  wire [29:0] _T_346; // @[FixedPoint.scala 18:52:@21125.4]
  wire  _T_370; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:101:@21193.4]
  wire  _T_374; // @[package.scala 96:25:@21201.4 package.scala 96:25:@21202.4]
  wire  _T_376; // @[implicits.scala 55:10:@21203.4]
  wire  _T_377; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:118:@21204.4]
  wire  _T_379; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:206:@21206.4]
  wire  _T_380; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:225:@21207.4]
  wire  x480_b255_D2; // @[package.scala 96:25:@21172.4 package.scala 96:25:@21173.4]
  wire  _T_381; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:251:@21208.4]
  wire  x478_b256_D2; // @[package.scala 96:25:@21154.4 package.scala 96:25:@21155.4]
  wire [31:0] x274_rdcol_number; // @[Math.scala 154:22:@21225.4 Math.scala 155:14:@21226.4]
  wire [31:0] _T_398; // @[Math.scala 406:49:@21234.4]
  wire [31:0] _T_400; // @[Math.scala 406:56:@21236.4]
  wire [31:0] _T_401; // @[Math.scala 406:56:@21237.4]
  wire  _T_406; // @[FixedPoint.scala 50:25:@21243.4]
  wire [1:0] _T_410; // @[Bitwise.scala 72:12:@21245.4]
  wire [29:0] _T_411; // @[FixedPoint.scala 18:52:@21246.4]
  wire  _T_430; // @[package.scala 96:25:@21295.4 package.scala 96:25:@21296.4]
  wire  _T_432; // @[implicits.scala 55:10:@21297.4]
  wire  _T_433; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:118:@21298.4]
  wire  _T_435; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:206:@21300.4]
  wire  _T_436; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:225:@21301.4]
  wire  _T_437; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:251:@21302.4]
  wire [31:0] x486_b253_D5_number; // @[package.scala 96:25:@21316.4 package.scala 96:25:@21317.4]
  wire [31:0] _T_454; // @[Math.scala 465:37:@21334.4]
  wire  x282; // @[Math.scala 465:44:@21336.4]
  wire [31:0] x487_x274_rdcol_D5_number; // @[package.scala 96:25:@21344.4 package.scala 96:25:@21345.4]
  wire [31:0] _T_465; // @[Math.scala 465:37:@21350.4]
  wire  x283; // @[Math.scala 465:44:@21352.4]
  wire  x488_x282_D1; // @[package.scala 96:25:@21360.4 package.scala 96:25:@21361.4]
  wire  x284; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 155:24:@21364.4]
  wire [31:0] x281_number; // @[Math.scala 370:22:@21328.4 Math.scala 371:14:@21329.4]
  wire [31:0] _T_482; // @[Math.scala 406:49:@21373.4]
  wire [31:0] _T_484; // @[Math.scala 406:56:@21375.4]
  wire [31:0] _T_485; // @[Math.scala 406:56:@21376.4]
  wire  _T_490; // @[FixedPoint.scala 50:25:@21382.4]
  wire [1:0] _T_494; // @[Bitwise.scala 72:12:@21384.4]
  wire [29:0] _T_495; // @[FixedPoint.scala 18:52:@21385.4]
  wire [31:0] x287_number; // @[Cat.scala 30:58:@21386.4]
  wire [39:0] _GEN_1; // @[Math.scala 450:32:@21391.4]
  wire [39:0] _T_500; // @[Math.scala 450:32:@21391.4]
  wire  _T_536; // @[package.scala 96:25:@21476.4 package.scala 96:25:@21477.4]
  wire  _T_538; // @[implicits.scala 55:10:@21478.4]
  wire  _T_539; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 190:194:@21479.4]
  wire  x491_x285_D17; // @[package.scala 96:25:@21428.4 package.scala 96:25:@21429.4]
  wire  _T_540; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 190:283:@21480.4]
  wire  x494_b255_D23; // @[package.scala 96:25:@21455.4 package.scala 96:25:@21456.4]
  wire  _T_541; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 190:326:@21481.4]
  wire  x493_b256_D23; // @[package.scala 96:25:@21446.4 package.scala 96:25:@21447.4]
  wire [31:0] x496_b254_D5_number; // @[package.scala 96:25:@21497.4 package.scala 96:25:@21498.4]
  wire [31:0] _T_554; // @[Math.scala 465:37:@21505.4]
  wire  x292; // @[Math.scala 465:44:@21507.4]
  wire  x293; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 200:59:@21510.4]
  wire  _T_587; // @[package.scala 96:25:@21570.4 package.scala 96:25:@21571.4]
  wire  _T_589; // @[implicits.scala 55:10:@21572.4]
  wire  _T_590; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:194:@21573.4]
  wire  x499_x294_D18; // @[package.scala 96:25:@21549.4 package.scala 96:25:@21550.4]
  wire  _T_591; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:283:@21574.4]
  wire  _T_592; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:291:@21575.4]
  wire [31:0] x298_rdcol_number; // @[Math.scala 154:22:@21594.4 Math.scala 155:14:@21595.4]
  wire [31:0] _T_607; // @[Math.scala 465:37:@21600.4]
  wire  x299; // @[Math.scala 465:44:@21602.4]
  wire  x300; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 225:59:@21605.4]
  wire [31:0] _T_623; // @[Math.scala 406:56:@21616.4]
  wire [31:0] _T_624; // @[Math.scala 406:56:@21617.4]
  wire  _T_629; // @[FixedPoint.scala 50:25:@21623.4]
  wire [1:0] _T_633; // @[Bitwise.scala 72:12:@21625.4]
  wire [29:0] _T_634; // @[FixedPoint.scala 18:52:@21626.4]
  wire  _T_662; // @[package.scala 96:25:@21685.4 package.scala 96:25:@21686.4]
  wire  _T_664; // @[implicits.scala 55:10:@21687.4]
  wire  _T_665; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:194:@21688.4]
  wire  x503_x301_D17; // @[package.scala 96:25:@21664.4 package.scala 96:25:@21665.4]
  wire  _T_666; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:283:@21689.4]
  wire  _T_667; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:291:@21690.4]
  wire [31:0] x307_rdcol_number; // @[Math.scala 154:22:@21709.4 Math.scala 155:14:@21710.4]
  wire [31:0] _T_682; // @[Math.scala 465:37:@21715.4]
  wire  x308; // @[Math.scala 465:44:@21717.4]
  wire  x309; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 254:59:@21720.4]
  wire [31:0] _T_698; // @[Math.scala 406:56:@21731.4]
  wire [31:0] _T_699; // @[Math.scala 406:56:@21732.4]
  wire  _T_704; // @[FixedPoint.scala 50:25:@21738.4]
  wire [1:0] _T_708; // @[Bitwise.scala 72:12:@21740.4]
  wire [29:0] _T_709; // @[FixedPoint.scala 18:52:@21741.4]
  wire  _T_737; // @[package.scala 96:25:@21800.4 package.scala 96:25:@21801.4]
  wire  _T_739; // @[implicits.scala 55:10:@21802.4]
  wire  _T_740; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 275:194:@21803.4]
  wire  x508_x310_D17; // @[package.scala 96:25:@21788.4 package.scala 96:25:@21789.4]
  wire  _T_741; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 275:283:@21804.4]
  wire  _T_742; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 275:291:@21805.4]
  wire [31:0] x316_rdrow_number; // @[Math.scala 195:22:@21824.4 Math.scala 196:14:@21825.4]
  wire [31:0] _T_764; // @[Math.scala 465:37:@21842.4]
  wire  x318; // @[Math.scala 465:44:@21844.4]
  wire  x319; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 285:24:@21847.4]
  wire [31:0] x317_number; // @[Math.scala 370:22:@21836.4 Math.scala 371:14:@21837.4]
  wire [31:0] _T_778; // @[Math.scala 406:49:@21856.4]
  wire [31:0] _T_780; // @[Math.scala 406:56:@21858.4]
  wire [31:0] _T_781; // @[Math.scala 406:56:@21859.4]
  wire  _T_788; // @[FixedPoint.scala 50:25:@21867.4]
  wire [1:0] _T_792; // @[Bitwise.scala 72:12:@21869.4]
  wire [29:0] _T_793; // @[FixedPoint.scala 18:52:@21870.4]
  wire [31:0] x322_number; // @[Cat.scala 30:58:@21871.4]
  wire [39:0] _GEN_2; // @[Math.scala 450:32:@21876.4]
  wire [39:0] _T_798; // @[Math.scala 450:32:@21876.4]
  wire  _T_822; // @[package.scala 96:25:@21925.4 package.scala 96:25:@21926.4]
  wire  _T_824; // @[implicits.scala 55:10:@21927.4]
  wire  _T_825; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:194:@21928.4]
  wire  x510_x320_D17; // @[package.scala 96:25:@21904.4 package.scala 96:25:@21905.4]
  wire  _T_826; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:283:@21929.4]
  wire  _T_827; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:291:@21930.4]
  wire  x512_x292_D1; // @[package.scala 96:25:@21946.4 package.scala 96:25:@21947.4]
  wire  x327; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 320:59:@21950.4]
  wire  _T_857; // @[package.scala 96:25:@21992.4 package.scala 96:25:@21993.4]
  wire  _T_859; // @[implicits.scala 55:10:@21994.4]
  wire  _T_860; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:194:@21995.4]
  wire  x514_x328_D17; // @[package.scala 96:25:@21980.4 package.scala 96:25:@21981.4]
  wire  _T_861; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:283:@21996.4]
  wire  _T_862; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:291:@21997.4]
  wire  x332; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 337:59:@22008.4]
  wire  _T_889; // @[package.scala 96:25:@22050.4 package.scala 96:25:@22051.4]
  wire  _T_891; // @[implicits.scala 55:10:@22052.4]
  wire  _T_892; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:194:@22053.4]
  wire  x516_x333_D17; // @[package.scala 96:25:@22038.4 package.scala 96:25:@22039.4]
  wire  _T_893; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:283:@22054.4]
  wire  _T_894; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:291:@22055.4]
  wire  x337; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 354:59:@22066.4]
  wire  _T_921; // @[package.scala 96:25:@22108.4 package.scala 96:25:@22109.4]
  wire  _T_923; // @[implicits.scala 55:10:@22110.4]
  wire  _T_924; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:194:@22111.4]
  wire  x518_x338_D17; // @[package.scala 96:25:@22096.4 package.scala 96:25:@22097.4]
  wire  _T_925; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:283:@22112.4]
  wire  _T_926; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:291:@22113.4]
  wire [31:0] x342_rdrow_number; // @[Math.scala 195:22:@22132.4 Math.scala 196:14:@22133.4]
  wire [31:0] _T_948; // @[Math.scala 465:37:@22150.4]
  wire  x344; // @[Math.scala 465:44:@22152.4]
  wire  x345; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 377:24:@22155.4]
  wire [31:0] x343_number; // @[Math.scala 370:22:@22144.4 Math.scala 371:14:@22145.4]
  wire [31:0] _T_962; // @[Math.scala 406:49:@22164.4]
  wire [31:0] _T_964; // @[Math.scala 406:56:@22166.4]
  wire [31:0] _T_965; // @[Math.scala 406:56:@22167.4]
  wire  _T_970; // @[FixedPoint.scala 50:25:@22173.4]
  wire [1:0] _T_974; // @[Bitwise.scala 72:12:@22175.4]
  wire [29:0] _T_975; // @[FixedPoint.scala 18:52:@22176.4]
  wire [31:0] x348_number; // @[Cat.scala 30:58:@22177.4]
  wire [39:0] _GEN_3; // @[Math.scala 450:32:@22182.4]
  wire [39:0] _T_980; // @[Math.scala 450:32:@22182.4]
  wire  _T_1001; // @[package.scala 96:25:@22222.4 package.scala 96:25:@22223.4]
  wire  _T_1003; // @[implicits.scala 55:10:@22224.4]
  wire  _T_1004; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 396:194:@22225.4]
  wire  x520_x346_D17; // @[package.scala 96:25:@22210.4 package.scala 96:25:@22211.4]
  wire  _T_1005; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 396:283:@22226.4]
  wire  _T_1006; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 396:291:@22227.4]
  wire  x353; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 400:24:@22238.4]
  wire  _T_1030; // @[package.scala 96:25:@22271.4 package.scala 96:25:@22272.4]
  wire  _T_1032; // @[implicits.scala 55:10:@22273.4]
  wire  _T_1033; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:194:@22274.4]
  wire  x521_x354_D17; // @[package.scala 96:25:@22259.4 package.scala 96:25:@22260.4]
  wire  _T_1034; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:283:@22275.4]
  wire  _T_1035; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:291:@22276.4]
  wire  x358; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 421:59:@22287.4]
  wire  _T_1061; // @[package.scala 96:25:@22322.4 package.scala 96:25:@22323.4]
  wire  _T_1063; // @[implicits.scala 55:10:@22324.4]
  wire  _T_1064; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:194:@22325.4]
  wire  x522_x359_D17; // @[package.scala 96:25:@22310.4 package.scala 96:25:@22311.4]
  wire  _T_1065; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:283:@22326.4]
  wire  _T_1066; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:291:@22327.4]
  wire  x363; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 438:59:@22338.4]
  wire  _T_1090; // @[package.scala 96:25:@22371.4 package.scala 96:25:@22372.4]
  wire  _T_1092; // @[implicits.scala 55:10:@22373.4]
  wire  _T_1093; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 449:194:@22374.4]
  wire  x523_x364_D17; // @[package.scala 96:25:@22359.4 package.scala 96:25:@22360.4]
  wire  _T_1094; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 449:283:@22375.4]
  wire  _T_1095; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 449:291:@22376.4]
  wire [7:0] x296_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 213:29:@21561.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:338:@21582.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@22388.4]
  wire [8:0] _T_1101; // @[Math.scala 450:32:@22388.4]
  wire [7:0] x325_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 310:29:@21916.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:408:@21937.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@22393.4]
  wire [8:0] _T_1105; // @[Math.scala 450:32:@22393.4]
  wire [7:0] x330_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 329:29:@21983.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:408:@22004.4]
  wire [9:0] _GEN_6; // @[Math.scala 450:32:@22398.4]
  wire [9:0] _T_1109; // @[Math.scala 450:32:@22398.4]
  wire [7:0] x335_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 346:29:@22041.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:408:@22062.4]
  wire [8:0] _GEN_7; // @[Math.scala 450:32:@22403.4]
  wire [8:0] _T_1113; // @[Math.scala 450:32:@22403.4]
  wire [7:0] x356_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 407:29:@22262.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:408:@22283.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@22408.4]
  wire [8:0] _T_1117; // @[Math.scala 450:32:@22408.4]
  wire [7:0] x380_sum_number; // @[Math.scala 154:22:@22560.4 Math.scala 155:14:@22561.4]
  wire [3:0] _T_1174; // @[FixedPoint.scala 18:52:@22566.4]
  wire [7:0] x305_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 242:29:@21676.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:338:@21697.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@22579.4]
  wire [8:0] _T_1181; // @[Math.scala 450:32:@22579.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@22584.4]
  wire [8:0] _T_1185; // @[Math.scala 450:32:@22584.4]
  wire [9:0] _GEN_11; // @[Math.scala 450:32:@22589.4]
  wire [9:0] _T_1189; // @[Math.scala 450:32:@22589.4]
  wire [7:0] x340_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 363:29:@22099.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:408:@22120.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@22594.4]
  wire [8:0] _T_1193; // @[Math.scala 450:32:@22594.4]
  wire [7:0] x361_rd_0_number; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 430:29:@22313.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:408:@22334.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@22599.4]
  wire [8:0] _T_1197; // @[Math.scala 450:32:@22599.4]
  wire [7:0] x394_sum_number; // @[Math.scala 154:22:@22753.4 Math.scala 155:14:@22754.4]
  wire [3:0] _T_1256; // @[FixedPoint.scala 18:52:@22759.4]
  wire [7:0] x541_x381_D1_number; // @[package.scala 96:25:@22785.4 package.scala 96:25:@22786.4]
  wire [7:0] x540_x395_D1_number; // @[package.scala 96:25:@22776.4 package.scala 96:25:@22777.4]
  wire  _T_1287; // @[package.scala 96:25:@22827.4 package.scala 96:25:@22828.4]
  wire  _T_1289; // @[implicits.scala 55:10:@22829.4]
  wire  x542_b255_D34; // @[package.scala 96:25:@22809.4 package.scala 96:25:@22810.4]
  wire  _T_1290; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 561:117:@22830.4]
  wire  x543_b256_D34; // @[package.scala 96:25:@22818.4 package.scala 96:25:@22819.4]
  wire  _T_1291; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 561:123:@22831.4]
  wire [31:0] x477_x468_D2_number; // @[package.scala 96:25:@21145.4 package.scala 96:25:@21146.4]
  wire [31:0] x481_x272_sum_D1_number; // @[package.scala 96:25:@21181.4 package.scala 96:25:@21182.4]
  wire [31:0] x482_x469_D2_number; // @[package.scala 96:25:@21190.4 package.scala 96:25:@21191.4]
  wire [31:0] x278_sum_number; // @[Math.scala 154:22:@21266.4 Math.scala 155:14:@21267.4]
  wire [31:0] x485_x470_D1_number; // @[package.scala 96:25:@21284.4 package.scala 96:25:@21285.4]
  wire [31:0] x490_x289_sum_D1_number; // @[package.scala 96:25:@21419.4 package.scala 96:25:@21420.4]
  wire [31:0] x492_x471_D2_number; // @[package.scala 96:25:@21437.4 package.scala 96:25:@21438.4]
  wire [31:0] x495_x470_D22_number; // @[package.scala 96:25:@21464.4 package.scala 96:25:@21465.4]
  wire [31:0] x498_x295_sum_D1_number; // @[package.scala 96:25:@21540.4 package.scala 96:25:@21541.4]
  wire [31:0] x500_x469_D23_number; // @[package.scala 96:25:@21558.4 package.scala 96:25:@21559.4]
  wire [31:0] x502_x472_D17_number; // @[package.scala 96:25:@21655.4 package.scala 96:25:@21656.4]
  wire [31:0] x504_x304_sum_D1_number; // @[package.scala 96:25:@21673.4 package.scala 96:25:@21674.4]
  wire [31:0] x506_x313_sum_D1_number; // @[package.scala 96:25:@21770.4 package.scala 96:25:@21771.4]
  wire [31:0] x507_x473_D17_number; // @[package.scala 96:25:@21779.4 package.scala 96:25:@21780.4]
  wire [31:0] x324_sum_number; // @[Math.scala 154:22:@21895.4 Math.scala 155:14:@21896.4]
  wire [31:0] x511_x474_D1_number; // @[package.scala 96:25:@21913.4 package.scala 96:25:@21914.4]
  wire [31:0] x329_sum_number; // @[Math.scala 154:22:@21971.4 Math.scala 155:14:@21972.4]
  wire [31:0] x334_sum_number; // @[Math.scala 154:22:@22029.4 Math.scala 155:14:@22030.4]
  wire [31:0] x339_sum_number; // @[Math.scala 154:22:@22087.4 Math.scala 155:14:@22088.4]
  wire [31:0] x350_sum_number; // @[Math.scala 154:22:@22192.4 Math.scala 155:14:@22193.4]
  wire [31:0] x519_x475_D1_number; // @[package.scala 96:25:@22201.4 package.scala 96:25:@22202.4]
  wire [31:0] x355_sum_number; // @[Math.scala 154:22:@22250.4 Math.scala 155:14:@22251.4]
  wire [31:0] x360_sum_number; // @[Math.scala 154:22:@22301.4 Math.scala 155:14:@22302.4]
  wire [31:0] x365_sum_number; // @[Math.scala 154:22:@22350.4 Math.scala 155:14:@22351.4]
  _ _ ( // @[Math.scala 709:24:@20890.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@20902.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x257_lb_0 x257_lb_0 ( // @[m_x257_lb_0.scala 39:17:@20912.4]
    .clock(x257_lb_0_clock),
    .reset(x257_lb_0_reset),
    .io_rPort_11_banks_1(x257_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x257_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x257_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x257_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x257_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x257_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x257_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x257_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x257_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x257_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x257_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x257_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x257_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x257_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x257_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x257_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x257_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x257_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x257_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x257_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x257_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x257_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x257_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x257_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x257_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x257_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x257_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x257_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x257_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x257_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x257_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x257_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x257_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x257_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x257_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x257_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x257_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x257_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x257_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x257_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x257_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x257_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x257_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x257_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x257_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x257_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x257_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x257_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x257_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x257_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x257_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x257_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x257_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x257_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x257_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x257_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x257_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x257_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x257_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x257_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x257_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x257_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x257_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x257_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x257_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x257_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x257_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x257_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x257_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x257_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x257_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x257_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x257_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x257_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x257_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x257_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x257_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x257_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x257_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x257_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x257_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x257_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_132 RetimeWrapper ( // @[package.scala 93:22:@21018.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x272_sum x272_sum_1 ( // @[Math.scala 150:24:@21130.4]
    .clock(x272_sum_1_clock),
    .reset(x272_sum_1_reset),
    .io_a(x272_sum_1_io_a),
    .io_b(x272_sum_1_io_b),
    .io_flow(x272_sum_1_io_flow),
    .io_result(x272_sum_1_io_result)
  );
  RetimeWrapper_134 RetimeWrapper_1 ( // @[package.scala 93:22:@21140.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_2 ( // @[package.scala 93:22:@21149.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_3 ( // @[package.scala 93:22:@21158.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_4 ( // @[package.scala 93:22:@21167.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_133 RetimeWrapper_5 ( // @[package.scala 93:22:@21176.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_134 RetimeWrapper_6 ( // @[package.scala 93:22:@21185.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_7 ( // @[package.scala 93:22:@21196.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x272_sum x274_rdcol_1 ( // @[Math.scala 150:24:@21219.4]
    .clock(x274_rdcol_1_clock),
    .reset(x274_rdcol_1_reset),
    .io_a(x274_rdcol_1_io_a),
    .io_b(x274_rdcol_1_io_b),
    .io_flow(x274_rdcol_1_io_flow),
    .io_result(x274_rdcol_1_io_result)
  );
  RetimeWrapper_133 RetimeWrapper_8 ( // @[package.scala 93:22:@21251.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x272_sum x278_sum_1 ( // @[Math.scala 150:24:@21260.4]
    .clock(x278_sum_1_clock),
    .reset(x278_sum_1_reset),
    .io_a(x278_sum_1_io_a),
    .io_b(x278_sum_1_io_b),
    .io_flow(x278_sum_1_io_flow),
    .io_result(x278_sum_1_io_result)
  );
  RetimeWrapper_136 RetimeWrapper_9 ( // @[package.scala 93:22:@21270.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_133 RetimeWrapper_10 ( // @[package.scala 93:22:@21279.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_11 ( // @[package.scala 93:22:@21290.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_147 RetimeWrapper_12 ( // @[package.scala 93:22:@21311.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  x281 x281_1 ( // @[Math.scala 366:24:@21322.4]
    .clock(x281_1_clock),
    .reset(x281_1_reset),
    .io_a(x281_1_io_a),
    .io_flow(x281_1_io_flow),
    .io_result(x281_1_io_result)
  );
  RetimeWrapper_147 RetimeWrapper_13 ( // @[package.scala 93:22:@21339.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@21355.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_151 RetimeWrapper_15 ( // @[package.scala 93:22:@21395.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  x272_sum x289_sum_1 ( // @[Math.scala 150:24:@21404.4]
    .clock(x289_sum_1_clock),
    .reset(x289_sum_1_reset),
    .io_a(x289_sum_1_io_a),
    .io_b(x289_sum_1_io_b),
    .io_flow(x289_sum_1_io_flow),
    .io_result(x289_sum_1_io_result)
  );
  RetimeWrapper_133 RetimeWrapper_16 ( // @[package.scala 93:22:@21414.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_154 RetimeWrapper_17 ( // @[package.scala 93:22:@21423.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_134 RetimeWrapper_18 ( // @[package.scala 93:22:@21432.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_19 ( // @[package.scala 93:22:@21441.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_20 ( // @[package.scala 93:22:@21450.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_158 RetimeWrapper_21 ( // @[package.scala 93:22:@21459.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_22 ( // @[package.scala 93:22:@21471.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_147 RetimeWrapper_23 ( // @[package.scala 93:22:@21492.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_161 RetimeWrapper_24 ( // @[package.scala 93:22:@21516.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x272_sum x295_sum_1 ( // @[Math.scala 150:24:@21525.4]
    .clock(x295_sum_1_clock),
    .reset(x295_sum_1_reset),
    .io_a(x295_sum_1_io_a),
    .io_b(x295_sum_1_io_b),
    .io_flow(x295_sum_1_io_flow),
    .io_result(x295_sum_1_io_result)
  );
  RetimeWrapper_133 RetimeWrapper_25 ( // @[package.scala 93:22:@21535.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_164 RetimeWrapper_26 ( // @[package.scala 93:22:@21544.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_27 ( // @[package.scala 93:22:@21553.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_28 ( // @[package.scala 93:22:@21565.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x272_sum x298_rdcol_1 ( // @[Math.scala 150:24:@21588.4]
    .clock(x298_rdcol_1_clock),
    .reset(x298_rdcol_1_reset),
    .io_a(x298_rdcol_1_io_a),
    .io_b(x298_rdcol_1_io_b),
    .io_flow(x298_rdcol_1_io_flow),
    .io_result(x298_rdcol_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_29 ( // @[package.scala 93:22:@21631.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  x272_sum x304_sum_1 ( // @[Math.scala 150:24:@21640.4]
    .clock(x304_sum_1_clock),
    .reset(x304_sum_1_reset),
    .io_a(x304_sum_1_io_a),
    .io_b(x304_sum_1_io_b),
    .io_flow(x304_sum_1_io_flow),
    .io_result(x304_sum_1_io_result)
  );
  RetimeWrapper_170 RetimeWrapper_30 ( // @[package.scala 93:22:@21650.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_154 RetimeWrapper_31 ( // @[package.scala 93:22:@21659.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_133 RetimeWrapper_32 ( // @[package.scala 93:22:@21668.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_33 ( // @[package.scala 93:22:@21680.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  x272_sum x307_rdcol_1 ( // @[Math.scala 150:24:@21703.4]
    .clock(x307_rdcol_1_clock),
    .reset(x307_rdcol_1_reset),
    .io_a(x307_rdcol_1_io_a),
    .io_b(x307_rdcol_1_io_b),
    .io_flow(x307_rdcol_1_io_flow),
    .io_result(x307_rdcol_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_34 ( // @[package.scala 93:22:@21746.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x272_sum x313_sum_1 ( // @[Math.scala 150:24:@21755.4]
    .clock(x313_sum_1_clock),
    .reset(x313_sum_1_reset),
    .io_a(x313_sum_1_io_a),
    .io_b(x313_sum_1_io_b),
    .io_flow(x313_sum_1_io_flow),
    .io_result(x313_sum_1_io_result)
  );
  RetimeWrapper_133 RetimeWrapper_35 ( // @[package.scala 93:22:@21765.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_36 ( // @[package.scala 93:22:@21774.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_154 RetimeWrapper_37 ( // @[package.scala 93:22:@21783.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_38 ( // @[package.scala 93:22:@21795.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  x316_rdrow x316_rdrow_1 ( // @[Math.scala 191:24:@21818.4]
    .clock(x316_rdrow_1_clock),
    .reset(x316_rdrow_1_reset),
    .io_a(x316_rdrow_1_io_a),
    .io_b(x316_rdrow_1_io_b),
    .io_flow(x316_rdrow_1_io_flow),
    .io_result(x316_rdrow_1_io_result)
  );
  x281 x317_1 ( // @[Math.scala 366:24:@21830.4]
    .clock(x317_1_clock),
    .reset(x317_1_reset),
    .io_a(x317_1_io_a),
    .io_flow(x317_1_io_flow),
    .io_result(x317_1_io_result)
  );
  RetimeWrapper_161 RetimeWrapper_39 ( // @[package.scala 93:22:@21880.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x272_sum x324_sum_1 ( // @[Math.scala 150:24:@21889.4]
    .clock(x324_sum_1_clock),
    .reset(x324_sum_1_reset),
    .io_a(x324_sum_1_io_a),
    .io_b(x324_sum_1_io_b),
    .io_flow(x324_sum_1_io_flow),
    .io_result(x324_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_40 ( // @[package.scala 93:22:@21899.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_133 RetimeWrapper_41 ( // @[package.scala 93:22:@21908.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_42 ( // @[package.scala 93:22:@21920.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper RetimeWrapper_43 ( // @[package.scala 93:22:@21941.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_158 RetimeWrapper_44 ( // @[package.scala 93:22:@21956.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  x272_sum x329_sum_1 ( // @[Math.scala 150:24:@21965.4]
    .clock(x329_sum_1_clock),
    .reset(x329_sum_1_reset),
    .io_a(x329_sum_1_io_a),
    .io_b(x329_sum_1_io_b),
    .io_flow(x329_sum_1_io_flow),
    .io_result(x329_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_45 ( // @[package.scala 93:22:@21975.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_46 ( // @[package.scala 93:22:@21987.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_47 ( // @[package.scala 93:22:@22014.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  x272_sum x334_sum_1 ( // @[Math.scala 150:24:@22023.4]
    .clock(x334_sum_1_clock),
    .reset(x334_sum_1_reset),
    .io_a(x334_sum_1_io_a),
    .io_b(x334_sum_1_io_b),
    .io_flow(x334_sum_1_io_flow),
    .io_result(x334_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_48 ( // @[package.scala 93:22:@22033.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_49 ( // @[package.scala 93:22:@22045.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_50 ( // @[package.scala 93:22:@22072.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x272_sum x339_sum_1 ( // @[Math.scala 150:24:@22081.4]
    .clock(x339_sum_1_clock),
    .reset(x339_sum_1_reset),
    .io_a(x339_sum_1_io_a),
    .io_b(x339_sum_1_io_b),
    .io_flow(x339_sum_1_io_flow),
    .io_result(x339_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_51 ( // @[package.scala 93:22:@22091.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_52 ( // @[package.scala 93:22:@22103.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x316_rdrow x342_rdrow_1 ( // @[Math.scala 191:24:@22126.4]
    .clock(x342_rdrow_1_clock),
    .reset(x342_rdrow_1_reset),
    .io_a(x342_rdrow_1_io_a),
    .io_b(x342_rdrow_1_io_b),
    .io_flow(x342_rdrow_1_io_flow),
    .io_result(x342_rdrow_1_io_result)
  );
  x281 x343_1 ( // @[Math.scala 366:24:@22138.4]
    .clock(x343_1_clock),
    .reset(x343_1_reset),
    .io_a(x343_1_io_a),
    .io_flow(x343_1_io_flow),
    .io_result(x343_1_io_result)
  );
  x272_sum x350_sum_1 ( // @[Math.scala 150:24:@22186.4]
    .clock(x350_sum_1_clock),
    .reset(x350_sum_1_reset),
    .io_a(x350_sum_1_io_a),
    .io_b(x350_sum_1_io_b),
    .io_flow(x350_sum_1_io_flow),
    .io_result(x350_sum_1_io_result)
  );
  RetimeWrapper_133 RetimeWrapper_53 ( // @[package.scala 93:22:@22196.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_154 RetimeWrapper_54 ( // @[package.scala 93:22:@22205.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_55 ( // @[package.scala 93:22:@22217.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x272_sum x355_sum_1 ( // @[Math.scala 150:24:@22244.4]
    .clock(x355_sum_1_clock),
    .reset(x355_sum_1_reset),
    .io_a(x355_sum_1_io_a),
    .io_b(x355_sum_1_io_b),
    .io_flow(x355_sum_1_io_flow),
    .io_result(x355_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_56 ( // @[package.scala 93:22:@22254.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_57 ( // @[package.scala 93:22:@22266.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x272_sum x360_sum_1 ( // @[Math.scala 150:24:@22295.4]
    .clock(x360_sum_1_clock),
    .reset(x360_sum_1_reset),
    .io_a(x360_sum_1_io_a),
    .io_b(x360_sum_1_io_b),
    .io_flow(x360_sum_1_io_flow),
    .io_result(x360_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_58 ( // @[package.scala 93:22:@22305.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_59 ( // @[package.scala 93:22:@22317.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  x272_sum x365_sum_1 ( // @[Math.scala 150:24:@22344.4]
    .clock(x365_sum_1_clock),
    .reset(x365_sum_1_reset),
    .io_a(x365_sum_1_io_a),
    .io_b(x365_sum_1_io_b),
    .io_flow(x365_sum_1_io_flow),
    .io_result(x365_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_60 ( // @[package.scala 93:22:@22354.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_156 RetimeWrapper_61 ( // @[package.scala 93:22:@22366.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_62 ( // @[package.scala 93:22:@22412.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_63 ( // @[package.scala 93:22:@22421.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x373_x11 x373_x11_1 ( // @[Math.scala 150:24:@22430.4]
    .clock(x373_x11_1_clock),
    .reset(x373_x11_1_reset),
    .io_a(x373_x11_1_io_a),
    .io_b(x373_x11_1_io_b),
    .io_flow(x373_x11_1_io_flow),
    .io_result(x373_x11_1_io_result)
  );
  RetimeWrapper_136 RetimeWrapper_64 ( // @[package.scala 93:22:@22440.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_65 ( // @[package.scala 93:22:@22449.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x373_x11 x374_x12_1 ( // @[Math.scala 150:24:@22458.4]
    .clock(x374_x12_1_clock),
    .reset(x374_x12_1_reset),
    .io_a(x374_x12_1_io_a),
    .io_b(x374_x12_1_io_b),
    .io_flow(x374_x12_1_io_flow),
    .io_result(x374_x12_1_io_result)
  );
  x373_x11 x375_x11_1 ( // @[Math.scala 150:24:@22468.4]
    .clock(x375_x11_1_clock),
    .reset(x375_x11_1_reset),
    .io_a(x375_x11_1_io_a),
    .io_b(x375_x11_1_io_b),
    .io_flow(x375_x11_1_io_flow),
    .io_result(x375_x11_1_io_result)
  );
  x373_x11 x376_x12_1 ( // @[Math.scala 150:24:@22478.4]
    .clock(x376_x12_1_clock),
    .reset(x376_x12_1_reset),
    .io_a(x376_x12_1_io_a),
    .io_b(x376_x12_1_io_b),
    .io_flow(x376_x12_1_io_flow),
    .io_result(x376_x12_1_io_result)
  );
  RetimeWrapper_224 RetimeWrapper_66 ( // @[package.scala 93:22:@22488.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_224 RetimeWrapper_67 ( // @[package.scala 93:22:@22497.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x377_x11 x377_x11_1 ( // @[Math.scala 150:24:@22506.4]
    .io_a(x377_x11_1_io_a),
    .io_b(x377_x11_1_io_b),
    .io_result(x377_x11_1_io_result)
  );
  x377_x11 x378_x12_1 ( // @[Math.scala 150:24:@22516.4]
    .io_a(x378_x12_1_io_a),
    .io_b(x378_x12_1_io_b),
    .io_result(x378_x12_1_io_result)
  );
  RetimeWrapper_226 RetimeWrapper_68 ( // @[package.scala 93:22:@22526.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  x377_x11 x379_x11_1 ( // @[Math.scala 150:24:@22535.4]
    .io_a(x379_x11_1_io_a),
    .io_b(x379_x11_1_io_b),
    .io_result(x379_x11_1_io_result)
  );
  RetimeWrapper_227 RetimeWrapper_69 ( // @[package.scala 93:22:@22545.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x377_x11 x380_sum_1 ( // @[Math.scala 150:24:@22554.4]
    .io_a(x380_sum_1_io_a),
    .io_b(x380_sum_1_io_b),
    .io_result(x380_sum_1_io_result)
  );
  RetimeWrapper_136 RetimeWrapper_70 ( // @[package.scala 93:22:@22568.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_71 ( // @[package.scala 93:22:@22603.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_72 ( // @[package.scala 93:22:@22612.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x373_x11 x387_x11_1 ( // @[Math.scala 150:24:@22621.4]
    .clock(x387_x11_1_clock),
    .reset(x387_x11_1_reset),
    .io_a(x387_x11_1_io_a),
    .io_b(x387_x11_1_io_b),
    .io_flow(x387_x11_1_io_flow),
    .io_result(x387_x11_1_io_result)
  );
  RetimeWrapper_136 RetimeWrapper_73 ( // @[package.scala 93:22:@22631.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_74 ( // @[package.scala 93:22:@22640.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x373_x11 x388_x12_1 ( // @[Math.scala 150:24:@22649.4]
    .clock(x388_x12_1_clock),
    .reset(x388_x12_1_reset),
    .io_a(x388_x12_1_io_a),
    .io_b(x388_x12_1_io_b),
    .io_flow(x388_x12_1_io_flow),
    .io_result(x388_x12_1_io_result)
  );
  x373_x11 x389_x11_1 ( // @[Math.scala 150:24:@22659.4]
    .clock(x389_x11_1_clock),
    .reset(x389_x11_1_reset),
    .io_a(x389_x11_1_io_a),
    .io_b(x389_x11_1_io_b),
    .io_flow(x389_x11_1_io_flow),
    .io_result(x389_x11_1_io_result)
  );
  x373_x11 x390_x12_1 ( // @[Math.scala 150:24:@22669.4]
    .clock(x390_x12_1_clock),
    .reset(x390_x12_1_reset),
    .io_a(x390_x12_1_io_a),
    .io_b(x390_x12_1_io_b),
    .io_flow(x390_x12_1_io_flow),
    .io_result(x390_x12_1_io_result)
  );
  RetimeWrapper_224 RetimeWrapper_75 ( // @[package.scala 93:22:@22679.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_224 RetimeWrapper_76 ( // @[package.scala 93:22:@22688.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x377_x11 x391_x11_1 ( // @[Math.scala 150:24:@22699.4]
    .io_a(x391_x11_1_io_a),
    .io_b(x391_x11_1_io_b),
    .io_result(x391_x11_1_io_result)
  );
  x377_x11 x392_x12_1 ( // @[Math.scala 150:24:@22709.4]
    .io_a(x392_x12_1_io_a),
    .io_b(x392_x12_1_io_b),
    .io_result(x392_x12_1_io_result)
  );
  RetimeWrapper_226 RetimeWrapper_77 ( // @[package.scala 93:22:@22719.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x377_x11 x393_x11_1 ( // @[Math.scala 150:24:@22728.4]
    .io_a(x393_x11_1_io_a),
    .io_b(x393_x11_1_io_b),
    .io_result(x393_x11_1_io_result)
  );
  RetimeWrapper_227 RetimeWrapper_78 ( // @[package.scala 93:22:@22738.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  x377_x11 x394_sum_1 ( // @[Math.scala 150:24:@22747.4]
    .io_a(x394_sum_1_io_a),
    .io_b(x394_sum_1_io_b),
    .io_result(x394_sum_1_io_result)
  );
  RetimeWrapper_136 RetimeWrapper_79 ( // @[package.scala 93:22:@22761.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_80 ( // @[package.scala 93:22:@22771.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_136 RetimeWrapper_81 ( // @[package.scala 93:22:@22780.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_82 ( // @[package.scala 93:22:@22795.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_83 ( // @[package.scala 93:22:@22804.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_84 ( // @[package.scala 93:22:@22813.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_85 ( // @[package.scala 93:22:@22822.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  assign b255 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 62:18:@20910.4]
  assign b256 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 63:18:@20911.4]
  assign _T_206 = b255 & b256; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 68:30:@21006.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 68:37:@21007.4]
  assign _T_211 = io_in_x244_TID == 8'h0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 70:76:@21012.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 70:62:@21013.4]
  assign _T_214 = io_in_x244_TDEST == 8'h0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 70:101:@21014.4]
  assign x476_x258_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@21023.4 package.scala 96:25:@21024.4]
  assign b253_number = __io_result; // @[Math.scala 712:22:@20895.4 Math.scala 713:14:@20896.4]
  assign _T_242 = $signed(b253_number); // @[Math.scala 499:52:@21039.4]
  assign x262 = $signed(32'sh1) == $signed(_T_242); // @[Math.scala 499:44:@21047.4]
  assign x263 = $signed(32'sh2) == $signed(_T_242); // @[Math.scala 499:44:@21054.4]
  assign x264 = $signed(32'sh3) == $signed(_T_242); // @[Math.scala 499:44:@21061.4]
  assign _T_289 = x262 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@21073.4]
  assign _T_291 = x263 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@21074.4]
  assign _T_293 = x264 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@21075.4]
  assign _T_295 = _T_289 | _T_291; // @[Mux.scala 19:72:@21077.4]
  assign x265_number = _T_295 | _T_293; // @[Mux.scala 19:72:@21078.4]
  assign _T_307 = $signed(x265_number); // @[Math.scala 406:49:@21088.4]
  assign _T_309 = $signed(_T_307) & $signed(32'sh3); // @[Math.scala 406:56:@21090.4]
  assign _T_310 = $signed(_T_309); // @[Math.scala 406:56:@21091.4]
  assign b254_number = __1_io_result; // @[Math.scala 712:22:@20907.4 Math.scala 713:14:@20908.4]
  assign _T_319 = $signed(b254_number); // @[Math.scala 406:49:@21099.4]
  assign _T_321 = $signed(_T_319) & $signed(32'sh3); // @[Math.scala 406:56:@21101.4]
  assign _T_322 = $signed(_T_321); // @[Math.scala 406:56:@21102.4]
  assign _T_327 = x265_number[31]; // @[FixedPoint.scala 50:25:@21108.4]
  assign _T_331 = _T_327 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21110.4]
  assign _T_332 = x265_number[31:2]; // @[FixedPoint.scala 18:52:@21111.4]
  assign x269_number = {_T_331,_T_332}; // @[Cat.scala 30:58:@21112.4]
  assign _GEN_0 = {{8'd0}, x269_number}; // @[Math.scala 450:32:@21117.4]
  assign _T_337 = _GEN_0 << 8; // @[Math.scala 450:32:@21117.4]
  assign _T_341 = b254_number[31]; // @[FixedPoint.scala 50:25:@21122.4]
  assign _T_345 = _T_341 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21124.4]
  assign _T_346 = b254_number[31:2]; // @[FixedPoint.scala 18:52:@21125.4]
  assign _T_370 = ~ io_sigsIn_break; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:101:@21193.4]
  assign _T_374 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@21201.4 package.scala 96:25:@21202.4]
  assign _T_376 = io_rr ? _T_374 : 1'h0; // @[implicits.scala 55:10:@21203.4]
  assign _T_377 = _T_370 & _T_376; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:118:@21204.4]
  assign _T_379 = _T_377 & _T_370; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:206:@21206.4]
  assign _T_380 = _T_379 & io_sigsIn_backpressure; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:225:@21207.4]
  assign x480_b255_D2 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@21172.4 package.scala 96:25:@21173.4]
  assign _T_381 = _T_380 & x480_b255_D2; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 119:251:@21208.4]
  assign x478_b256_D2 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@21154.4 package.scala 96:25:@21155.4]
  assign x274_rdcol_number = x274_rdcol_1_io_result; // @[Math.scala 154:22:@21225.4 Math.scala 155:14:@21226.4]
  assign _T_398 = $signed(x274_rdcol_number); // @[Math.scala 406:49:@21234.4]
  assign _T_400 = $signed(_T_398) & $signed(32'sh3); // @[Math.scala 406:56:@21236.4]
  assign _T_401 = $signed(_T_400); // @[Math.scala 406:56:@21237.4]
  assign _T_406 = x274_rdcol_number[31]; // @[FixedPoint.scala 50:25:@21243.4]
  assign _T_410 = _T_406 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21245.4]
  assign _T_411 = x274_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@21246.4]
  assign _T_430 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@21295.4 package.scala 96:25:@21296.4]
  assign _T_432 = io_rr ? _T_430 : 1'h0; // @[implicits.scala 55:10:@21297.4]
  assign _T_433 = _T_370 & _T_432; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:118:@21298.4]
  assign _T_435 = _T_433 & _T_370; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:206:@21300.4]
  assign _T_436 = _T_435 & io_sigsIn_backpressure; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:225:@21301.4]
  assign _T_437 = _T_436 & x480_b255_D2; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 140:251:@21302.4]
  assign x486_b253_D5_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@21316.4 package.scala 96:25:@21317.4]
  assign _T_454 = $signed(x486_b253_D5_number); // @[Math.scala 465:37:@21334.4]
  assign x282 = $signed(_T_454) < $signed(32'sh0); // @[Math.scala 465:44:@21336.4]
  assign x487_x274_rdcol_D5_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@21344.4 package.scala 96:25:@21345.4]
  assign _T_465 = $signed(x487_x274_rdcol_D5_number); // @[Math.scala 465:37:@21350.4]
  assign x283 = $signed(_T_465) < $signed(32'sh0); // @[Math.scala 465:44:@21352.4]
  assign x488_x282_D1 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@21360.4 package.scala 96:25:@21361.4]
  assign x284 = x488_x282_D1 | x283; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 155:24:@21364.4]
  assign x281_number = x281_1_io_result; // @[Math.scala 370:22:@21328.4 Math.scala 371:14:@21329.4]
  assign _T_482 = $signed(x281_number); // @[Math.scala 406:49:@21373.4]
  assign _T_484 = $signed(_T_482) & $signed(32'sh3); // @[Math.scala 406:56:@21375.4]
  assign _T_485 = $signed(_T_484); // @[Math.scala 406:56:@21376.4]
  assign _T_490 = x281_number[31]; // @[FixedPoint.scala 50:25:@21382.4]
  assign _T_494 = _T_490 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21384.4]
  assign _T_495 = x281_number[31:2]; // @[FixedPoint.scala 18:52:@21385.4]
  assign x287_number = {_T_494,_T_495}; // @[Cat.scala 30:58:@21386.4]
  assign _GEN_1 = {{8'd0}, x287_number}; // @[Math.scala 450:32:@21391.4]
  assign _T_500 = _GEN_1 << 8; // @[Math.scala 450:32:@21391.4]
  assign _T_536 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@21476.4 package.scala 96:25:@21477.4]
  assign _T_538 = io_rr ? _T_536 : 1'h0; // @[implicits.scala 55:10:@21478.4]
  assign _T_539 = _T_370 & _T_538; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 190:194:@21479.4]
  assign x491_x285_D17 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@21428.4 package.scala 96:25:@21429.4]
  assign _T_540 = _T_539 & x491_x285_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 190:283:@21480.4]
  assign x494_b255_D23 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@21455.4 package.scala 96:25:@21456.4]
  assign _T_541 = _T_540 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 190:326:@21481.4]
  assign x493_b256_D23 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@21446.4 package.scala 96:25:@21447.4]
  assign x496_b254_D5_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@21497.4 package.scala 96:25:@21498.4]
  assign _T_554 = $signed(x496_b254_D5_number); // @[Math.scala 465:37:@21505.4]
  assign x292 = $signed(_T_554) < $signed(32'sh0); // @[Math.scala 465:44:@21507.4]
  assign x293 = x282 | x292; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 200:59:@21510.4]
  assign _T_587 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@21570.4 package.scala 96:25:@21571.4]
  assign _T_589 = io_rr ? _T_587 : 1'h0; // @[implicits.scala 55:10:@21572.4]
  assign _T_590 = _T_370 & _T_589; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:194:@21573.4]
  assign x499_x294_D18 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@21549.4 package.scala 96:25:@21550.4]
  assign _T_591 = _T_590 & x499_x294_D18; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:283:@21574.4]
  assign _T_592 = _T_591 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:291:@21575.4]
  assign x298_rdcol_number = x298_rdcol_1_io_result; // @[Math.scala 154:22:@21594.4 Math.scala 155:14:@21595.4]
  assign _T_607 = $signed(x298_rdcol_number); // @[Math.scala 465:37:@21600.4]
  assign x299 = $signed(_T_607) < $signed(32'sh0); // @[Math.scala 465:44:@21602.4]
  assign x300 = x488_x282_D1 | x299; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 225:59:@21605.4]
  assign _T_623 = $signed(_T_607) & $signed(32'sh3); // @[Math.scala 406:56:@21616.4]
  assign _T_624 = $signed(_T_623); // @[Math.scala 406:56:@21617.4]
  assign _T_629 = x298_rdcol_number[31]; // @[FixedPoint.scala 50:25:@21623.4]
  assign _T_633 = _T_629 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21625.4]
  assign _T_634 = x298_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@21626.4]
  assign _T_662 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@21685.4 package.scala 96:25:@21686.4]
  assign _T_664 = io_rr ? _T_662 : 1'h0; // @[implicits.scala 55:10:@21687.4]
  assign _T_665 = _T_370 & _T_664; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:194:@21688.4]
  assign x503_x301_D17 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@21664.4 package.scala 96:25:@21665.4]
  assign _T_666 = _T_665 & x503_x301_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:283:@21689.4]
  assign _T_667 = _T_666 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:291:@21690.4]
  assign x307_rdcol_number = x307_rdcol_1_io_result; // @[Math.scala 154:22:@21709.4 Math.scala 155:14:@21710.4]
  assign _T_682 = $signed(x307_rdcol_number); // @[Math.scala 465:37:@21715.4]
  assign x308 = $signed(_T_682) < $signed(32'sh0); // @[Math.scala 465:44:@21717.4]
  assign x309 = x488_x282_D1 | x308; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 254:59:@21720.4]
  assign _T_698 = $signed(_T_682) & $signed(32'sh3); // @[Math.scala 406:56:@21731.4]
  assign _T_699 = $signed(_T_698); // @[Math.scala 406:56:@21732.4]
  assign _T_704 = x307_rdcol_number[31]; // @[FixedPoint.scala 50:25:@21738.4]
  assign _T_708 = _T_704 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21740.4]
  assign _T_709 = x307_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@21741.4]
  assign _T_737 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@21800.4 package.scala 96:25:@21801.4]
  assign _T_739 = io_rr ? _T_737 : 1'h0; // @[implicits.scala 55:10:@21802.4]
  assign _T_740 = _T_370 & _T_739; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 275:194:@21803.4]
  assign x508_x310_D17 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@21788.4 package.scala 96:25:@21789.4]
  assign _T_741 = _T_740 & x508_x310_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 275:283:@21804.4]
  assign _T_742 = _T_741 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 275:291:@21805.4]
  assign x316_rdrow_number = x316_rdrow_1_io_result; // @[Math.scala 195:22:@21824.4 Math.scala 196:14:@21825.4]
  assign _T_764 = $signed(x316_rdrow_number); // @[Math.scala 465:37:@21842.4]
  assign x318 = $signed(_T_764) < $signed(32'sh0); // @[Math.scala 465:44:@21844.4]
  assign x319 = x318 | x283; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 285:24:@21847.4]
  assign x317_number = x317_1_io_result; // @[Math.scala 370:22:@21836.4 Math.scala 371:14:@21837.4]
  assign _T_778 = $signed(x317_number); // @[Math.scala 406:49:@21856.4]
  assign _T_780 = $signed(_T_778) & $signed(32'sh3); // @[Math.scala 406:56:@21858.4]
  assign _T_781 = $signed(_T_780); // @[Math.scala 406:56:@21859.4]
  assign _T_788 = x317_number[31]; // @[FixedPoint.scala 50:25:@21867.4]
  assign _T_792 = _T_788 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21869.4]
  assign _T_793 = x317_number[31:2]; // @[FixedPoint.scala 18:52:@21870.4]
  assign x322_number = {_T_792,_T_793}; // @[Cat.scala 30:58:@21871.4]
  assign _GEN_2 = {{8'd0}, x322_number}; // @[Math.scala 450:32:@21876.4]
  assign _T_798 = _GEN_2 << 8; // @[Math.scala 450:32:@21876.4]
  assign _T_822 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@21925.4 package.scala 96:25:@21926.4]
  assign _T_824 = io_rr ? _T_822 : 1'h0; // @[implicits.scala 55:10:@21927.4]
  assign _T_825 = _T_370 & _T_824; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:194:@21928.4]
  assign x510_x320_D17 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@21904.4 package.scala 96:25:@21905.4]
  assign _T_826 = _T_825 & x510_x320_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:283:@21929.4]
  assign _T_827 = _T_826 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:291:@21930.4]
  assign x512_x292_D1 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@21946.4 package.scala 96:25:@21947.4]
  assign x327 = x318 | x512_x292_D1; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 320:59:@21950.4]
  assign _T_857 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@21992.4 package.scala 96:25:@21993.4]
  assign _T_859 = io_rr ? _T_857 : 1'h0; // @[implicits.scala 55:10:@21994.4]
  assign _T_860 = _T_370 & _T_859; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:194:@21995.4]
  assign x514_x328_D17 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@21980.4 package.scala 96:25:@21981.4]
  assign _T_861 = _T_860 & x514_x328_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:283:@21996.4]
  assign _T_862 = _T_861 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:291:@21997.4]
  assign x332 = x318 | x299; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 337:59:@22008.4]
  assign _T_889 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@22050.4 package.scala 96:25:@22051.4]
  assign _T_891 = io_rr ? _T_889 : 1'h0; // @[implicits.scala 55:10:@22052.4]
  assign _T_892 = _T_370 & _T_891; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:194:@22053.4]
  assign x516_x333_D17 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@22038.4 package.scala 96:25:@22039.4]
  assign _T_893 = _T_892 & x516_x333_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:283:@22054.4]
  assign _T_894 = _T_893 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:291:@22055.4]
  assign x337 = x318 | x308; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 354:59:@22066.4]
  assign _T_921 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@22108.4 package.scala 96:25:@22109.4]
  assign _T_923 = io_rr ? _T_921 : 1'h0; // @[implicits.scala 55:10:@22110.4]
  assign _T_924 = _T_370 & _T_923; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:194:@22111.4]
  assign x518_x338_D17 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@22096.4 package.scala 96:25:@22097.4]
  assign _T_925 = _T_924 & x518_x338_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:283:@22112.4]
  assign _T_926 = _T_925 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:291:@22113.4]
  assign x342_rdrow_number = x342_rdrow_1_io_result; // @[Math.scala 195:22:@22132.4 Math.scala 196:14:@22133.4]
  assign _T_948 = $signed(x342_rdrow_number); // @[Math.scala 465:37:@22150.4]
  assign x344 = $signed(_T_948) < $signed(32'sh0); // @[Math.scala 465:44:@22152.4]
  assign x345 = x344 | x283; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 377:24:@22155.4]
  assign x343_number = x343_1_io_result; // @[Math.scala 370:22:@22144.4 Math.scala 371:14:@22145.4]
  assign _T_962 = $signed(x343_number); // @[Math.scala 406:49:@22164.4]
  assign _T_964 = $signed(_T_962) & $signed(32'sh3); // @[Math.scala 406:56:@22166.4]
  assign _T_965 = $signed(_T_964); // @[Math.scala 406:56:@22167.4]
  assign _T_970 = x343_number[31]; // @[FixedPoint.scala 50:25:@22173.4]
  assign _T_974 = _T_970 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@22175.4]
  assign _T_975 = x343_number[31:2]; // @[FixedPoint.scala 18:52:@22176.4]
  assign x348_number = {_T_974,_T_975}; // @[Cat.scala 30:58:@22177.4]
  assign _GEN_3 = {{8'd0}, x348_number}; // @[Math.scala 450:32:@22182.4]
  assign _T_980 = _GEN_3 << 8; // @[Math.scala 450:32:@22182.4]
  assign _T_1001 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@22222.4 package.scala 96:25:@22223.4]
  assign _T_1003 = io_rr ? _T_1001 : 1'h0; // @[implicits.scala 55:10:@22224.4]
  assign _T_1004 = _T_370 & _T_1003; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 396:194:@22225.4]
  assign x520_x346_D17 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@22210.4 package.scala 96:25:@22211.4]
  assign _T_1005 = _T_1004 & x520_x346_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 396:283:@22226.4]
  assign _T_1006 = _T_1005 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 396:291:@22227.4]
  assign x353 = x344 | x512_x292_D1; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 400:24:@22238.4]
  assign _T_1030 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@22271.4 package.scala 96:25:@22272.4]
  assign _T_1032 = io_rr ? _T_1030 : 1'h0; // @[implicits.scala 55:10:@22273.4]
  assign _T_1033 = _T_370 & _T_1032; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:194:@22274.4]
  assign x521_x354_D17 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@22259.4 package.scala 96:25:@22260.4]
  assign _T_1034 = _T_1033 & x521_x354_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:283:@22275.4]
  assign _T_1035 = _T_1034 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:291:@22276.4]
  assign x358 = x344 | x299; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 421:59:@22287.4]
  assign _T_1061 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@22322.4 package.scala 96:25:@22323.4]
  assign _T_1063 = io_rr ? _T_1061 : 1'h0; // @[implicits.scala 55:10:@22324.4]
  assign _T_1064 = _T_370 & _T_1063; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:194:@22325.4]
  assign x522_x359_D17 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@22310.4 package.scala 96:25:@22311.4]
  assign _T_1065 = _T_1064 & x522_x359_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:283:@22326.4]
  assign _T_1066 = _T_1065 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:291:@22327.4]
  assign x363 = x344 | x308; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 438:59:@22338.4]
  assign _T_1090 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@22371.4 package.scala 96:25:@22372.4]
  assign _T_1092 = io_rr ? _T_1090 : 1'h0; // @[implicits.scala 55:10:@22373.4]
  assign _T_1093 = _T_370 & _T_1092; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 449:194:@22374.4]
  assign x523_x364_D17 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@22359.4 package.scala 96:25:@22360.4]
  assign _T_1094 = _T_1093 & x523_x364_D17; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 449:283:@22375.4]
  assign _T_1095 = _T_1094 & x494_b255_D23; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 449:291:@22376.4]
  assign x296_rd_0_number = x257_lb_0_io_rPort_5_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 213:29:@21561.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 217:338:@21582.4]
  assign _GEN_4 = {{1'd0}, x296_rd_0_number}; // @[Math.scala 450:32:@22388.4]
  assign _T_1101 = _GEN_4 << 1; // @[Math.scala 450:32:@22388.4]
  assign x325_rd_0_number = x257_lb_0_io_rPort_1_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 310:29:@21916.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 314:408:@21937.4]
  assign _GEN_5 = {{1'd0}, x325_rd_0_number}; // @[Math.scala 450:32:@22393.4]
  assign _T_1105 = _GEN_5 << 1; // @[Math.scala 450:32:@22393.4]
  assign x330_rd_0_number = x257_lb_0_io_rPort_7_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 329:29:@21983.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 333:408:@22004.4]
  assign _GEN_6 = {{2'd0}, x330_rd_0_number}; // @[Math.scala 450:32:@22398.4]
  assign _T_1109 = _GEN_6 << 2; // @[Math.scala 450:32:@22398.4]
  assign x335_rd_0_number = x257_lb_0_io_rPort_6_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 346:29:@22041.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 350:408:@22062.4]
  assign _GEN_7 = {{1'd0}, x335_rd_0_number}; // @[Math.scala 450:32:@22403.4]
  assign _T_1113 = _GEN_7 << 1; // @[Math.scala 450:32:@22403.4]
  assign x356_rd_0_number = x257_lb_0_io_rPort_4_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 407:29:@22262.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 411:408:@22283.4]
  assign _GEN_8 = {{1'd0}, x356_rd_0_number}; // @[Math.scala 450:32:@22408.4]
  assign _T_1117 = _GEN_8 << 1; // @[Math.scala 450:32:@22408.4]
  assign x380_sum_number = x380_sum_1_io_result; // @[Math.scala 154:22:@22560.4 Math.scala 155:14:@22561.4]
  assign _T_1174 = x380_sum_number[7:4]; // @[FixedPoint.scala 18:52:@22566.4]
  assign x305_rd_0_number = x257_lb_0_io_rPort_11_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 242:29:@21676.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 246:338:@21697.4]
  assign _GEN_9 = {{1'd0}, x305_rd_0_number}; // @[Math.scala 450:32:@22579.4]
  assign _T_1181 = _GEN_9 << 1; // @[Math.scala 450:32:@22579.4]
  assign _GEN_10 = {{1'd0}, x330_rd_0_number}; // @[Math.scala 450:32:@22584.4]
  assign _T_1185 = _GEN_10 << 1; // @[Math.scala 450:32:@22584.4]
  assign _GEN_11 = {{2'd0}, x335_rd_0_number}; // @[Math.scala 450:32:@22589.4]
  assign _T_1189 = _GEN_11 << 2; // @[Math.scala 450:32:@22589.4]
  assign x340_rd_0_number = x257_lb_0_io_rPort_0_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 363:29:@22099.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 367:408:@22120.4]
  assign _GEN_12 = {{1'd0}, x340_rd_0_number}; // @[Math.scala 450:32:@22594.4]
  assign _T_1193 = _GEN_12 << 1; // @[Math.scala 450:32:@22594.4]
  assign x361_rd_0_number = x257_lb_0_io_rPort_3_output_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 430:29:@22313.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 434:408:@22334.4]
  assign _GEN_13 = {{1'd0}, x361_rd_0_number}; // @[Math.scala 450:32:@22599.4]
  assign _T_1197 = _GEN_13 << 1; // @[Math.scala 450:32:@22599.4]
  assign x394_sum_number = x394_sum_1_io_result; // @[Math.scala 154:22:@22753.4 Math.scala 155:14:@22754.4]
  assign _T_1256 = x394_sum_number[7:4]; // @[FixedPoint.scala 18:52:@22759.4]
  assign x541_x381_D1_number = RetimeWrapper_81_io_out; // @[package.scala 96:25:@22785.4 package.scala 96:25:@22786.4]
  assign x540_x395_D1_number = RetimeWrapper_80_io_out; // @[package.scala 96:25:@22776.4 package.scala 96:25:@22777.4]
  assign _T_1287 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@22827.4 package.scala 96:25:@22828.4]
  assign _T_1289 = io_rr ? _T_1287 : 1'h0; // @[implicits.scala 55:10:@22829.4]
  assign x542_b255_D34 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@22809.4 package.scala 96:25:@22810.4]
  assign _T_1290 = _T_1289 & x542_b255_D34; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 561:117:@22830.4]
  assign x543_b256_D34 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@22818.4 package.scala 96:25:@22819.4]
  assign _T_1291 = _T_1290 & x543_b256_D34; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 561:123:@22831.4]
  assign x477_x468_D2_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@21145.4 package.scala 96:25:@21146.4]
  assign x481_x272_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@21181.4 package.scala 96:25:@21182.4]
  assign x482_x469_D2_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@21190.4 package.scala 96:25:@21191.4]
  assign x278_sum_number = x278_sum_1_io_result; // @[Math.scala 154:22:@21266.4 Math.scala 155:14:@21267.4]
  assign x485_x470_D1_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@21284.4 package.scala 96:25:@21285.4]
  assign x490_x289_sum_D1_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@21419.4 package.scala 96:25:@21420.4]
  assign x492_x471_D2_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@21437.4 package.scala 96:25:@21438.4]
  assign x495_x470_D22_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@21464.4 package.scala 96:25:@21465.4]
  assign x498_x295_sum_D1_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@21540.4 package.scala 96:25:@21541.4]
  assign x500_x469_D23_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@21558.4 package.scala 96:25:@21559.4]
  assign x502_x472_D17_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@21655.4 package.scala 96:25:@21656.4]
  assign x504_x304_sum_D1_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@21673.4 package.scala 96:25:@21674.4]
  assign x506_x313_sum_D1_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@21770.4 package.scala 96:25:@21771.4]
  assign x507_x473_D17_number = RetimeWrapper_36_io_out; // @[package.scala 96:25:@21779.4 package.scala 96:25:@21780.4]
  assign x324_sum_number = x324_sum_1_io_result; // @[Math.scala 154:22:@21895.4 Math.scala 155:14:@21896.4]
  assign x511_x474_D1_number = RetimeWrapper_41_io_out; // @[package.scala 96:25:@21913.4 package.scala 96:25:@21914.4]
  assign x329_sum_number = x329_sum_1_io_result; // @[Math.scala 154:22:@21971.4 Math.scala 155:14:@21972.4]
  assign x334_sum_number = x334_sum_1_io_result; // @[Math.scala 154:22:@22029.4 Math.scala 155:14:@22030.4]
  assign x339_sum_number = x339_sum_1_io_result; // @[Math.scala 154:22:@22087.4 Math.scala 155:14:@22088.4]
  assign x350_sum_number = x350_sum_1_io_result; // @[Math.scala 154:22:@22192.4 Math.scala 155:14:@22193.4]
  assign x519_x475_D1_number = RetimeWrapper_53_io_out; // @[package.scala 96:25:@22201.4 package.scala 96:25:@22202.4]
  assign x355_sum_number = x355_sum_1_io_result; // @[Math.scala 154:22:@22250.4 Math.scala 155:14:@22251.4]
  assign x360_sum_number = x360_sum_1_io_result; // @[Math.scala 154:22:@22301.4 Math.scala 155:14:@22302.4]
  assign x365_sum_number = x365_sum_1_io_result; // @[Math.scala 154:22:@22350.4 Math.scala 155:14:@22351.4]
  assign io_in_x244_TREADY = _T_212 & _T_214; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 68:22:@21008.4 sm_x400_inr_Foreach_SAMPLER_BOX.scala 70:22:@21016.4]
  assign io_in_x245_TVALID = _T_1291 & io_sigsIn_backpressure; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 561:22:@22833.4]
  assign io_in_x245_TDATA = {{240'd0}, RetimeWrapper_82_io_out}; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 562:24:@22834.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@20893.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@20905.4]
  assign x257_lb_0_clock = clock; // @[:@20913.4]
  assign x257_lb_0_reset = reset; // @[:@20914.4]
  assign x257_lb_0_io_rPort_11_banks_1 = x502_x472_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@21693.4]
  assign x257_lb_0_io_rPort_11_banks_0 = x492_x471_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21692.4]
  assign x257_lb_0_io_rPort_11_ofs_0 = x504_x304_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@21694.4]
  assign x257_lb_0_io_rPort_11_en_0 = _T_667 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@21696.4]
  assign x257_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21695.4]
  assign x257_lb_0_io_rPort_10_banks_1 = x495_x470_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@21484.4]
  assign x257_lb_0_io_rPort_10_banks_0 = x492_x471_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21483.4]
  assign x257_lb_0_io_rPort_10_ofs_0 = x490_x289_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@21485.4]
  assign x257_lb_0_io_rPort_10_en_0 = _T_541 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@21487.4]
  assign x257_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21486.4]
  assign x257_lb_0_io_rPort_9_banks_1 = x495_x470_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@22230.4]
  assign x257_lb_0_io_rPort_9_banks_0 = x519_x475_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@22229.4]
  assign x257_lb_0_io_rPort_9_ofs_0 = x350_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@22231.4]
  assign x257_lb_0_io_rPort_9_en_0 = _T_1006 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@22233.4]
  assign x257_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@22232.4]
  assign x257_lb_0_io_rPort_8_banks_1 = x507_x473_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@21808.4]
  assign x257_lb_0_io_rPort_8_banks_0 = x492_x471_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21807.4]
  assign x257_lb_0_io_rPort_8_ofs_0 = x506_x313_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@21809.4]
  assign x257_lb_0_io_rPort_8_en_0 = _T_742 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@21811.4]
  assign x257_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21810.4]
  assign x257_lb_0_io_rPort_7_banks_1 = x500_x469_D23_number[2:0]; // @[MemInterfaceType.scala 106:58:@22000.4]
  assign x257_lb_0_io_rPort_7_banks_0 = x511_x474_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21999.4]
  assign x257_lb_0_io_rPort_7_ofs_0 = x329_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@22001.4]
  assign x257_lb_0_io_rPort_7_en_0 = _T_862 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@22003.4]
  assign x257_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@22002.4]
  assign x257_lb_0_io_rPort_6_banks_1 = x502_x472_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@22058.4]
  assign x257_lb_0_io_rPort_6_banks_0 = x511_x474_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@22057.4]
  assign x257_lb_0_io_rPort_6_ofs_0 = x334_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@22059.4]
  assign x257_lb_0_io_rPort_6_en_0 = _T_894 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@22061.4]
  assign x257_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@22060.4]
  assign x257_lb_0_io_rPort_5_banks_1 = x500_x469_D23_number[2:0]; // @[MemInterfaceType.scala 106:58:@21578.4]
  assign x257_lb_0_io_rPort_5_banks_0 = x492_x471_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21577.4]
  assign x257_lb_0_io_rPort_5_ofs_0 = x498_x295_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@21579.4]
  assign x257_lb_0_io_rPort_5_en_0 = _T_592 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@21581.4]
  assign x257_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21580.4]
  assign x257_lb_0_io_rPort_4_banks_1 = x500_x469_D23_number[2:0]; // @[MemInterfaceType.scala 106:58:@22279.4]
  assign x257_lb_0_io_rPort_4_banks_0 = x519_x475_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@22278.4]
  assign x257_lb_0_io_rPort_4_ofs_0 = x355_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@22280.4]
  assign x257_lb_0_io_rPort_4_en_0 = _T_1035 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@22282.4]
  assign x257_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@22281.4]
  assign x257_lb_0_io_rPort_3_banks_1 = x502_x472_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@22330.4]
  assign x257_lb_0_io_rPort_3_banks_0 = x519_x475_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@22329.4]
  assign x257_lb_0_io_rPort_3_ofs_0 = x360_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@22331.4]
  assign x257_lb_0_io_rPort_3_en_0 = _T_1066 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@22333.4]
  assign x257_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@22332.4]
  assign x257_lb_0_io_rPort_2_banks_1 = x507_x473_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@22379.4]
  assign x257_lb_0_io_rPort_2_banks_0 = x519_x475_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@22378.4]
  assign x257_lb_0_io_rPort_2_ofs_0 = x365_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@22380.4]
  assign x257_lb_0_io_rPort_2_en_0 = _T_1095 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@22382.4]
  assign x257_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@22381.4]
  assign x257_lb_0_io_rPort_1_banks_1 = x495_x470_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@21933.4]
  assign x257_lb_0_io_rPort_1_banks_0 = x511_x474_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21932.4]
  assign x257_lb_0_io_rPort_1_ofs_0 = x324_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@21934.4]
  assign x257_lb_0_io_rPort_1_en_0 = _T_827 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@21936.4]
  assign x257_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21935.4]
  assign x257_lb_0_io_rPort_0_banks_1 = x507_x473_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@22116.4]
  assign x257_lb_0_io_rPort_0_banks_0 = x511_x474_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@22115.4]
  assign x257_lb_0_io_rPort_0_ofs_0 = x339_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@22117.4]
  assign x257_lb_0_io_rPort_0_en_0 = _T_926 & x493_b256_D23; // @[MemInterfaceType.scala 110:79:@22119.4]
  assign x257_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@22118.4]
  assign x257_lb_0_io_wPort_1_banks_1 = x485_x470_D1_number[2:0]; // @[MemInterfaceType.scala 88:58:@21305.4]
  assign x257_lb_0_io_wPort_1_banks_0 = x477_x468_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@21304.4]
  assign x257_lb_0_io_wPort_1_ofs_0 = x278_sum_number[8:0]; // @[MemInterfaceType.scala 89:54:@21306.4]
  assign x257_lb_0_io_wPort_1_data_0 = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 90:56:@21307.4]
  assign x257_lb_0_io_wPort_1_en_0 = _T_437 & x478_b256_D2; // @[MemInterfaceType.scala 93:57:@21309.4]
  assign x257_lb_0_io_wPort_0_banks_1 = x482_x469_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@21211.4]
  assign x257_lb_0_io_wPort_0_banks_0 = x477_x468_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@21210.4]
  assign x257_lb_0_io_wPort_0_ofs_0 = x481_x272_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@21212.4]
  assign x257_lb_0_io_wPort_0_data_0 = RetimeWrapper_3_io_out; // @[MemInterfaceType.scala 90:56:@21213.4]
  assign x257_lb_0_io_wPort_0_en_0 = _T_381 & x478_b256_D2; // @[MemInterfaceType.scala 93:57:@21215.4]
  assign RetimeWrapper_clock = clock; // @[:@21019.4]
  assign RetimeWrapper_reset = reset; // @[:@21020.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21022.4]
  assign RetimeWrapper_io_in = io_in_x244_TDATA[15:0]; // @[package.scala 94:16:@21021.4]
  assign x272_sum_1_clock = clock; // @[:@21131.4]
  assign x272_sum_1_reset = reset; // @[:@21132.4]
  assign x272_sum_1_io_a = _T_337[31:0]; // @[Math.scala 151:17:@21133.4]
  assign x272_sum_1_io_b = {_T_345,_T_346}; // @[Math.scala 152:17:@21134.4]
  assign x272_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21135.4]
  assign RetimeWrapper_1_clock = clock; // @[:@21141.4]
  assign RetimeWrapper_1_reset = reset; // @[:@21142.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21144.4]
  assign RetimeWrapper_1_io_in = $unsigned(_T_310); // @[package.scala 94:16:@21143.4]
  assign RetimeWrapper_2_clock = clock; // @[:@21150.4]
  assign RetimeWrapper_2_reset = reset; // @[:@21151.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21153.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@21152.4]
  assign RetimeWrapper_3_clock = clock; // @[:@21159.4]
  assign RetimeWrapper_3_reset = reset; // @[:@21160.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21162.4]
  assign RetimeWrapper_3_io_in = x476_x258_D1_0_number[7:0]; // @[package.scala 94:16:@21161.4]
  assign RetimeWrapper_4_clock = clock; // @[:@21168.4]
  assign RetimeWrapper_4_reset = reset; // @[:@21169.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21171.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@21170.4]
  assign RetimeWrapper_5_clock = clock; // @[:@21177.4]
  assign RetimeWrapper_5_reset = reset; // @[:@21178.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21180.4]
  assign RetimeWrapper_5_io_in = x272_sum_1_io_result; // @[package.scala 94:16:@21179.4]
  assign RetimeWrapper_6_clock = clock; // @[:@21186.4]
  assign RetimeWrapper_6_reset = reset; // @[:@21187.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21189.4]
  assign RetimeWrapper_6_io_in = $unsigned(_T_322); // @[package.scala 94:16:@21188.4]
  assign RetimeWrapper_7_clock = clock; // @[:@21197.4]
  assign RetimeWrapper_7_reset = reset; // @[:@21198.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21200.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21199.4]
  assign x274_rdcol_1_clock = clock; // @[:@21220.4]
  assign x274_rdcol_1_reset = reset; // @[:@21221.4]
  assign x274_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@21222.4]
  assign x274_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@21223.4]
  assign x274_rdcol_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21224.4]
  assign RetimeWrapper_8_clock = clock; // @[:@21252.4]
  assign RetimeWrapper_8_reset = reset; // @[:@21253.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21255.4]
  assign RetimeWrapper_8_io_in = _T_337[31:0]; // @[package.scala 94:16:@21254.4]
  assign x278_sum_1_clock = clock; // @[:@21261.4]
  assign x278_sum_1_reset = reset; // @[:@21262.4]
  assign x278_sum_1_io_a = RetimeWrapper_8_io_out; // @[Math.scala 151:17:@21263.4]
  assign x278_sum_1_io_b = {_T_410,_T_411}; // @[Math.scala 152:17:@21264.4]
  assign x278_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21265.4]
  assign RetimeWrapper_9_clock = clock; // @[:@21271.4]
  assign RetimeWrapper_9_reset = reset; // @[:@21272.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21274.4]
  assign RetimeWrapper_9_io_in = x476_x258_D1_0_number[15:8]; // @[package.scala 94:16:@21273.4]
  assign RetimeWrapper_10_clock = clock; // @[:@21280.4]
  assign RetimeWrapper_10_reset = reset; // @[:@21281.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21283.4]
  assign RetimeWrapper_10_io_in = $unsigned(_T_401); // @[package.scala 94:16:@21282.4]
  assign RetimeWrapper_11_clock = clock; // @[:@21291.4]
  assign RetimeWrapper_11_reset = reset; // @[:@21292.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21294.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21293.4]
  assign RetimeWrapper_12_clock = clock; // @[:@21312.4]
  assign RetimeWrapper_12_reset = reset; // @[:@21313.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21315.4]
  assign RetimeWrapper_12_io_in = __io_result; // @[package.scala 94:16:@21314.4]
  assign x281_1_clock = clock; // @[:@21323.4]
  assign x281_1_reset = reset; // @[:@21324.4]
  assign x281_1_io_a = RetimeWrapper_12_io_out; // @[Math.scala 367:17:@21325.4]
  assign x281_1_io_flow = io_in_x245_TREADY; // @[Math.scala 369:20:@21327.4]
  assign RetimeWrapper_13_clock = clock; // @[:@21340.4]
  assign RetimeWrapper_13_reset = reset; // @[:@21341.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21343.4]
  assign RetimeWrapper_13_io_in = x274_rdcol_1_io_result; // @[package.scala 94:16:@21342.4]
  assign RetimeWrapper_14_clock = clock; // @[:@21356.4]
  assign RetimeWrapper_14_reset = reset; // @[:@21357.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21359.4]
  assign RetimeWrapper_14_io_in = $signed(_T_454) < $signed(32'sh0); // @[package.scala 94:16:@21358.4]
  assign RetimeWrapper_15_clock = clock; // @[:@21396.4]
  assign RetimeWrapper_15_reset = reset; // @[:@21397.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21399.4]
  assign RetimeWrapper_15_io_in = {_T_410,_T_411}; // @[package.scala 94:16:@21398.4]
  assign x289_sum_1_clock = clock; // @[:@21405.4]
  assign x289_sum_1_reset = reset; // @[:@21406.4]
  assign x289_sum_1_io_a = _T_500[31:0]; // @[Math.scala 151:17:@21407.4]
  assign x289_sum_1_io_b = RetimeWrapper_15_io_out; // @[Math.scala 152:17:@21408.4]
  assign x289_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21409.4]
  assign RetimeWrapper_16_clock = clock; // @[:@21415.4]
  assign RetimeWrapper_16_reset = reset; // @[:@21416.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21418.4]
  assign RetimeWrapper_16_io_in = x289_sum_1_io_result; // @[package.scala 94:16:@21417.4]
  assign RetimeWrapper_17_clock = clock; // @[:@21424.4]
  assign RetimeWrapper_17_reset = reset; // @[:@21425.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21427.4]
  assign RetimeWrapper_17_io_in = ~ x284; // @[package.scala 94:16:@21426.4]
  assign RetimeWrapper_18_clock = clock; // @[:@21433.4]
  assign RetimeWrapper_18_reset = reset; // @[:@21434.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21436.4]
  assign RetimeWrapper_18_io_in = $unsigned(_T_485); // @[package.scala 94:16:@21435.4]
  assign RetimeWrapper_19_clock = clock; // @[:@21442.4]
  assign RetimeWrapper_19_reset = reset; // @[:@21443.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21445.4]
  assign RetimeWrapper_19_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@21444.4]
  assign RetimeWrapper_20_clock = clock; // @[:@21451.4]
  assign RetimeWrapper_20_reset = reset; // @[:@21452.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21454.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@21453.4]
  assign RetimeWrapper_21_clock = clock; // @[:@21460.4]
  assign RetimeWrapper_21_reset = reset; // @[:@21461.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21463.4]
  assign RetimeWrapper_21_io_in = $unsigned(_T_401); // @[package.scala 94:16:@21462.4]
  assign RetimeWrapper_22_clock = clock; // @[:@21472.4]
  assign RetimeWrapper_22_reset = reset; // @[:@21473.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21475.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21474.4]
  assign RetimeWrapper_23_clock = clock; // @[:@21493.4]
  assign RetimeWrapper_23_reset = reset; // @[:@21494.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21496.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@21495.4]
  assign RetimeWrapper_24_clock = clock; // @[:@21517.4]
  assign RetimeWrapper_24_reset = reset; // @[:@21518.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21520.4]
  assign RetimeWrapper_24_io_in = {_T_345,_T_346}; // @[package.scala 94:16:@21519.4]
  assign x295_sum_1_clock = clock; // @[:@21526.4]
  assign x295_sum_1_reset = reset; // @[:@21527.4]
  assign x295_sum_1_io_a = _T_500[31:0]; // @[Math.scala 151:17:@21528.4]
  assign x295_sum_1_io_b = RetimeWrapper_24_io_out; // @[Math.scala 152:17:@21529.4]
  assign x295_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21530.4]
  assign RetimeWrapper_25_clock = clock; // @[:@21536.4]
  assign RetimeWrapper_25_reset = reset; // @[:@21537.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21539.4]
  assign RetimeWrapper_25_io_in = x295_sum_1_io_result; // @[package.scala 94:16:@21538.4]
  assign RetimeWrapper_26_clock = clock; // @[:@21545.4]
  assign RetimeWrapper_26_reset = reset; // @[:@21546.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21548.4]
  assign RetimeWrapper_26_io_in = ~ x293; // @[package.scala 94:16:@21547.4]
  assign RetimeWrapper_27_clock = clock; // @[:@21554.4]
  assign RetimeWrapper_27_reset = reset; // @[:@21555.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21557.4]
  assign RetimeWrapper_27_io_in = $unsigned(_T_322); // @[package.scala 94:16:@21556.4]
  assign RetimeWrapper_28_clock = clock; // @[:@21566.4]
  assign RetimeWrapper_28_reset = reset; // @[:@21567.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21569.4]
  assign RetimeWrapper_28_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21568.4]
  assign x298_rdcol_1_clock = clock; // @[:@21589.4]
  assign x298_rdcol_1_reset = reset; // @[:@21590.4]
  assign x298_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@21591.4]
  assign x298_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@21592.4]
  assign x298_rdcol_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21593.4]
  assign RetimeWrapper_29_clock = clock; // @[:@21632.4]
  assign RetimeWrapper_29_reset = reset; // @[:@21633.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21635.4]
  assign RetimeWrapper_29_io_in = {_T_633,_T_634}; // @[package.scala 94:16:@21634.4]
  assign x304_sum_1_clock = clock; // @[:@21641.4]
  assign x304_sum_1_reset = reset; // @[:@21642.4]
  assign x304_sum_1_io_a = _T_500[31:0]; // @[Math.scala 151:17:@21643.4]
  assign x304_sum_1_io_b = RetimeWrapper_29_io_out; // @[Math.scala 152:17:@21644.4]
  assign x304_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21645.4]
  assign RetimeWrapper_30_clock = clock; // @[:@21651.4]
  assign RetimeWrapper_30_reset = reset; // @[:@21652.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21654.4]
  assign RetimeWrapper_30_io_in = $unsigned(_T_624); // @[package.scala 94:16:@21653.4]
  assign RetimeWrapper_31_clock = clock; // @[:@21660.4]
  assign RetimeWrapper_31_reset = reset; // @[:@21661.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21663.4]
  assign RetimeWrapper_31_io_in = ~ x300; // @[package.scala 94:16:@21662.4]
  assign RetimeWrapper_32_clock = clock; // @[:@21669.4]
  assign RetimeWrapper_32_reset = reset; // @[:@21670.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21672.4]
  assign RetimeWrapper_32_io_in = x304_sum_1_io_result; // @[package.scala 94:16:@21671.4]
  assign RetimeWrapper_33_clock = clock; // @[:@21681.4]
  assign RetimeWrapper_33_reset = reset; // @[:@21682.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21684.4]
  assign RetimeWrapper_33_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21683.4]
  assign x307_rdcol_1_clock = clock; // @[:@21704.4]
  assign x307_rdcol_1_reset = reset; // @[:@21705.4]
  assign x307_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@21706.4]
  assign x307_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@21707.4]
  assign x307_rdcol_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21708.4]
  assign RetimeWrapper_34_clock = clock; // @[:@21747.4]
  assign RetimeWrapper_34_reset = reset; // @[:@21748.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21750.4]
  assign RetimeWrapper_34_io_in = {_T_708,_T_709}; // @[package.scala 94:16:@21749.4]
  assign x313_sum_1_clock = clock; // @[:@21756.4]
  assign x313_sum_1_reset = reset; // @[:@21757.4]
  assign x313_sum_1_io_a = _T_500[31:0]; // @[Math.scala 151:17:@21758.4]
  assign x313_sum_1_io_b = RetimeWrapper_34_io_out; // @[Math.scala 152:17:@21759.4]
  assign x313_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21760.4]
  assign RetimeWrapper_35_clock = clock; // @[:@21766.4]
  assign RetimeWrapper_35_reset = reset; // @[:@21767.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21769.4]
  assign RetimeWrapper_35_io_in = x313_sum_1_io_result; // @[package.scala 94:16:@21768.4]
  assign RetimeWrapper_36_clock = clock; // @[:@21775.4]
  assign RetimeWrapper_36_reset = reset; // @[:@21776.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21778.4]
  assign RetimeWrapper_36_io_in = $unsigned(_T_699); // @[package.scala 94:16:@21777.4]
  assign RetimeWrapper_37_clock = clock; // @[:@21784.4]
  assign RetimeWrapper_37_reset = reset; // @[:@21785.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21787.4]
  assign RetimeWrapper_37_io_in = ~ x309; // @[package.scala 94:16:@21786.4]
  assign RetimeWrapper_38_clock = clock; // @[:@21796.4]
  assign RetimeWrapper_38_reset = reset; // @[:@21797.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21799.4]
  assign RetimeWrapper_38_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21798.4]
  assign x316_rdrow_1_clock = clock; // @[:@21819.4]
  assign x316_rdrow_1_reset = reset; // @[:@21820.4]
  assign x316_rdrow_1_io_a = RetimeWrapper_12_io_out; // @[Math.scala 192:17:@21821.4]
  assign x316_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@21822.4]
  assign x316_rdrow_1_io_flow = io_in_x245_TREADY; // @[Math.scala 194:20:@21823.4]
  assign x317_1_clock = clock; // @[:@21831.4]
  assign x317_1_reset = reset; // @[:@21832.4]
  assign x317_1_io_a = x316_rdrow_1_io_result; // @[Math.scala 367:17:@21833.4]
  assign x317_1_io_flow = io_in_x245_TREADY; // @[Math.scala 369:20:@21835.4]
  assign RetimeWrapper_39_clock = clock; // @[:@21881.4]
  assign RetimeWrapper_39_reset = reset; // @[:@21882.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21884.4]
  assign RetimeWrapper_39_io_in = {_T_410,_T_411}; // @[package.scala 94:16:@21883.4]
  assign x324_sum_1_clock = clock; // @[:@21890.4]
  assign x324_sum_1_reset = reset; // @[:@21891.4]
  assign x324_sum_1_io_a = _T_798[31:0]; // @[Math.scala 151:17:@21892.4]
  assign x324_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@21893.4]
  assign x324_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21894.4]
  assign RetimeWrapper_40_clock = clock; // @[:@21900.4]
  assign RetimeWrapper_40_reset = reset; // @[:@21901.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21903.4]
  assign RetimeWrapper_40_io_in = ~ x319; // @[package.scala 94:16:@21902.4]
  assign RetimeWrapper_41_clock = clock; // @[:@21909.4]
  assign RetimeWrapper_41_reset = reset; // @[:@21910.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21912.4]
  assign RetimeWrapper_41_io_in = $unsigned(_T_781); // @[package.scala 94:16:@21911.4]
  assign RetimeWrapper_42_clock = clock; // @[:@21921.4]
  assign RetimeWrapper_42_reset = reset; // @[:@21922.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21924.4]
  assign RetimeWrapper_42_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21923.4]
  assign RetimeWrapper_43_clock = clock; // @[:@21942.4]
  assign RetimeWrapper_43_reset = reset; // @[:@21943.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21945.4]
  assign RetimeWrapper_43_io_in = $signed(_T_554) < $signed(32'sh0); // @[package.scala 94:16:@21944.4]
  assign RetimeWrapper_44_clock = clock; // @[:@21957.4]
  assign RetimeWrapper_44_reset = reset; // @[:@21958.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21960.4]
  assign RetimeWrapper_44_io_in = {_T_345,_T_346}; // @[package.scala 94:16:@21959.4]
  assign x329_sum_1_clock = clock; // @[:@21966.4]
  assign x329_sum_1_reset = reset; // @[:@21967.4]
  assign x329_sum_1_io_a = _T_798[31:0]; // @[Math.scala 151:17:@21968.4]
  assign x329_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@21969.4]
  assign x329_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@21970.4]
  assign RetimeWrapper_45_clock = clock; // @[:@21976.4]
  assign RetimeWrapper_45_reset = reset; // @[:@21977.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21979.4]
  assign RetimeWrapper_45_io_in = ~ x327; // @[package.scala 94:16:@21978.4]
  assign RetimeWrapper_46_clock = clock; // @[:@21988.4]
  assign RetimeWrapper_46_reset = reset; // @[:@21989.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21991.4]
  assign RetimeWrapper_46_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21990.4]
  assign RetimeWrapper_47_clock = clock; // @[:@22015.4]
  assign RetimeWrapper_47_reset = reset; // @[:@22016.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22018.4]
  assign RetimeWrapper_47_io_in = {_T_633,_T_634}; // @[package.scala 94:16:@22017.4]
  assign x334_sum_1_clock = clock; // @[:@22024.4]
  assign x334_sum_1_reset = reset; // @[:@22025.4]
  assign x334_sum_1_io_a = _T_798[31:0]; // @[Math.scala 151:17:@22026.4]
  assign x334_sum_1_io_b = RetimeWrapper_47_io_out; // @[Math.scala 152:17:@22027.4]
  assign x334_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22028.4]
  assign RetimeWrapper_48_clock = clock; // @[:@22034.4]
  assign RetimeWrapper_48_reset = reset; // @[:@22035.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22037.4]
  assign RetimeWrapper_48_io_in = ~ x332; // @[package.scala 94:16:@22036.4]
  assign RetimeWrapper_49_clock = clock; // @[:@22046.4]
  assign RetimeWrapper_49_reset = reset; // @[:@22047.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22049.4]
  assign RetimeWrapper_49_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22048.4]
  assign RetimeWrapper_50_clock = clock; // @[:@22073.4]
  assign RetimeWrapper_50_reset = reset; // @[:@22074.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22076.4]
  assign RetimeWrapper_50_io_in = {_T_708,_T_709}; // @[package.scala 94:16:@22075.4]
  assign x339_sum_1_clock = clock; // @[:@22082.4]
  assign x339_sum_1_reset = reset; // @[:@22083.4]
  assign x339_sum_1_io_a = _T_798[31:0]; // @[Math.scala 151:17:@22084.4]
  assign x339_sum_1_io_b = RetimeWrapper_50_io_out; // @[Math.scala 152:17:@22085.4]
  assign x339_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22086.4]
  assign RetimeWrapper_51_clock = clock; // @[:@22092.4]
  assign RetimeWrapper_51_reset = reset; // @[:@22093.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22095.4]
  assign RetimeWrapper_51_io_in = ~ x337; // @[package.scala 94:16:@22094.4]
  assign RetimeWrapper_52_clock = clock; // @[:@22104.4]
  assign RetimeWrapper_52_reset = reset; // @[:@22105.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22107.4]
  assign RetimeWrapper_52_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22106.4]
  assign x342_rdrow_1_clock = clock; // @[:@22127.4]
  assign x342_rdrow_1_reset = reset; // @[:@22128.4]
  assign x342_rdrow_1_io_a = RetimeWrapper_12_io_out; // @[Math.scala 192:17:@22129.4]
  assign x342_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@22130.4]
  assign x342_rdrow_1_io_flow = io_in_x245_TREADY; // @[Math.scala 194:20:@22131.4]
  assign x343_1_clock = clock; // @[:@22139.4]
  assign x343_1_reset = reset; // @[:@22140.4]
  assign x343_1_io_a = x342_rdrow_1_io_result; // @[Math.scala 367:17:@22141.4]
  assign x343_1_io_flow = io_in_x245_TREADY; // @[Math.scala 369:20:@22143.4]
  assign x350_sum_1_clock = clock; // @[:@22187.4]
  assign x350_sum_1_reset = reset; // @[:@22188.4]
  assign x350_sum_1_io_a = _T_980[31:0]; // @[Math.scala 151:17:@22189.4]
  assign x350_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@22190.4]
  assign x350_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22191.4]
  assign RetimeWrapper_53_clock = clock; // @[:@22197.4]
  assign RetimeWrapper_53_reset = reset; // @[:@22198.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22200.4]
  assign RetimeWrapper_53_io_in = $unsigned(_T_965); // @[package.scala 94:16:@22199.4]
  assign RetimeWrapper_54_clock = clock; // @[:@22206.4]
  assign RetimeWrapper_54_reset = reset; // @[:@22207.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22209.4]
  assign RetimeWrapper_54_io_in = ~ x345; // @[package.scala 94:16:@22208.4]
  assign RetimeWrapper_55_clock = clock; // @[:@22218.4]
  assign RetimeWrapper_55_reset = reset; // @[:@22219.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22221.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22220.4]
  assign x355_sum_1_clock = clock; // @[:@22245.4]
  assign x355_sum_1_reset = reset; // @[:@22246.4]
  assign x355_sum_1_io_a = _T_980[31:0]; // @[Math.scala 151:17:@22247.4]
  assign x355_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@22248.4]
  assign x355_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22249.4]
  assign RetimeWrapper_56_clock = clock; // @[:@22255.4]
  assign RetimeWrapper_56_reset = reset; // @[:@22256.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22258.4]
  assign RetimeWrapper_56_io_in = ~ x353; // @[package.scala 94:16:@22257.4]
  assign RetimeWrapper_57_clock = clock; // @[:@22267.4]
  assign RetimeWrapper_57_reset = reset; // @[:@22268.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22270.4]
  assign RetimeWrapper_57_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22269.4]
  assign x360_sum_1_clock = clock; // @[:@22296.4]
  assign x360_sum_1_reset = reset; // @[:@22297.4]
  assign x360_sum_1_io_a = _T_980[31:0]; // @[Math.scala 151:17:@22298.4]
  assign x360_sum_1_io_b = RetimeWrapper_47_io_out; // @[Math.scala 152:17:@22299.4]
  assign x360_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22300.4]
  assign RetimeWrapper_58_clock = clock; // @[:@22306.4]
  assign RetimeWrapper_58_reset = reset; // @[:@22307.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22309.4]
  assign RetimeWrapper_58_io_in = ~ x358; // @[package.scala 94:16:@22308.4]
  assign RetimeWrapper_59_clock = clock; // @[:@22318.4]
  assign RetimeWrapper_59_reset = reset; // @[:@22319.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22321.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22320.4]
  assign x365_sum_1_clock = clock; // @[:@22345.4]
  assign x365_sum_1_reset = reset; // @[:@22346.4]
  assign x365_sum_1_io_a = _T_980[31:0]; // @[Math.scala 151:17:@22347.4]
  assign x365_sum_1_io_b = RetimeWrapper_50_io_out; // @[Math.scala 152:17:@22348.4]
  assign x365_sum_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22349.4]
  assign RetimeWrapper_60_clock = clock; // @[:@22355.4]
  assign RetimeWrapper_60_reset = reset; // @[:@22356.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22358.4]
  assign RetimeWrapper_60_io_in = ~ x363; // @[package.scala 94:16:@22357.4]
  assign RetimeWrapper_61_clock = clock; // @[:@22367.4]
  assign RetimeWrapper_61_reset = reset; // @[:@22368.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22370.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22369.4]
  assign RetimeWrapper_62_clock = clock; // @[:@22413.4]
  assign RetimeWrapper_62_reset = reset; // @[:@22414.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22416.4]
  assign RetimeWrapper_62_io_in = _T_1101[7:0]; // @[package.scala 94:16:@22415.4]
  assign RetimeWrapper_63_clock = clock; // @[:@22422.4]
  assign RetimeWrapper_63_reset = reset; // @[:@22423.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22425.4]
  assign RetimeWrapper_63_io_in = x257_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@22424.4]
  assign x373_x11_1_clock = clock; // @[:@22431.4]
  assign x373_x11_1_reset = reset; // @[:@22432.4]
  assign x373_x11_1_io_a = RetimeWrapper_63_io_out; // @[Math.scala 151:17:@22433.4]
  assign x373_x11_1_io_b = RetimeWrapper_62_io_out; // @[Math.scala 152:17:@22434.4]
  assign x373_x11_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22435.4]
  assign RetimeWrapper_64_clock = clock; // @[:@22441.4]
  assign RetimeWrapper_64_reset = reset; // @[:@22442.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22444.4]
  assign RetimeWrapper_64_io_in = _T_1105[7:0]; // @[package.scala 94:16:@22443.4]
  assign RetimeWrapper_65_clock = clock; // @[:@22450.4]
  assign RetimeWrapper_65_reset = reset; // @[:@22451.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22453.4]
  assign RetimeWrapper_65_io_in = x257_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@22452.4]
  assign x374_x12_1_clock = clock; // @[:@22459.4]
  assign x374_x12_1_reset = reset; // @[:@22460.4]
  assign x374_x12_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@22461.4]
  assign x374_x12_1_io_b = RetimeWrapper_64_io_out; // @[Math.scala 152:17:@22462.4]
  assign x374_x12_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22463.4]
  assign x375_x11_1_clock = clock; // @[:@22469.4]
  assign x375_x11_1_reset = reset; // @[:@22470.4]
  assign x375_x11_1_io_a = _T_1109[7:0]; // @[Math.scala 151:17:@22471.4]
  assign x375_x11_1_io_b = _T_1113[7:0]; // @[Math.scala 152:17:@22472.4]
  assign x375_x11_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22473.4]
  assign x376_x12_1_clock = clock; // @[:@22479.4]
  assign x376_x12_1_reset = reset; // @[:@22480.4]
  assign x376_x12_1_io_a = x257_lb_0_io_rPort_9_output_0; // @[Math.scala 151:17:@22481.4]
  assign x376_x12_1_io_b = _T_1117[7:0]; // @[Math.scala 152:17:@22482.4]
  assign x376_x12_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22483.4]
  assign RetimeWrapper_66_clock = clock; // @[:@22489.4]
  assign RetimeWrapper_66_reset = reset; // @[:@22490.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22492.4]
  assign RetimeWrapper_66_io_in = x373_x11_1_io_result; // @[package.scala 94:16:@22491.4]
  assign RetimeWrapper_67_clock = clock; // @[:@22498.4]
  assign RetimeWrapper_67_reset = reset; // @[:@22499.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22501.4]
  assign RetimeWrapper_67_io_in = x374_x12_1_io_result; // @[package.scala 94:16:@22500.4]
  assign x377_x11_1_io_a = RetimeWrapper_66_io_out; // @[Math.scala 151:17:@22509.4]
  assign x377_x11_1_io_b = RetimeWrapper_67_io_out; // @[Math.scala 152:17:@22510.4]
  assign x378_x12_1_io_a = x375_x11_1_io_result; // @[Math.scala 151:17:@22519.4]
  assign x378_x12_1_io_b = x376_x12_1_io_result; // @[Math.scala 152:17:@22520.4]
  assign RetimeWrapper_68_clock = clock; // @[:@22527.4]
  assign RetimeWrapper_68_reset = reset; // @[:@22528.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22530.4]
  assign RetimeWrapper_68_io_in = x378_x12_1_io_result; // @[package.scala 94:16:@22529.4]
  assign x379_x11_1_io_a = x377_x11_1_io_result; // @[Math.scala 151:17:@22538.4]
  assign x379_x11_1_io_b = RetimeWrapper_68_io_out; // @[Math.scala 152:17:@22539.4]
  assign RetimeWrapper_69_clock = clock; // @[:@22546.4]
  assign RetimeWrapper_69_reset = reset; // @[:@22547.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22549.4]
  assign RetimeWrapper_69_io_in = x257_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@22548.4]
  assign x380_sum_1_io_a = x379_x11_1_io_result; // @[Math.scala 151:17:@22557.4]
  assign x380_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@22558.4]
  assign RetimeWrapper_70_clock = clock; // @[:@22569.4]
  assign RetimeWrapper_70_reset = reset; // @[:@22570.4]
  assign RetimeWrapper_70_io_flow = io_in_x245_TREADY; // @[package.scala 95:18:@22572.4]
  assign RetimeWrapper_70_io_in = {4'h0,_T_1174}; // @[package.scala 94:16:@22571.4]
  assign RetimeWrapper_71_clock = clock; // @[:@22604.4]
  assign RetimeWrapper_71_reset = reset; // @[:@22605.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22607.4]
  assign RetimeWrapper_71_io_in = _T_1181[7:0]; // @[package.scala 94:16:@22606.4]
  assign RetimeWrapper_72_clock = clock; // @[:@22613.4]
  assign RetimeWrapper_72_reset = reset; // @[:@22614.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22616.4]
  assign RetimeWrapper_72_io_in = x257_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@22615.4]
  assign x387_x11_1_clock = clock; // @[:@22622.4]
  assign x387_x11_1_reset = reset; // @[:@22623.4]
  assign x387_x11_1_io_a = RetimeWrapper_72_io_out; // @[Math.scala 151:17:@22624.4]
  assign x387_x11_1_io_b = RetimeWrapper_71_io_out; // @[Math.scala 152:17:@22625.4]
  assign x387_x11_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22626.4]
  assign RetimeWrapper_73_clock = clock; // @[:@22632.4]
  assign RetimeWrapper_73_reset = reset; // @[:@22633.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22635.4]
  assign RetimeWrapper_73_io_in = x257_lb_0_io_rPort_8_output_0; // @[package.scala 94:16:@22634.4]
  assign RetimeWrapper_74_clock = clock; // @[:@22641.4]
  assign RetimeWrapper_74_reset = reset; // @[:@22642.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22644.4]
  assign RetimeWrapper_74_io_in = _T_1185[7:0]; // @[package.scala 94:16:@22643.4]
  assign x388_x12_1_clock = clock; // @[:@22650.4]
  assign x388_x12_1_reset = reset; // @[:@22651.4]
  assign x388_x12_1_io_a = RetimeWrapper_73_io_out; // @[Math.scala 151:17:@22652.4]
  assign x388_x12_1_io_b = RetimeWrapper_74_io_out; // @[Math.scala 152:17:@22653.4]
  assign x388_x12_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22654.4]
  assign x389_x11_1_clock = clock; // @[:@22660.4]
  assign x389_x11_1_reset = reset; // @[:@22661.4]
  assign x389_x11_1_io_a = _T_1189[7:0]; // @[Math.scala 151:17:@22662.4]
  assign x389_x11_1_io_b = _T_1193[7:0]; // @[Math.scala 152:17:@22663.4]
  assign x389_x11_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22664.4]
  assign x390_x12_1_clock = clock; // @[:@22670.4]
  assign x390_x12_1_reset = reset; // @[:@22671.4]
  assign x390_x12_1_io_a = x257_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@22672.4]
  assign x390_x12_1_io_b = _T_1197[7:0]; // @[Math.scala 152:17:@22673.4]
  assign x390_x12_1_io_flow = io_in_x245_TREADY; // @[Math.scala 153:20:@22674.4]
  assign RetimeWrapper_75_clock = clock; // @[:@22680.4]
  assign RetimeWrapper_75_reset = reset; // @[:@22681.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22683.4]
  assign RetimeWrapper_75_io_in = x387_x11_1_io_result; // @[package.scala 94:16:@22682.4]
  assign RetimeWrapper_76_clock = clock; // @[:@22689.4]
  assign RetimeWrapper_76_reset = reset; // @[:@22690.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22692.4]
  assign RetimeWrapper_76_io_in = x388_x12_1_io_result; // @[package.scala 94:16:@22691.4]
  assign x391_x11_1_io_a = RetimeWrapper_75_io_out; // @[Math.scala 151:17:@22702.4]
  assign x391_x11_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@22703.4]
  assign x392_x12_1_io_a = x389_x11_1_io_result; // @[Math.scala 151:17:@22712.4]
  assign x392_x12_1_io_b = x390_x12_1_io_result; // @[Math.scala 152:17:@22713.4]
  assign RetimeWrapper_77_clock = clock; // @[:@22720.4]
  assign RetimeWrapper_77_reset = reset; // @[:@22721.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22723.4]
  assign RetimeWrapper_77_io_in = x392_x12_1_io_result; // @[package.scala 94:16:@22722.4]
  assign x393_x11_1_io_a = x391_x11_1_io_result; // @[Math.scala 151:17:@22731.4]
  assign x393_x11_1_io_b = RetimeWrapper_77_io_out; // @[Math.scala 152:17:@22732.4]
  assign RetimeWrapper_78_clock = clock; // @[:@22739.4]
  assign RetimeWrapper_78_reset = reset; // @[:@22740.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22742.4]
  assign RetimeWrapper_78_io_in = x257_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@22741.4]
  assign x394_sum_1_io_a = x393_x11_1_io_result; // @[Math.scala 151:17:@22750.4]
  assign x394_sum_1_io_b = RetimeWrapper_78_io_out; // @[Math.scala 152:17:@22751.4]
  assign RetimeWrapper_79_clock = clock; // @[:@22762.4]
  assign RetimeWrapper_79_reset = reset; // @[:@22763.4]
  assign RetimeWrapper_79_io_flow = io_in_x245_TREADY; // @[package.scala 95:18:@22765.4]
  assign RetimeWrapper_79_io_in = {4'h0,_T_1256}; // @[package.scala 94:16:@22764.4]
  assign RetimeWrapper_80_clock = clock; // @[:@22772.4]
  assign RetimeWrapper_80_reset = reset; // @[:@22773.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22775.4]
  assign RetimeWrapper_80_io_in = RetimeWrapper_79_io_out; // @[package.scala 94:16:@22774.4]
  assign RetimeWrapper_81_clock = clock; // @[:@22781.4]
  assign RetimeWrapper_81_reset = reset; // @[:@22782.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22784.4]
  assign RetimeWrapper_81_io_in = RetimeWrapper_70_io_out; // @[package.scala 94:16:@22783.4]
  assign RetimeWrapper_82_clock = clock; // @[:@22796.4]
  assign RetimeWrapper_82_reset = reset; // @[:@22797.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22799.4]
  assign RetimeWrapper_82_io_in = {x541_x381_D1_number,x540_x395_D1_number}; // @[package.scala 94:16:@22798.4]
  assign RetimeWrapper_83_clock = clock; // @[:@22805.4]
  assign RetimeWrapper_83_reset = reset; // @[:@22806.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22808.4]
  assign RetimeWrapper_83_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@22807.4]
  assign RetimeWrapper_84_clock = clock; // @[:@22814.4]
  assign RetimeWrapper_84_reset = reset; // @[:@22815.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22817.4]
  assign RetimeWrapper_84_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@22816.4]
  assign RetimeWrapper_85_clock = clock; // @[:@22823.4]
  assign RetimeWrapper_85_reset = reset; // @[:@22824.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22826.4]
  assign RetimeWrapper_85_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22825.4]
endmodule
module x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1( // @[:@22844.2]
  input          clock, // @[:@22845.4]
  input          reset, // @[:@22846.4]
  input          io_in_x244_TVALID, // @[:@22847.4]
  output         io_in_x244_TREADY, // @[:@22847.4]
  input  [255:0] io_in_x244_TDATA, // @[:@22847.4]
  input  [7:0]   io_in_x244_TID, // @[:@22847.4]
  input  [7:0]   io_in_x244_TDEST, // @[:@22847.4]
  output         io_in_x245_TVALID, // @[:@22847.4]
  input          io_in_x245_TREADY, // @[:@22847.4]
  output [255:0] io_in_x245_TDATA, // @[:@22847.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@22847.4]
  input          io_sigsIn_smChildAcks_0, // @[:@22847.4]
  output         io_sigsOut_smDoneIn_0, // @[:@22847.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@22847.4]
  input          io_rr // @[:@22847.4]
);
  wire  x252_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire  x252_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire  x252_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire  x252_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire [31:0] x252_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire [31:0] x252_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire  x252_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire  x252_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire  x252_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@22857.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@22987.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@22987.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@22987.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@22987.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@22987.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@22995.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@22995.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@22995.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@22995.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@22995.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TREADY; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire [255:0] x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TDATA; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire [7:0] x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TID; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire [7:0] x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TDEST; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TVALID; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TREADY; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire [255:0] x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TDATA; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire [31:0] x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire [31:0] x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
  wire  _T_239; // @[package.scala 96:25:@22950.4 package.scala 96:25:@22951.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x401_outr_UnitPipe.scala 68:66:@22956.4]
  wire  _T_252; // @[package.scala 96:25:@22992.4 package.scala 96:25:@22993.4]
  wire  _T_258; // @[package.scala 96:25:@23000.4 package.scala 96:25:@23001.4]
  wire  _T_261; // @[SpatialBlocks.scala 138:93:@23003.4]
  wire  x400_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@23004.4]
  wire  _T_263; // @[SpatialBlocks.scala 157:36:@23012.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:78:@23013.4]
  wire  _T_271; // @[SpatialBlocks.scala 159:58:@23025.4]
  x252_ctrchain x252_ctrchain ( // @[SpatialBlocks.scala 37:22:@22857.4]
    .clock(x252_ctrchain_clock),
    .reset(x252_ctrchain_reset),
    .io_input_reset(x252_ctrchain_io_input_reset),
    .io_input_enable(x252_ctrchain_io_input_enable),
    .io_output_counts_1(x252_ctrchain_io_output_counts_1),
    .io_output_counts_0(x252_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x252_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x252_ctrchain_io_output_oobs_1),
    .io_output_done(x252_ctrchain_io_output_done)
  );
  x400_inr_Foreach_SAMPLER_BOX_sm x400_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 32:18:@22917.4]
    .clock(x400_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x400_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x400_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x400_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x400_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x400_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x400_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x400_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x400_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@22945.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@22987.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@22995.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1 x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 574:24:@23030.4]
    .clock(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x244_TREADY(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TREADY),
    .io_in_x244_TDATA(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TDATA),
    .io_in_x244_TID(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TID),
    .io_in_x244_TDEST(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TDEST),
    .io_in_x245_TVALID(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TVALID),
    .io_in_x245_TREADY(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TREADY),
    .io_in_x245_TDATA(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TDATA),
    .io_sigsIn_backpressure(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@22950.4 package.scala 96:25:@22951.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x244_TVALID | x400_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x401_outr_UnitPipe.scala 68:66:@22956.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@22992.4 package.scala 96:25:@22993.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@23000.4 package.scala 96:25:@23001.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 138:93:@23003.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 138:90:@23004.4]
  assign _T_263 = x400_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@23012.4]
  assign _T_264 = ~ x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@23013.4]
  assign _T_271 = x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@23025.4]
  assign io_in_x244_TREADY = x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TREADY; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 48:23:@23088.4]
  assign io_in_x245_TVALID = x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TVALID; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 49:23:@23098.4]
  assign io_in_x245_TDATA = x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TDATA; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 49:23:@23096.4]
  assign io_sigsOut_smDoneIn_0 = x400_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@23010.4]
  assign io_sigsOut_smCtrCopyDone_0 = x400_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 168:125:@23029.4]
  assign x252_ctrchain_clock = clock; // @[:@22858.4]
  assign x252_ctrchain_reset = reset; // @[:@22859.4]
  assign x252_ctrchain_io_input_reset = x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@23028.4]
  assign x252_ctrchain_io_input_enable = _T_271 & x400_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@22980.4 SpatialBlocks.scala 159:42:@23027.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@22918.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@22919.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sm_io_enable = x400_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x400_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@23007.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x401_outr_UnitPipe.scala 66:50:@22953.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@23009.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x245_TREADY | x400_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@22981.4]
  assign x400_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x401_outr_UnitPipe.scala 70:48:@22959.4]
  assign RetimeWrapper_clock = clock; // @[:@22946.4]
  assign RetimeWrapper_reset = reset; // @[:@22947.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@22949.4]
  assign RetimeWrapper_io_in = x252_ctrchain_io_output_done; // @[package.scala 94:16:@22948.4]
  assign RetimeWrapper_1_clock = clock; // @[:@22988.4]
  assign RetimeWrapper_1_reset = reset; // @[:@22989.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@22991.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@22990.4]
  assign RetimeWrapper_2_clock = clock; // @[:@22996.4]
  assign RetimeWrapper_2_reset = reset; // @[:@22997.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@22999.4]
  assign RetimeWrapper_2_io_in = x400_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@22998.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@23031.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@23032.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TDATA = io_in_x244_TDATA; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 48:23:@23087.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TID = io_in_x244_TID; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 48:23:@23083.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x244_TDEST = io_in_x244_TDEST; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 48:23:@23082.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x245_TREADY = io_in_x245_TREADY; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 49:23:@23097.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x245_TREADY | x400_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 579:22:@23115.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 579:22:@23113.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x400_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 579:22:@23111.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x252_ctrchain_io_output_counts_1; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 579:22:@23106.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x252_ctrchain_io_output_counts_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 579:22:@23105.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x252_ctrchain_io_output_oobs_0; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 579:22:@23103.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x252_ctrchain_io_output_oobs_1; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 579:22:@23104.4]
  assign x400_inr_Foreach_SAMPLER_BOX_kernelx400_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x400_inr_Foreach_SAMPLER_BOX.scala 578:18:@23099.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@23129.2]
  input          clock, // @[:@23130.4]
  input          reset, // @[:@23131.4]
  input          io_in_x244_TVALID, // @[:@23132.4]
  output         io_in_x244_TREADY, // @[:@23132.4]
  input  [255:0] io_in_x244_TDATA, // @[:@23132.4]
  input  [7:0]   io_in_x244_TID, // @[:@23132.4]
  input  [7:0]   io_in_x244_TDEST, // @[:@23132.4]
  output         io_in_x245_TVALID, // @[:@23132.4]
  input          io_in_x245_TREADY, // @[:@23132.4]
  output [255:0] io_in_x245_TDATA, // @[:@23132.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@23132.4]
  input          io_sigsIn_smChildAcks_0, // @[:@23132.4]
  output         io_sigsOut_smDoneIn_0, // @[:@23132.4]
  input          io_rr // @[:@23132.4]
);
  wire  x401_outr_UnitPipe_sm_clock; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_reset; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_io_enable; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_io_done; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_io_parentAck; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_io_childAck_0; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  x401_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23326.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23326.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23326.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@23326.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@23326.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@23334.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@23334.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@23334.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@23334.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@23334.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_clock; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_reset; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TVALID; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TREADY; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire [255:0] x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TDATA; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire [7:0] x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TID; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire [7:0] x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TDEST; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TVALID; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TREADY; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire [255:0] x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TDATA; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_rr; // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
  wire  _T_246; // @[package.scala 96:25:@23331.4 package.scala 96:25:@23332.4]
  wire  _T_252; // @[package.scala 96:25:@23339.4 package.scala 96:25:@23340.4]
  wire  _T_255; // @[SpatialBlocks.scala 138:93:@23342.4]
  x401_outr_UnitPipe_sm x401_outr_UnitPipe_sm ( // @[sm_x401_outr_UnitPipe.scala 32:18:@23274.4]
    .clock(x401_outr_UnitPipe_sm_clock),
    .reset(x401_outr_UnitPipe_sm_reset),
    .io_enable(x401_outr_UnitPipe_sm_io_enable),
    .io_done(x401_outr_UnitPipe_sm_io_done),
    .io_parentAck(x401_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x401_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x401_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x401_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x401_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@23326.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@23334.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1 x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1 ( // @[sm_x401_outr_UnitPipe.scala 75:24:@23364.4]
    .clock(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_clock),
    .reset(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_reset),
    .io_in_x244_TVALID(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TVALID),
    .io_in_x244_TREADY(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TREADY),
    .io_in_x244_TDATA(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TDATA),
    .io_in_x244_TID(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TID),
    .io_in_x244_TDEST(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TDEST),
    .io_in_x245_TVALID(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TVALID),
    .io_in_x245_TREADY(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TREADY),
    .io_in_x245_TDATA(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TDATA),
    .io_sigsIn_smEnableOuts_0(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@23331.4 package.scala 96:25:@23332.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@23339.4 package.scala 96:25:@23340.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 138:93:@23342.4]
  assign io_in_x244_TREADY = x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TREADY; // @[sm_x401_outr_UnitPipe.scala 48:23:@23420.4]
  assign io_in_x245_TVALID = x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TVALID; // @[sm_x401_outr_UnitPipe.scala 49:23:@23430.4]
  assign io_in_x245_TDATA = x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TDATA; // @[sm_x401_outr_UnitPipe.scala 49:23:@23428.4]
  assign io_sigsOut_smDoneIn_0 = x401_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@23349.4]
  assign x401_outr_UnitPipe_sm_clock = clock; // @[:@23275.4]
  assign x401_outr_UnitPipe_sm_reset = reset; // @[:@23276.4]
  assign x401_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 140:18:@23346.4]
  assign x401_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@23348.4]
  assign x401_outr_UnitPipe_sm_io_doneIn_0 = x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@23318.4]
  assign x401_outr_UnitPipe_sm_io_ctrCopyDone_0 = x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@23363.4]
  assign RetimeWrapper_clock = clock; // @[:@23327.4]
  assign RetimeWrapper_reset = reset; // @[:@23328.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23330.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@23329.4]
  assign RetimeWrapper_1_clock = clock; // @[:@23335.4]
  assign RetimeWrapper_1_reset = reset; // @[:@23336.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@23338.4]
  assign RetimeWrapper_1_io_in = x401_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@23337.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_clock = clock; // @[:@23365.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_reset = reset; // @[:@23366.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TVALID = io_in_x244_TVALID; // @[sm_x401_outr_UnitPipe.scala 48:23:@23421.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TDATA = io_in_x244_TDATA; // @[sm_x401_outr_UnitPipe.scala 48:23:@23419.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TID = io_in_x244_TID; // @[sm_x401_outr_UnitPipe.scala 48:23:@23415.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x244_TDEST = io_in_x244_TDEST; // @[sm_x401_outr_UnitPipe.scala 48:23:@23414.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_in_x245_TREADY = io_in_x245_TREADY; // @[sm_x401_outr_UnitPipe.scala 49:23:@23429.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x401_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x401_outr_UnitPipe.scala 80:22:@23439.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x401_outr_UnitPipe_sm_io_childAck_0; // @[sm_x401_outr_UnitPipe.scala 80:22:@23437.4]
  assign x401_outr_UnitPipe_kernelx401_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x401_outr_UnitPipe.scala 79:18:@23431.4]
endmodule
module AccelUnit( // @[:@23459.2]
  input          clock, // @[:@23460.4]
  input          reset, // @[:@23461.4]
  input          io_enable, // @[:@23462.4]
  output         io_done, // @[:@23462.4]
  input          io_reset, // @[:@23462.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@23462.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@23462.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@23462.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@23462.4]
  output         io_memStreams_loads_0_data_ready, // @[:@23462.4]
  input          io_memStreams_loads_0_data_valid, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@23462.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@23462.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@23462.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@23462.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@23462.4]
  input          io_memStreams_stores_0_data_ready, // @[:@23462.4]
  output         io_memStreams_stores_0_data_valid, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@23462.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@23462.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@23462.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@23462.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@23462.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@23462.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@23462.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@23462.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@23462.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@23462.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@23462.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@23462.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@23462.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@23462.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@23462.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@23462.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@23462.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@23462.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@23462.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@23462.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@23462.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@23462.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@23462.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@23462.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@23462.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@23462.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@23462.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@23462.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@23462.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@23462.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@23462.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@23462.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@23462.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@23462.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@23462.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@23462.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@23462.4]
  output         io_heap_0_req_valid, // @[:@23462.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@23462.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@23462.4]
  input          io_heap_0_resp_valid, // @[:@23462.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@23462.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@23462.4]
  input  [63:0]  io_argIns_0, // @[:@23462.4]
  input  [63:0]  io_argIns_1, // @[:@23462.4]
  input          io_argOuts_0_port_ready, // @[:@23462.4]
  output         io_argOuts_0_port_valid, // @[:@23462.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@23462.4]
  input  [63:0]  io_argOuts_0_echo // @[:@23462.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@23625.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@23625.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@23625.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@23625.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23643.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23643.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23643.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@23643.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@23643.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@23652.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@23652.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@23652.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@23652.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@23652.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@23652.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@23691.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@23723.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@23723.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@23723.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@23723.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@23723.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_in_x244_TVALID; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_in_x244_TREADY; // @[sm_RootController.scala 73:24:@23785.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x244_TDATA; // @[sm_RootController.scala 73:24:@23785.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x244_TID; // @[sm_RootController.scala 73:24:@23785.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x244_TDEST; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_in_x245_TVALID; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_in_x245_TREADY; // @[sm_RootController.scala 73:24:@23785.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x245_TDATA; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@23785.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@23785.4]
  wire  _T_599; // @[package.scala 96:25:@23648.4 package.scala 96:25:@23649.4]
  wire  _T_664; // @[Main.scala 41:50:@23719.4]
  wire  _T_665; // @[Main.scala 41:59:@23720.4]
  wire  _T_677; // @[package.scala 100:49:@23740.4]
  reg  _T_680; // @[package.scala 48:56:@23741.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@23625.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@23643.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@23652.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@23691.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@23723.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@23785.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x244_TVALID(RootController_kernelRootController_concrete1_io_in_x244_TVALID),
    .io_in_x244_TREADY(RootController_kernelRootController_concrete1_io_in_x244_TREADY),
    .io_in_x244_TDATA(RootController_kernelRootController_concrete1_io_in_x244_TDATA),
    .io_in_x244_TID(RootController_kernelRootController_concrete1_io_in_x244_TID),
    .io_in_x244_TDEST(RootController_kernelRootController_concrete1_io_in_x244_TDEST),
    .io_in_x245_TVALID(RootController_kernelRootController_concrete1_io_in_x245_TVALID),
    .io_in_x245_TREADY(RootController_kernelRootController_concrete1_io_in_x245_TREADY),
    .io_in_x245_TDATA(RootController_kernelRootController_concrete1_io_in_x245_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@23648.4 package.scala 96:25:@23649.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@23719.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@23720.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@23740.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@23739.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x244_TREADY; // @[sm_RootController.scala 48:23:@23841.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x245_TVALID; // @[sm_RootController.scala 49:23:@23851.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x245_TDATA; // @[sm_RootController.scala 49:23:@23849.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:23:@23848.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:23:@23847.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:23:@23846.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:23:@23845.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:23:@23844.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:23:@23843.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@23626.4]
  assign SingleCounter_reset = reset; // @[:@23627.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@23641.4]
  assign RetimeWrapper_clock = clock; // @[:@23644.4]
  assign RetimeWrapper_reset = reset; // @[:@23645.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23647.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@23646.4]
  assign SRFF_clock = clock; // @[:@23653.4]
  assign SRFF_reset = reset; // @[:@23654.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@23879.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@23737.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@23738.4]
  assign RootController_sm_clock = clock; // @[:@23692.4]
  assign RootController_sm_reset = reset; // @[:@23693.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@23736.4 SpatialBlocks.scala 140:18:@23770.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@23764.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@23744.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@23761.4]
  assign RetimeWrapper_1_clock = clock; // @[:@23724.4]
  assign RetimeWrapper_1_reset = reset; // @[:@23725.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@23727.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@23726.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@23786.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@23787.4]
  assign RootController_kernelRootController_concrete1_io_in_x244_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 48:23:@23842.4]
  assign RootController_kernelRootController_concrete1_io_in_x244_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:23:@23840.4]
  assign RootController_kernelRootController_concrete1_io_in_x244_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:23:@23836.4]
  assign RootController_kernelRootController_concrete1_io_in_x244_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:23:@23835.4]
  assign RootController_kernelRootController_concrete1_io_in_x245_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:23:@23850.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 78:22:@23860.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 78:22:@23858.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 77:18:@23852.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@23881.2]
  input         clock, // @[:@23882.4]
  input         reset, // @[:@23883.4]
  input  [31:0] io_raddr, // @[:@23884.4]
  input         io_wen, // @[:@23884.4]
  input  [31:0] io_waddr, // @[:@23884.4]
  input  [63:0] io_wdata, // @[:@23884.4]
  output [63:0] io_rdata // @[:@23884.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@23886.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@23886.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@23886.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@23886.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@23886.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@23886.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@23886.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@23886.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@23886.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@23886.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@23886.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@23886.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@23887.4]
  assign accel_reset = reset; // @[:@23888.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
