// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLKclock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x744_TREADY(dontcare), // @[:@1298.4]
    .io_in_x744_TDATA({I_0,I_1,I_2,I_3,I_4,I_5,I_6,I_7}), // @[:@1298.4]
    .io_in_x744_TID(8'h0),
    .io_in_x744_TDEST(8'h0),
    .io_in_x745_TVALID(valid_down), // @[:@1298.4]
    .io_in_x745_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0,O_4_0_0,O_5_0_0,O_6_0_0,O_7_0_0}), // @[:@1298.4]
    .io_in_x745_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x752_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 311:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 315:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 315:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh3b); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh3b); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [7:0]  io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@512.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@512.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@512.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@532.4]
  assign SRAMVerilogSim_wdata = 8'h0; // @[SRAM.scala 190:20:@526.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@527.4]
  assign SRAMVerilogSim_wen = 1'h0; // @[SRAM.scala 188:18:@524.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@529.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@528.4]
  assign SRAMVerilogSim_waddr = 21'h0; // @[SRAM.scala 189:20:@525.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@523.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@546.2]
  input         clock, // @[:@547.4]
  input         reset, // @[:@548.4]
  input         io_flow, // @[:@549.4]
  input  [20:0] io_in, // @[:@549.4]
  output [20:0] io_out // @[:@549.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@551.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@551.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@564.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@563.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@562.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@561.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@560.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@558.4]
endmodule
module Mem1D( // @[:@566.2]
  input         clock, // @[:@567.4]
  input         reset, // @[:@568.4]
  input  [20:0] io_r_ofs_0, // @[:@569.4]
  input         io_r_backpressure, // @[:@569.4]
  output [7:0]  io_output // @[:@569.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@573.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@573.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@573.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@573.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@576.4]
  SRAM SRAM ( // @[MemPrimitives.scala 705:21:@573.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@576.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@589.4]
  assign SRAM_clock = clock; // @[:@574.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@583.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@588.4]
  assign RetimeWrapper_clock = clock; // @[:@577.4]
  assign RetimeWrapper_reset = reset; // @[:@578.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@580.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@579.4]
endmodule
module StickySelects( // @[:@591.2]
  input   io_ins_0, // @[:@594.4]
  output  io_outs_0 // @[:@594.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@596.4]
endmodule
module RetimeWrapper_6( // @[:@610.2]
  input   clock, // @[:@611.4]
  input   reset, // @[:@612.4]
  input   io_flow, // @[:@613.4]
  input   io_in, // @[:@613.4]
  output  io_out // @[:@613.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@615.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@615.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@628.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@627.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@626.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@625.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@624.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@622.4]
endmodule
module x746_outbuf_0( // @[:@630.2]
  input         clock, // @[:@631.4]
  input         reset, // @[:@632.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@633.4]
  input         io_rPort_0_en_0, // @[:@633.4]
  input         io_rPort_0_backpressure, // @[:@633.4]
  output [7:0]  io_rPort_0_output_0 // @[:@633.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@648.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@648.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@648.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@688.4]
  wire  _T_76; // @[MemPrimitives.scala 123:41:@678.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@680.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@648.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@674.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@688.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@678.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@680.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@695.4]
  assign Mem1D_clock = clock; // @[:@649.4]
  assign Mem1D_reset = reset; // @[:@650.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 127:28:@684.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 128:32:@685.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@677.4]
  assign RetimeWrapper_clock = clock; // @[:@689.4]
  assign RetimeWrapper_reset = reset; // @[:@690.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@692.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@691.4]
endmodule
module x1251_sm( // @[:@839.2]
  input   clock, // @[:@840.4]
  input   reset, // @[:@841.4]
  input   io_enable, // @[:@842.4]
  output  io_done, // @[:@842.4]
  input   io_ctrDone, // @[:@842.4]
  output  io_ctrInc, // @[:@842.4]
  input   io_parentAck, // @[:@842.4]
  input   io_doneIn_0, // @[:@842.4]
  input   io_doneIn_1, // @[:@842.4]
  output  io_enableOut_0, // @[:@842.4]
  output  io_enableOut_1, // @[:@842.4]
  output  io_childAck_0, // @[:@842.4]
  output  io_childAck_1 // @[:@842.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@845.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@848.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@851.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@854.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@886.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1004.4]
  wire  allDone; // @[Controllers.scala 80:47:@857.4]
  wire  synchronize; // @[Controllers.scala 146:56:@911.4]
  wire  _T_127; // @[Controllers.scala 150:35:@913.4]
  wire  _T_129; // @[Controllers.scala 150:60:@914.4]
  wire  _T_130; // @[Controllers.scala 150:58:@915.4]
  wire  _T_132; // @[Controllers.scala 150:76:@916.4]
  wire  _T_133; // @[Controllers.scala 150:74:@917.4]
  wire  _T_135; // @[Controllers.scala 150:97:@918.4]
  wire  _T_136; // @[Controllers.scala 150:95:@919.4]
  wire  _T_152; // @[Controllers.scala 150:35:@937.4]
  wire  _T_154; // @[Controllers.scala 150:60:@938.4]
  wire  _T_155; // @[Controllers.scala 150:58:@939.4]
  wire  _T_157; // @[Controllers.scala 150:76:@940.4]
  wire  _T_158; // @[Controllers.scala 150:74:@941.4]
  wire  _T_161; // @[Controllers.scala 150:95:@943.4]
  wire  _T_179; // @[Controllers.scala 213:68:@965.4]
  wire  _T_181; // @[Controllers.scala 213:90:@967.4]
  wire  _T_183; // @[Controllers.scala 213:132:@969.4]
  wire  _T_184; // @[Controllers.scala 213:130:@970.4]
  wire  _T_185; // @[Controllers.scala 213:156:@971.4]
  wire  _T_187; // @[Controllers.scala 213:68:@974.4]
  wire  _T_189; // @[Controllers.scala 213:90:@976.4]
  wire  _T_196; // @[package.scala 100:49:@982.4]
  reg  _T_199; // @[package.scala 48:56:@983.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@985.4]
  reg  _T_213; // @[package.scala 48:56:@1001.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@845.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@848.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@851.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@854.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@883.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@886.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@987.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1004.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@857.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@911.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@913.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@914.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@915.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@916.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@917.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@918.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@919.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@937.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@938.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@939.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@940.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@941.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@943.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@965.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@967.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@969.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@970.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@971.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@974.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@976.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@982.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@985.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1011.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@910.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@973.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@981.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@962.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@964.4]
  assign active_0_clock = clock; // @[:@846.4]
  assign active_0_reset = reset; // @[:@847.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@922.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@926.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@860.4]
  assign active_1_clock = clock; // @[:@849.4]
  assign active_1_reset = reset; // @[:@850.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@946.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@950.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@861.4]
  assign done_0_clock = clock; // @[:@852.4]
  assign done_0_reset = reset; // @[:@853.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@936.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@872.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@862.4]
  assign done_1_clock = clock; // @[:@855.4]
  assign done_1_reset = reset; // @[:@856.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@960.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@881.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@863.4]
  assign iterDone_0_clock = clock; // @[:@884.4]
  assign iterDone_0_reset = reset; // @[:@885.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@932.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@899.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@889.4]
  assign iterDone_1_clock = clock; // @[:@887.4]
  assign iterDone_1_reset = reset; // @[:@888.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@956.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@908.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@890.4]
  assign RetimeWrapper_clock = clock; // @[:@988.4]
  assign RetimeWrapper_reset = reset; // @[:@989.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@991.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@990.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1005.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1006.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1008.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1007.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x1158_outr_UnitPipe_sm( // @[:@1428.2]
  input   clock, // @[:@1429.4]
  input   reset, // @[:@1430.4]
  input   io_enable, // @[:@1431.4]
  output  io_done, // @[:@1431.4]
  input   io_parentAck, // @[:@1431.4]
  input   io_doneIn_0, // @[:@1431.4]
  input   io_doneIn_1, // @[:@1431.4]
  output  io_enableOut_0, // @[:@1431.4]
  output  io_enableOut_1, // @[:@1431.4]
  output  io_childAck_0, // @[:@1431.4]
  output  io_childAck_1, // @[:@1431.4]
  input   io_ctrCopyDone_0, // @[:@1431.4]
  input   io_ctrCopyDone_1 // @[:@1431.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1434.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1437.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1440.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1443.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1475.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1681.4]
  wire  allDone; // @[Controllers.scala 80:47:@1446.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1500.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1501.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1502.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1503.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1504.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1507.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1509.4]
  wire  _T_148; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1524.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1525.4]
  wire  _T_160; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  wire  _T_178; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1556.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1557.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1569.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1570.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1571.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1572.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1573.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1576.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1578.4]
  wire  _T_216; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1593.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1594.4]
  wire  _T_228; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  wire  _T_246; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1625.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1626.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1642.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1644.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1646.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1651.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1653.4]
  wire  _T_282; // @[package.scala 100:49:@1659.4]
  reg  _T_285; // @[package.scala 48:56:@1660.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1662.4]
  reg  _T_299; // @[package.scala 48:56:@1678.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1434.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1437.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1440.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1443.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1472.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1475.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1516.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1530.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1548.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1585.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1599.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1617.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1664.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1681.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1446.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1500.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1501.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1502.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1503.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1504.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1507.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1509.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1524.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1525.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1556.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1557.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1569.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1570.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1571.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1572.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1573.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1576.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1578.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1593.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1594.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1625.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1626.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1642.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1644.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1646.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1651.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1653.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1659.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1662.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1688.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1650.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1658.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1639.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1641.4]
  assign active_0_clock = clock; // @[:@1435.4]
  assign active_0_reset = reset; // @[:@1436.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1511.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1515.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1449.4]
  assign active_1_clock = clock; // @[:@1438.4]
  assign active_1_reset = reset; // @[:@1439.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1580.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1584.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1450.4]
  assign done_0_clock = clock; // @[:@1441.4]
  assign done_0_reset = reset; // @[:@1442.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1561.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1461.4 Controllers.scala 170:32:@1568.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1451.4]
  assign done_1_clock = clock; // @[:@1444.4]
  assign done_1_reset = reset; // @[:@1445.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1630.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1470.4 Controllers.scala 170:32:@1637.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1452.4]
  assign iterDone_0_clock = clock; // @[:@1473.4]
  assign iterDone_0_reset = reset; // @[:@1474.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1529.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1488.4 Controllers.scala 168:36:@1545.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1478.4]
  assign iterDone_1_clock = clock; // @[:@1476.4]
  assign iterDone_1_reset = reset; // @[:@1477.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1598.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1497.4 Controllers.scala 168:36:@1614.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1479.4]
  assign RetimeWrapper_clock = clock; // @[:@1517.4]
  assign RetimeWrapper_reset = reset; // @[:@1518.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1520.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1519.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1531.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1532.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1534.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1533.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1549.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1550.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1552.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1551.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1586.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1587.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1589.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1588.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1600.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1601.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1603.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1602.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1618.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1619.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1621.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1620.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1665.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1666.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1668.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1667.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1682.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1683.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1685.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1684.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1917.2]
  input   clock, // @[:@1918.4]
  input   reset, // @[:@1919.4]
  input   io_input_inc_en_0, // @[:@1920.4]
  input   io_input_dinc_en_0, // @[:@1920.4]
  output  io_output_full // @[:@1920.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1922.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1923.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1924.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1925.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1925.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1926.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1927.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1928.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1928.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1929.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1930.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1923.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1924.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1925.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1925.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1926.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1927.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1928.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1928.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1929.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1930.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1944.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x747_fifoinraw_0( // @[:@2067.2]
  input   clock, // @[:@2068.4]
  input   reset // @[:@2069.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2114.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2114.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2115.4]
  assign elements_reset = reset; // @[:@2116.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 384:79:@2126.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2127.4]
endmodule
module x748_fifoinpacked_0( // @[:@2490.2]
  input   clock, // @[:@2491.4]
  input   reset, // @[:@2492.4]
  input   io_wPort_0_en_0, // @[:@2493.4]
  output  io_full, // @[:@2493.4]
  input   io_active_0_in, // @[:@2493.4]
  output  io_active_0_out // @[:@2493.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2537.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2537.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 429:39:@2611.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 427:129:@2609.4]
  assign elements_clock = clock; // @[:@2538.4]
  assign elements_reset = reset; // @[:@2539.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 384:79:@2549.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2550.4]
endmodule
module FF_7( // @[:@3040.2]
  input         clock, // @[:@3041.4]
  input         reset, // @[:@3042.4]
  output [12:0] io_rPort_0_output_0, // @[:@3043.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3043.4]
  input         io_wPort_0_reset, // @[:@3043.4]
  input         io_wPort_0_en_0 // @[:@3043.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 311:19:@3058.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 315:32:@3060.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 315:12:@3061.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@3060.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 315:12:@3061.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@3063.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3078.2]
  input         clock, // @[:@3079.4]
  input         reset, // @[:@3080.4]
  input         io_setup_saturate, // @[:@3081.4]
  input         io_input_reset, // @[:@3081.4]
  input         io_input_enable, // @[:@3081.4]
  output [12:0] io_output_count_0, // @[:@3081.4]
  output        io_output_oobs_0, // @[:@3081.4]
  output        io_output_done, // @[:@3081.4]
  output        io_output_saturated // @[:@3081.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3094.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3110.4]
  wire  _T_36; // @[Counter.scala 264:45:@3113.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3138.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3139.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3140.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3141.4]
  wire  _T_57; // @[Counter.scala 293:18:@3143.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3151.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3153.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3154.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3155.4]
  wire  _T_75; // @[Counter.scala 322:102:@3159.4]
  wire  _T_77; // @[Counter.scala 322:130:@3160.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3094.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3110.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3113.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3138.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3139.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3140.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3141.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3143.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3151.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3153.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3154.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3155.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3159.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3160.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3158.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3162.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3164.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3167.4]
  assign bases_0_clock = clock; // @[:@3095.4]
  assign bases_0_reset = reset; // @[:@3096.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3157.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3136.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3137.4]
  assign SRFF_clock = clock; // @[:@3111.4]
  assign SRFF_reset = reset; // @[:@3112.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3115.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3117.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3118.4]
endmodule
module SingleCounter_2( // @[:@3207.2]
  input         clock, // @[:@3208.4]
  input         reset, // @[:@3209.4]
  input         io_setup_saturate, // @[:@3210.4]
  input         io_input_reset, // @[:@3210.4]
  input         io_input_enable, // @[:@3210.4]
  output [12:0] io_output_count_0, // @[:@3210.4]
  output        io_output_oobs_0, // @[:@3210.4]
  output        io_output_done // @[:@3210.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3223.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3239.4]
  wire  _T_36; // @[Counter.scala 264:45:@3242.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3267.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3268.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3269.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3270.4]
  wire  _T_57; // @[Counter.scala 293:18:@3272.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3280.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3282.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3283.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3284.4]
  wire  _T_75; // @[Counter.scala 322:102:@3288.4]
  wire  _T_77; // @[Counter.scala 322:130:@3289.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3223.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3239.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3242.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3267.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh8); // @[Counter.scala 291:33:@3268.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh8); // @[Counter.scala 291:33:@3269.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3270.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3272.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3280.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3282.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3283.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3284.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3288.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3289.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3287.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3291.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3293.4]
  assign bases_0_clock = clock; // @[:@3224.4]
  assign bases_0_reset = reset; // @[:@3225.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3286.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3265.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3266.4]
  assign SRFF_clock = clock; // @[:@3240.4]
  assign SRFF_reset = reset; // @[:@3241.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3244.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3246.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3247.4]
endmodule
module x752_ctrchain( // @[:@3298.2]
  input         clock, // @[:@3299.4]
  input         reset, // @[:@3300.4]
  input         io_input_reset, // @[:@3301.4]
  input         io_input_enable, // @[:@3301.4]
  output [12:0] io_output_counts_1, // @[:@3301.4]
  output [12:0] io_output_counts_0, // @[:@3301.4]
  output        io_output_oobs_0, // @[:@3301.4]
  output        io_output_oobs_1, // @[:@3301.4]
  output        io_output_done // @[:@3301.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3303.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3306.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3306.4]
  wire  isDone; // @[Counter.scala 541:51:@3323.4]
  reg  wasDone; // @[Counter.scala 542:24:@3324.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3332.4]
  wire  _T_66; // @[Counter.scala 546:80:@3333.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3338.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3339.4]
  wire  _T_74; // @[Counter.scala 551:19:@3340.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3303.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3306.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3323.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3332.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3333.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3339.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3340.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3345.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3342.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3344.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3347.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3335.4]
  assign ctrs_0_clock = clock; // @[:@3304.4]
  assign ctrs_0_reset = reset; // @[:@3305.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3320.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3312.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3319.4]
  assign ctrs_1_clock = clock; // @[:@3307.4]
  assign ctrs_1_reset = reset; // @[:@3308.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3322.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3316.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3317.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3387.2]
  input   clock, // @[:@3388.4]
  input   reset, // @[:@3389.4]
  input   io_flow, // @[:@3390.4]
  input   io_in, // @[:@3390.4]
  output  io_out // @[:@3390.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3392.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3405.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3404.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3403.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3402.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3401.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3399.4]
endmodule
module RetimeWrapper_25( // @[:@3515.2]
  input   clock, // @[:@3516.4]
  input   reset, // @[:@3517.4]
  input   io_flow, // @[:@3518.4]
  input   io_in, // @[:@3518.4]
  output  io_out // @[:@3518.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3520.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3533.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3532.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3531.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3530.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3529.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3527.4]
endmodule
module x794_inr_Foreach_sm( // @[:@3535.2]
  input   clock, // @[:@3536.4]
  input   reset, // @[:@3537.4]
  input   io_enable, // @[:@3538.4]
  output  io_done, // @[:@3538.4]
  output  io_doneLatch, // @[:@3538.4]
  input   io_ctrDone, // @[:@3538.4]
  output  io_datapathEn, // @[:@3538.4]
  output  io_ctrInc, // @[:@3538.4]
  output  io_ctrRst, // @[:@3538.4]
  input   io_parentAck, // @[:@3538.4]
  input   io_backpressure, // @[:@3538.4]
  input   io_break // @[:@3538.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3540.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3540.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3543.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3543.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3635.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3548.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3549.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3550.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3551.4]
  wire  _T_100; // @[package.scala 100:49:@3568.4]
  reg  _T_103; // @[package.scala 48:56:@3569.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  wire  _T_110; // @[package.scala 100:49:@3584.4]
  reg  _T_113; // @[package.scala 48:56:@3585.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3587.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3592.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3593.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3596.4]
  wire  _T_124; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  wire  _T_126; // @[package.scala 100:49:@3606.4]
  reg  _T_129; // @[package.scala 48:56:@3607.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3629.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3631.4]
  reg  _T_153; // @[package.scala 48:56:@3632.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3642.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3643.4]
  SRFF active ( // @[Controllers.scala 261:22:@3540.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3543.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3577.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3599.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3611.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3619.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3635.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3548.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3549.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3550.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3551.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3568.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3584.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3587.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3592.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3593.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3596.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3606.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3631.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3642.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3643.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3610.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3645.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3595.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3598.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3590.4]
  assign active_clock = clock; // @[:@3541.4]
  assign active_reset = reset; // @[:@3542.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3553.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3557.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3558.4]
  assign done_clock = clock; // @[:@3544.4]
  assign done_reset = reset; // @[:@3545.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3573.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3566.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3567.4]
  assign RetimeWrapper_clock = clock; // @[:@3578.4]
  assign RetimeWrapper_reset = reset; // @[:@3579.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3581.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3580.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3600.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3601.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3603.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3602.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3612.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3613.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3615.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3614.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3620.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3621.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3623.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3622.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3636.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3637.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3639.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3638.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3752.2]
  input  [31:0] io_a, // @[:@3755.4]
  output [31:0] io_b // @[:@3755.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3768.4]
endmodule
module _( // @[:@3770.2]
  input  [31:0] io_b, // @[:@3773.4]
  output [31:0] io_result // @[:@3773.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3778.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3778.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3778.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3791.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3786.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@3834.2]
  input  [31:0] io_a, // @[:@3837.4]
  output [32:0] io_b // @[:@3837.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3847.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3847.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@3852.4]
endmodule
module __2( // @[:@3854.2]
  input  [31:0] io_b, // @[:@3857.4]
  output [32:0] io_result // @[:@3857.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3862.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3862.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3862.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3875.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3870.4]
endmodule
module RetimeWrapper_29( // @[:@3932.2]
  input         clock, // @[:@3933.4]
  input         reset, // @[:@3934.4]
  input         io_flow, // @[:@3935.4]
  input  [31:0] io_in, // @[:@3935.4]
  output [31:0] io_out // @[:@3935.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3937.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3950.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3949.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3948.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3947.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3946.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3944.4]
endmodule
module fix2fixBox( // @[:@3952.2]
  input         clock, // @[:@3953.4]
  input         reset, // @[:@3954.4]
  input  [32:0] io_a, // @[:@3955.4]
  input         io_flow, // @[:@3955.4]
  output [31:0] io_b // @[:@3955.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3968.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3968.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3975.4]
  assign RetimeWrapper_clock = clock; // @[:@3969.4]
  assign RetimeWrapper_reset = reset; // @[:@3970.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3972.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3971.4]
endmodule
module x1207_sub( // @[:@3977.2]
  input         clock, // @[:@3978.4]
  input         reset, // @[:@3979.4]
  input  [31:0] io_a, // @[:@3980.4]
  input  [31:0] io_b, // @[:@3980.4]
  input         io_flow, // @[:@3980.4]
  output [31:0] io_result // @[:@3980.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@3988.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@3988.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@3995.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@3995.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4014.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4014.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4014.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@4002.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@4003.4]
  __2 _ ( // @[Math.scala 709:24:@3988.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@3995.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@4014.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@4002.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@4003.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4022.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@3991.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@3998.4]
  assign fix2fixBox_clock = clock; // @[:@4015.4]
  assign fix2fixBox_reset = reset; // @[:@4016.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4017.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4020.4]
endmodule
module x758_sum( // @[:@4199.2]
  input         clock, // @[:@4200.4]
  input         reset, // @[:@4201.4]
  input  [31:0] io_a, // @[:@4202.4]
  input  [31:0] io_b, // @[:@4202.4]
  input         io_flow, // @[:@4202.4]
  output [31:0] io_result // @[:@4202.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@4210.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@4210.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@4217.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@4217.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4235.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4235.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4235.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4224.4]
  __2 _ ( // @[Math.scala 709:24:@4210.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@4217.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@4235.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4224.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4243.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@4213.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@4220.4]
  assign fix2fixBox_clock = clock; // @[:@4236.4]
  assign fix2fixBox_reset = reset; // @[:@4237.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4238.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4241.4]
endmodule
module x794_inr_Foreach_kernelx794_inr_Foreach_concrete1( // @[:@7693.2]
  input         clock, // @[:@7694.4]
  input         reset, // @[:@7695.4]
  output        io_in_x748_fifoinpacked_0_wPort_0_en_0, // @[:@7696.4]
  input         io_in_x748_fifoinpacked_0_full, // @[:@7696.4]
  output        io_in_x748_fifoinpacked_0_active_0_in, // @[:@7696.4]
  input         io_in_x748_fifoinpacked_0_active_0_out, // @[:@7696.4]
  input         io_sigsIn_backpressure, // @[:@7696.4]
  input         io_sigsIn_datapathEn, // @[:@7696.4]
  input         io_sigsIn_break, // @[:@7696.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@7696.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@7696.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@7696.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@7696.4]
  input         io_rr // @[:@7696.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@7730.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@7730.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@7742.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@7742.4]
  wire  x1207_sub_1_clock; // @[Math.scala 191:24:@7769.4]
  wire  x1207_sub_1_reset; // @[Math.scala 191:24:@7769.4]
  wire [31:0] x1207_sub_1_io_a; // @[Math.scala 191:24:@7769.4]
  wire [31:0] x1207_sub_1_io_b; // @[Math.scala 191:24:@7769.4]
  wire  x1207_sub_1_io_flow; // @[Math.scala 191:24:@7769.4]
  wire [31:0] x1207_sub_1_io_result; // @[Math.scala 191:24:@7769.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7779.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7779.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7779.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7779.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7779.4]
  wire  x758_sum_1_clock; // @[Math.scala 150:24:@7788.4]
  wire  x758_sum_1_reset; // @[Math.scala 150:24:@7788.4]
  wire [31:0] x758_sum_1_io_a; // @[Math.scala 150:24:@7788.4]
  wire [31:0] x758_sum_1_io_b; // @[Math.scala 150:24:@7788.4]
  wire  x758_sum_1_io_flow; // @[Math.scala 150:24:@7788.4]
  wire [31:0] x758_sum_1_io_result; // @[Math.scala 150:24:@7788.4]
  wire  x759_sum_1_clock; // @[Math.scala 150:24:@7800.4]
  wire  x759_sum_1_reset; // @[Math.scala 150:24:@7800.4]
  wire [31:0] x759_sum_1_io_a; // @[Math.scala 150:24:@7800.4]
  wire [31:0] x759_sum_1_io_b; // @[Math.scala 150:24:@7800.4]
  wire  x759_sum_1_io_flow; // @[Math.scala 150:24:@7800.4]
  wire [31:0] x759_sum_1_io_result; // @[Math.scala 150:24:@7800.4]
  wire  x1209_sum_1_clock; // @[Math.scala 150:24:@7815.4]
  wire  x1209_sum_1_reset; // @[Math.scala 150:24:@7815.4]
  wire [31:0] x1209_sum_1_io_a; // @[Math.scala 150:24:@7815.4]
  wire [31:0] x1209_sum_1_io_b; // @[Math.scala 150:24:@7815.4]
  wire  x1209_sum_1_io_flow; // @[Math.scala 150:24:@7815.4]
  wire [31:0] x1209_sum_1_io_result; // @[Math.scala 150:24:@7815.4]
  wire  x763_sum_1_clock; // @[Math.scala 150:24:@7847.4]
  wire  x763_sum_1_reset; // @[Math.scala 150:24:@7847.4]
  wire [31:0] x763_sum_1_io_a; // @[Math.scala 150:24:@7847.4]
  wire [31:0] x763_sum_1_io_b; // @[Math.scala 150:24:@7847.4]
  wire  x763_sum_1_io_flow; // @[Math.scala 150:24:@7847.4]
  wire [31:0] x763_sum_1_io_result; // @[Math.scala 150:24:@7847.4]
  wire  x1212_sum_1_clock; // @[Math.scala 150:24:@7862.4]
  wire  x1212_sum_1_reset; // @[Math.scala 150:24:@7862.4]
  wire [31:0] x1212_sum_1_io_a; // @[Math.scala 150:24:@7862.4]
  wire [31:0] x1212_sum_1_io_b; // @[Math.scala 150:24:@7862.4]
  wire  x1212_sum_1_io_flow; // @[Math.scala 150:24:@7862.4]
  wire [31:0] x1212_sum_1_io_result; // @[Math.scala 150:24:@7862.4]
  wire  x767_sum_1_clock; // @[Math.scala 150:24:@7894.4]
  wire  x767_sum_1_reset; // @[Math.scala 150:24:@7894.4]
  wire [31:0] x767_sum_1_io_a; // @[Math.scala 150:24:@7894.4]
  wire [31:0] x767_sum_1_io_b; // @[Math.scala 150:24:@7894.4]
  wire  x767_sum_1_io_flow; // @[Math.scala 150:24:@7894.4]
  wire [31:0] x767_sum_1_io_result; // @[Math.scala 150:24:@7894.4]
  wire  x1215_sum_1_clock; // @[Math.scala 150:24:@7909.4]
  wire  x1215_sum_1_reset; // @[Math.scala 150:24:@7909.4]
  wire [31:0] x1215_sum_1_io_a; // @[Math.scala 150:24:@7909.4]
  wire [31:0] x1215_sum_1_io_b; // @[Math.scala 150:24:@7909.4]
  wire  x1215_sum_1_io_flow; // @[Math.scala 150:24:@7909.4]
  wire [31:0] x1215_sum_1_io_result; // @[Math.scala 150:24:@7909.4]
  wire  x771_sum_1_clock; // @[Math.scala 150:24:@7941.4]
  wire  x771_sum_1_reset; // @[Math.scala 150:24:@7941.4]
  wire [31:0] x771_sum_1_io_a; // @[Math.scala 150:24:@7941.4]
  wire [31:0] x771_sum_1_io_b; // @[Math.scala 150:24:@7941.4]
  wire  x771_sum_1_io_flow; // @[Math.scala 150:24:@7941.4]
  wire [31:0] x771_sum_1_io_result; // @[Math.scala 150:24:@7941.4]
  wire  x1218_sum_1_clock; // @[Math.scala 150:24:@7956.4]
  wire  x1218_sum_1_reset; // @[Math.scala 150:24:@7956.4]
  wire [31:0] x1218_sum_1_io_a; // @[Math.scala 150:24:@7956.4]
  wire [31:0] x1218_sum_1_io_b; // @[Math.scala 150:24:@7956.4]
  wire  x1218_sum_1_io_flow; // @[Math.scala 150:24:@7956.4]
  wire [31:0] x1218_sum_1_io_result; // @[Math.scala 150:24:@7956.4]
  wire  x775_sum_1_clock; // @[Math.scala 150:24:@7988.4]
  wire  x775_sum_1_reset; // @[Math.scala 150:24:@7988.4]
  wire [31:0] x775_sum_1_io_a; // @[Math.scala 150:24:@7988.4]
  wire [31:0] x775_sum_1_io_b; // @[Math.scala 150:24:@7988.4]
  wire  x775_sum_1_io_flow; // @[Math.scala 150:24:@7988.4]
  wire [31:0] x775_sum_1_io_result; // @[Math.scala 150:24:@7988.4]
  wire  x1221_sum_1_clock; // @[Math.scala 150:24:@8003.4]
  wire  x1221_sum_1_reset; // @[Math.scala 150:24:@8003.4]
  wire [31:0] x1221_sum_1_io_a; // @[Math.scala 150:24:@8003.4]
  wire [31:0] x1221_sum_1_io_b; // @[Math.scala 150:24:@8003.4]
  wire  x1221_sum_1_io_flow; // @[Math.scala 150:24:@8003.4]
  wire [31:0] x1221_sum_1_io_result; // @[Math.scala 150:24:@8003.4]
  wire  x779_sum_1_clock; // @[Math.scala 150:24:@8035.4]
  wire  x779_sum_1_reset; // @[Math.scala 150:24:@8035.4]
  wire [31:0] x779_sum_1_io_a; // @[Math.scala 150:24:@8035.4]
  wire [31:0] x779_sum_1_io_b; // @[Math.scala 150:24:@8035.4]
  wire  x779_sum_1_io_flow; // @[Math.scala 150:24:@8035.4]
  wire [31:0] x779_sum_1_io_result; // @[Math.scala 150:24:@8035.4]
  wire  x1224_sum_1_clock; // @[Math.scala 150:24:@8050.4]
  wire  x1224_sum_1_reset; // @[Math.scala 150:24:@8050.4]
  wire [31:0] x1224_sum_1_io_a; // @[Math.scala 150:24:@8050.4]
  wire [31:0] x1224_sum_1_io_b; // @[Math.scala 150:24:@8050.4]
  wire  x1224_sum_1_io_flow; // @[Math.scala 150:24:@8050.4]
  wire [31:0] x1224_sum_1_io_result; // @[Math.scala 150:24:@8050.4]
  wire  x783_sum_1_clock; // @[Math.scala 150:24:@8082.4]
  wire  x783_sum_1_reset; // @[Math.scala 150:24:@8082.4]
  wire [31:0] x783_sum_1_io_a; // @[Math.scala 150:24:@8082.4]
  wire [31:0] x783_sum_1_io_b; // @[Math.scala 150:24:@8082.4]
  wire  x783_sum_1_io_flow; // @[Math.scala 150:24:@8082.4]
  wire [31:0] x783_sum_1_io_result; // @[Math.scala 150:24:@8082.4]
  wire  x1227_sum_1_clock; // @[Math.scala 150:24:@8097.4]
  wire  x1227_sum_1_reset; // @[Math.scala 150:24:@8097.4]
  wire [31:0] x1227_sum_1_io_a; // @[Math.scala 150:24:@8097.4]
  wire [31:0] x1227_sum_1_io_b; // @[Math.scala 150:24:@8097.4]
  wire  x1227_sum_1_io_flow; // @[Math.scala 150:24:@8097.4]
  wire [31:0] x1227_sum_1_io_result; // @[Math.scala 150:24:@8097.4]
  wire  x787_sum_1_clock; // @[Math.scala 150:24:@8129.4]
  wire  x787_sum_1_reset; // @[Math.scala 150:24:@8129.4]
  wire [31:0] x787_sum_1_io_a; // @[Math.scala 150:24:@8129.4]
  wire [31:0] x787_sum_1_io_b; // @[Math.scala 150:24:@8129.4]
  wire  x787_sum_1_io_flow; // @[Math.scala 150:24:@8129.4]
  wire [31:0] x787_sum_1_io_result; // @[Math.scala 150:24:@8129.4]
  wire  x1230_sum_1_clock; // @[Math.scala 150:24:@8144.4]
  wire  x1230_sum_1_reset; // @[Math.scala 150:24:@8144.4]
  wire [31:0] x1230_sum_1_io_a; // @[Math.scala 150:24:@8144.4]
  wire [31:0] x1230_sum_1_io_b; // @[Math.scala 150:24:@8144.4]
  wire  x1230_sum_1_io_flow; // @[Math.scala 150:24:@8144.4]
  wire [31:0] x1230_sum_1_io_result; // @[Math.scala 150:24:@8144.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@8192.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@8192.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@8192.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@8192.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@8192.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@8201.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@8201.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@8201.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@8201.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@8201.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@8212.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@8212.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@8212.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@8212.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@8212.4]
  wire  _T_328; // @[sm_x794_inr_Foreach.scala 64:22:@7755.4]
  wire  _T_329; // @[sm_x794_inr_Foreach.scala 64:59:@7756.4]
  wire [31:0] b753_number; // @[Math.scala 712:22:@7735.4 Math.scala 713:14:@7736.4]
  wire [42:0] _GEN_0; // @[Math.scala 450:32:@7760.4]
  wire [42:0] _T_333; // @[Math.scala 450:32:@7760.4]
  wire [38:0] _GEN_1; // @[Math.scala 450:32:@7765.4]
  wire [38:0] _T_337; // @[Math.scala 450:32:@7765.4]
  wire [31:0] x759_sum_number; // @[Math.scala 154:22:@7806.4 Math.scala 155:14:@7807.4]
  wire [33:0] _GEN_2; // @[Math.scala 450:32:@7811.4]
  wire [33:0] _T_357; // @[Math.scala 450:32:@7811.4]
  wire [31:0] x763_sum_number; // @[Math.scala 154:22:@7853.4 Math.scala 155:14:@7854.4]
  wire [33:0] _GEN_3; // @[Math.scala 450:32:@7858.4]
  wire [33:0] _T_386; // @[Math.scala 450:32:@7858.4]
  wire [31:0] x767_sum_number; // @[Math.scala 154:22:@7900.4 Math.scala 155:14:@7901.4]
  wire [33:0] _GEN_4; // @[Math.scala 450:32:@7905.4]
  wire [33:0] _T_415; // @[Math.scala 450:32:@7905.4]
  wire [31:0] x771_sum_number; // @[Math.scala 154:22:@7947.4 Math.scala 155:14:@7948.4]
  wire [33:0] _GEN_5; // @[Math.scala 450:32:@7952.4]
  wire [33:0] _T_444; // @[Math.scala 450:32:@7952.4]
  wire [31:0] x775_sum_number; // @[Math.scala 154:22:@7994.4 Math.scala 155:14:@7995.4]
  wire [33:0] _GEN_6; // @[Math.scala 450:32:@7999.4]
  wire [33:0] _T_473; // @[Math.scala 450:32:@7999.4]
  wire [31:0] x779_sum_number; // @[Math.scala 154:22:@8041.4 Math.scala 155:14:@8042.4]
  wire [33:0] _GEN_7; // @[Math.scala 450:32:@8046.4]
  wire [33:0] _T_502; // @[Math.scala 450:32:@8046.4]
  wire [31:0] x783_sum_number; // @[Math.scala 154:22:@8088.4 Math.scala 155:14:@8089.4]
  wire [33:0] _GEN_8; // @[Math.scala 450:32:@8093.4]
  wire [33:0] _T_531; // @[Math.scala 450:32:@8093.4]
  wire [31:0] x787_sum_number; // @[Math.scala 154:22:@8135.4 Math.scala 155:14:@8136.4]
  wire [33:0] _GEN_9; // @[Math.scala 450:32:@8140.4]
  wire [33:0] _T_560; // @[Math.scala 450:32:@8140.4]
  wire  _T_608; // @[sm_x794_inr_Foreach.scala 171:135:@8209.4]
  wire  _T_612; // @[package.scala 96:25:@8217.4 package.scala 96:25:@8218.4]
  wire  _T_614; // @[implicits.scala 55:10:@8219.4]
  wire  _T_615; // @[sm_x794_inr_Foreach.scala 171:152:@8220.4]
  wire  _T_617; // @[sm_x794_inr_Foreach.scala 171:240:@8222.4]
  wire  _T_618; // @[sm_x794_inr_Foreach.scala 171:259:@8223.4]
  wire  x1254_b755_D4; // @[package.scala 96:25:@8197.4 package.scala 96:25:@8198.4]
  wire  _T_621; // @[sm_x794_inr_Foreach.scala 171:295:@8225.4]
  wire  x1255_b756_D4; // @[package.scala 96:25:@8206.4 package.scala 96:25:@8207.4]
  _ _ ( // @[Math.scala 709:24:@7730.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@7742.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x1207_sub x1207_sub_1 ( // @[Math.scala 191:24:@7769.4]
    .clock(x1207_sub_1_clock),
    .reset(x1207_sub_1_reset),
    .io_a(x1207_sub_1_io_a),
    .io_b(x1207_sub_1_io_b),
    .io_flow(x1207_sub_1_io_flow),
    .io_result(x1207_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@7779.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x758_sum x758_sum_1 ( // @[Math.scala 150:24:@7788.4]
    .clock(x758_sum_1_clock),
    .reset(x758_sum_1_reset),
    .io_a(x758_sum_1_io_a),
    .io_b(x758_sum_1_io_b),
    .io_flow(x758_sum_1_io_flow),
    .io_result(x758_sum_1_io_result)
  );
  x758_sum x759_sum_1 ( // @[Math.scala 150:24:@7800.4]
    .clock(x759_sum_1_clock),
    .reset(x759_sum_1_reset),
    .io_a(x759_sum_1_io_a),
    .io_b(x759_sum_1_io_b),
    .io_flow(x759_sum_1_io_flow),
    .io_result(x759_sum_1_io_result)
  );
  x758_sum x1209_sum_1 ( // @[Math.scala 150:24:@7815.4]
    .clock(x1209_sum_1_clock),
    .reset(x1209_sum_1_reset),
    .io_a(x1209_sum_1_io_a),
    .io_b(x1209_sum_1_io_b),
    .io_flow(x1209_sum_1_io_flow),
    .io_result(x1209_sum_1_io_result)
  );
  x758_sum x763_sum_1 ( // @[Math.scala 150:24:@7847.4]
    .clock(x763_sum_1_clock),
    .reset(x763_sum_1_reset),
    .io_a(x763_sum_1_io_a),
    .io_b(x763_sum_1_io_b),
    .io_flow(x763_sum_1_io_flow),
    .io_result(x763_sum_1_io_result)
  );
  x758_sum x1212_sum_1 ( // @[Math.scala 150:24:@7862.4]
    .clock(x1212_sum_1_clock),
    .reset(x1212_sum_1_reset),
    .io_a(x1212_sum_1_io_a),
    .io_b(x1212_sum_1_io_b),
    .io_flow(x1212_sum_1_io_flow),
    .io_result(x1212_sum_1_io_result)
  );
  x758_sum x767_sum_1 ( // @[Math.scala 150:24:@7894.4]
    .clock(x767_sum_1_clock),
    .reset(x767_sum_1_reset),
    .io_a(x767_sum_1_io_a),
    .io_b(x767_sum_1_io_b),
    .io_flow(x767_sum_1_io_flow),
    .io_result(x767_sum_1_io_result)
  );
  x758_sum x1215_sum_1 ( // @[Math.scala 150:24:@7909.4]
    .clock(x1215_sum_1_clock),
    .reset(x1215_sum_1_reset),
    .io_a(x1215_sum_1_io_a),
    .io_b(x1215_sum_1_io_b),
    .io_flow(x1215_sum_1_io_flow),
    .io_result(x1215_sum_1_io_result)
  );
  x758_sum x771_sum_1 ( // @[Math.scala 150:24:@7941.4]
    .clock(x771_sum_1_clock),
    .reset(x771_sum_1_reset),
    .io_a(x771_sum_1_io_a),
    .io_b(x771_sum_1_io_b),
    .io_flow(x771_sum_1_io_flow),
    .io_result(x771_sum_1_io_result)
  );
  x758_sum x1218_sum_1 ( // @[Math.scala 150:24:@7956.4]
    .clock(x1218_sum_1_clock),
    .reset(x1218_sum_1_reset),
    .io_a(x1218_sum_1_io_a),
    .io_b(x1218_sum_1_io_b),
    .io_flow(x1218_sum_1_io_flow),
    .io_result(x1218_sum_1_io_result)
  );
  x758_sum x775_sum_1 ( // @[Math.scala 150:24:@7988.4]
    .clock(x775_sum_1_clock),
    .reset(x775_sum_1_reset),
    .io_a(x775_sum_1_io_a),
    .io_b(x775_sum_1_io_b),
    .io_flow(x775_sum_1_io_flow),
    .io_result(x775_sum_1_io_result)
  );
  x758_sum x1221_sum_1 ( // @[Math.scala 150:24:@8003.4]
    .clock(x1221_sum_1_clock),
    .reset(x1221_sum_1_reset),
    .io_a(x1221_sum_1_io_a),
    .io_b(x1221_sum_1_io_b),
    .io_flow(x1221_sum_1_io_flow),
    .io_result(x1221_sum_1_io_result)
  );
  x758_sum x779_sum_1 ( // @[Math.scala 150:24:@8035.4]
    .clock(x779_sum_1_clock),
    .reset(x779_sum_1_reset),
    .io_a(x779_sum_1_io_a),
    .io_b(x779_sum_1_io_b),
    .io_flow(x779_sum_1_io_flow),
    .io_result(x779_sum_1_io_result)
  );
  x758_sum x1224_sum_1 ( // @[Math.scala 150:24:@8050.4]
    .clock(x1224_sum_1_clock),
    .reset(x1224_sum_1_reset),
    .io_a(x1224_sum_1_io_a),
    .io_b(x1224_sum_1_io_b),
    .io_flow(x1224_sum_1_io_flow),
    .io_result(x1224_sum_1_io_result)
  );
  x758_sum x783_sum_1 ( // @[Math.scala 150:24:@8082.4]
    .clock(x783_sum_1_clock),
    .reset(x783_sum_1_reset),
    .io_a(x783_sum_1_io_a),
    .io_b(x783_sum_1_io_b),
    .io_flow(x783_sum_1_io_flow),
    .io_result(x783_sum_1_io_result)
  );
  x758_sum x1227_sum_1 ( // @[Math.scala 150:24:@8097.4]
    .clock(x1227_sum_1_clock),
    .reset(x1227_sum_1_reset),
    .io_a(x1227_sum_1_io_a),
    .io_b(x1227_sum_1_io_b),
    .io_flow(x1227_sum_1_io_flow),
    .io_result(x1227_sum_1_io_result)
  );
  x758_sum x787_sum_1 ( // @[Math.scala 150:24:@8129.4]
    .clock(x787_sum_1_clock),
    .reset(x787_sum_1_reset),
    .io_a(x787_sum_1_io_a),
    .io_b(x787_sum_1_io_b),
    .io_flow(x787_sum_1_io_flow),
    .io_result(x787_sum_1_io_result)
  );
  x758_sum x1230_sum_1 ( // @[Math.scala 150:24:@8144.4]
    .clock(x1230_sum_1_clock),
    .reset(x1230_sum_1_reset),
    .io_a(x1230_sum_1_io_a),
    .io_b(x1230_sum_1_io_b),
    .io_flow(x1230_sum_1_io_flow),
    .io_result(x1230_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@8192.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@8201.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@8212.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_328 = ~ io_in_x748_fifoinpacked_0_full; // @[sm_x794_inr_Foreach.scala 64:22:@7755.4]
  assign _T_329 = ~ io_in_x748_fifoinpacked_0_active_0_out; // @[sm_x794_inr_Foreach.scala 64:59:@7756.4]
  assign b753_number = __io_result; // @[Math.scala 712:22:@7735.4 Math.scala 713:14:@7736.4]
  assign _GEN_0 = {{11'd0}, b753_number}; // @[Math.scala 450:32:@7760.4]
  assign _T_333 = _GEN_0 << 11; // @[Math.scala 450:32:@7760.4]
  assign _GEN_1 = {{7'd0}, b753_number}; // @[Math.scala 450:32:@7765.4]
  assign _T_337 = _GEN_1 << 7; // @[Math.scala 450:32:@7765.4]
  assign x759_sum_number = x759_sum_1_io_result; // @[Math.scala 154:22:@7806.4 Math.scala 155:14:@7807.4]
  assign _GEN_2 = {{2'd0}, x759_sum_number}; // @[Math.scala 450:32:@7811.4]
  assign _T_357 = _GEN_2 << 2; // @[Math.scala 450:32:@7811.4]
  assign x763_sum_number = x763_sum_1_io_result; // @[Math.scala 154:22:@7853.4 Math.scala 155:14:@7854.4]
  assign _GEN_3 = {{2'd0}, x763_sum_number}; // @[Math.scala 450:32:@7858.4]
  assign _T_386 = _GEN_3 << 2; // @[Math.scala 450:32:@7858.4]
  assign x767_sum_number = x767_sum_1_io_result; // @[Math.scala 154:22:@7900.4 Math.scala 155:14:@7901.4]
  assign _GEN_4 = {{2'd0}, x767_sum_number}; // @[Math.scala 450:32:@7905.4]
  assign _T_415 = _GEN_4 << 2; // @[Math.scala 450:32:@7905.4]
  assign x771_sum_number = x771_sum_1_io_result; // @[Math.scala 154:22:@7947.4 Math.scala 155:14:@7948.4]
  assign _GEN_5 = {{2'd0}, x771_sum_number}; // @[Math.scala 450:32:@7952.4]
  assign _T_444 = _GEN_5 << 2; // @[Math.scala 450:32:@7952.4]
  assign x775_sum_number = x775_sum_1_io_result; // @[Math.scala 154:22:@7994.4 Math.scala 155:14:@7995.4]
  assign _GEN_6 = {{2'd0}, x775_sum_number}; // @[Math.scala 450:32:@7999.4]
  assign _T_473 = _GEN_6 << 2; // @[Math.scala 450:32:@7999.4]
  assign x779_sum_number = x779_sum_1_io_result; // @[Math.scala 154:22:@8041.4 Math.scala 155:14:@8042.4]
  assign _GEN_7 = {{2'd0}, x779_sum_number}; // @[Math.scala 450:32:@8046.4]
  assign _T_502 = _GEN_7 << 2; // @[Math.scala 450:32:@8046.4]
  assign x783_sum_number = x783_sum_1_io_result; // @[Math.scala 154:22:@8088.4 Math.scala 155:14:@8089.4]
  assign _GEN_8 = {{2'd0}, x783_sum_number}; // @[Math.scala 450:32:@8093.4]
  assign _T_531 = _GEN_8 << 2; // @[Math.scala 450:32:@8093.4]
  assign x787_sum_number = x787_sum_1_io_result; // @[Math.scala 154:22:@8135.4 Math.scala 155:14:@8136.4]
  assign _GEN_9 = {{2'd0}, x787_sum_number}; // @[Math.scala 450:32:@8140.4]
  assign _T_560 = _GEN_9 << 2; // @[Math.scala 450:32:@8140.4]
  assign _T_608 = ~ io_sigsIn_break; // @[sm_x794_inr_Foreach.scala 171:135:@8209.4]
  assign _T_612 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@8217.4 package.scala 96:25:@8218.4]
  assign _T_614 = io_rr ? _T_612 : 1'h0; // @[implicits.scala 55:10:@8219.4]
  assign _T_615 = _T_608 & _T_614; // @[sm_x794_inr_Foreach.scala 171:152:@8220.4]
  assign _T_617 = _T_615 & _T_608; // @[sm_x794_inr_Foreach.scala 171:240:@8222.4]
  assign _T_618 = _T_617 & io_sigsIn_backpressure; // @[sm_x794_inr_Foreach.scala 171:259:@8223.4]
  assign x1254_b755_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@8197.4 package.scala 96:25:@8198.4]
  assign _T_621 = _T_618 & x1254_b755_D4; // @[sm_x794_inr_Foreach.scala 171:295:@8225.4]
  assign x1255_b756_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@8206.4 package.scala 96:25:@8207.4]
  assign io_in_x748_fifoinpacked_0_wPort_0_en_0 = _T_621 & x1255_b756_D4; // @[MemInterfaceType.scala 93:57:@8229.4]
  assign io_in_x748_fifoinpacked_0_active_0_in = x1254_b755_D4 & x1255_b756_D4; // @[MemInterfaceType.scala 147:18:@8232.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@7733.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@7745.4]
  assign x1207_sub_1_clock = clock; // @[:@7770.4]
  assign x1207_sub_1_reset = reset; // @[:@7771.4]
  assign x1207_sub_1_io_a = _T_333[31:0]; // @[Math.scala 192:17:@7772.4]
  assign x1207_sub_1_io_b = _T_337[31:0]; // @[Math.scala 193:17:@7773.4]
  assign x1207_sub_1_io_flow = _T_328 | _T_329; // @[Math.scala 194:20:@7774.4]
  assign RetimeWrapper_clock = clock; // @[:@7780.4]
  assign RetimeWrapper_reset = reset; // @[:@7781.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@7783.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@7782.4]
  assign x758_sum_1_clock = clock; // @[:@7789.4]
  assign x758_sum_1_reset = reset; // @[:@7790.4]
  assign x758_sum_1_io_a = x1207_sub_1_io_result; // @[Math.scala 151:17:@7791.4]
  assign x758_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@7792.4]
  assign x758_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7793.4]
  assign x759_sum_1_clock = clock; // @[:@7801.4]
  assign x759_sum_1_reset = reset; // @[:@7802.4]
  assign x759_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@7803.4]
  assign x759_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@7804.4]
  assign x759_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7805.4]
  assign x1209_sum_1_clock = clock; // @[:@7816.4]
  assign x1209_sum_1_reset = reset; // @[:@7817.4]
  assign x1209_sum_1_io_a = _T_357[31:0]; // @[Math.scala 151:17:@7818.4]
  assign x1209_sum_1_io_b = x759_sum_1_io_result; // @[Math.scala 152:17:@7819.4]
  assign x1209_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7820.4]
  assign x763_sum_1_clock = clock; // @[:@7848.4]
  assign x763_sum_1_reset = reset; // @[:@7849.4]
  assign x763_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@7850.4]
  assign x763_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@7851.4]
  assign x763_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7852.4]
  assign x1212_sum_1_clock = clock; // @[:@7863.4]
  assign x1212_sum_1_reset = reset; // @[:@7864.4]
  assign x1212_sum_1_io_a = _T_386[31:0]; // @[Math.scala 151:17:@7865.4]
  assign x1212_sum_1_io_b = x763_sum_1_io_result; // @[Math.scala 152:17:@7866.4]
  assign x1212_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7867.4]
  assign x767_sum_1_clock = clock; // @[:@7895.4]
  assign x767_sum_1_reset = reset; // @[:@7896.4]
  assign x767_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@7897.4]
  assign x767_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@7898.4]
  assign x767_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7899.4]
  assign x1215_sum_1_clock = clock; // @[:@7910.4]
  assign x1215_sum_1_reset = reset; // @[:@7911.4]
  assign x1215_sum_1_io_a = _T_415[31:0]; // @[Math.scala 151:17:@7912.4]
  assign x1215_sum_1_io_b = x767_sum_1_io_result; // @[Math.scala 152:17:@7913.4]
  assign x1215_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7914.4]
  assign x771_sum_1_clock = clock; // @[:@7942.4]
  assign x771_sum_1_reset = reset; // @[:@7943.4]
  assign x771_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@7944.4]
  assign x771_sum_1_io_b = 32'h4; // @[Math.scala 152:17:@7945.4]
  assign x771_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7946.4]
  assign x1218_sum_1_clock = clock; // @[:@7957.4]
  assign x1218_sum_1_reset = reset; // @[:@7958.4]
  assign x1218_sum_1_io_a = _T_444[31:0]; // @[Math.scala 151:17:@7959.4]
  assign x1218_sum_1_io_b = x771_sum_1_io_result; // @[Math.scala 152:17:@7960.4]
  assign x1218_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7961.4]
  assign x775_sum_1_clock = clock; // @[:@7989.4]
  assign x775_sum_1_reset = reset; // @[:@7990.4]
  assign x775_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@7991.4]
  assign x775_sum_1_io_b = 32'h5; // @[Math.scala 152:17:@7992.4]
  assign x775_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@7993.4]
  assign x1221_sum_1_clock = clock; // @[:@8004.4]
  assign x1221_sum_1_reset = reset; // @[:@8005.4]
  assign x1221_sum_1_io_a = _T_473[31:0]; // @[Math.scala 151:17:@8006.4]
  assign x1221_sum_1_io_b = x775_sum_1_io_result; // @[Math.scala 152:17:@8007.4]
  assign x1221_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@8008.4]
  assign x779_sum_1_clock = clock; // @[:@8036.4]
  assign x779_sum_1_reset = reset; // @[:@8037.4]
  assign x779_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@8038.4]
  assign x779_sum_1_io_b = 32'h6; // @[Math.scala 152:17:@8039.4]
  assign x779_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@8040.4]
  assign x1224_sum_1_clock = clock; // @[:@8051.4]
  assign x1224_sum_1_reset = reset; // @[:@8052.4]
  assign x1224_sum_1_io_a = _T_502[31:0]; // @[Math.scala 151:17:@8053.4]
  assign x1224_sum_1_io_b = x779_sum_1_io_result; // @[Math.scala 152:17:@8054.4]
  assign x1224_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@8055.4]
  assign x783_sum_1_clock = clock; // @[:@8083.4]
  assign x783_sum_1_reset = reset; // @[:@8084.4]
  assign x783_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@8085.4]
  assign x783_sum_1_io_b = 32'h7; // @[Math.scala 152:17:@8086.4]
  assign x783_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@8087.4]
  assign x1227_sum_1_clock = clock; // @[:@8098.4]
  assign x1227_sum_1_reset = reset; // @[:@8099.4]
  assign x1227_sum_1_io_a = _T_531[31:0]; // @[Math.scala 151:17:@8100.4]
  assign x1227_sum_1_io_b = x783_sum_1_io_result; // @[Math.scala 152:17:@8101.4]
  assign x1227_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@8102.4]
  assign x787_sum_1_clock = clock; // @[:@8130.4]
  assign x787_sum_1_reset = reset; // @[:@8131.4]
  assign x787_sum_1_io_a = x758_sum_1_io_result; // @[Math.scala 151:17:@8132.4]
  assign x787_sum_1_io_b = 32'h8; // @[Math.scala 152:17:@8133.4]
  assign x787_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@8134.4]
  assign x1230_sum_1_clock = clock; // @[:@8145.4]
  assign x1230_sum_1_reset = reset; // @[:@8146.4]
  assign x1230_sum_1_io_a = _T_560[31:0]; // @[Math.scala 151:17:@8147.4]
  assign x1230_sum_1_io_b = x787_sum_1_io_result; // @[Math.scala 152:17:@8148.4]
  assign x1230_sum_1_io_flow = _T_328 | _T_329; // @[Math.scala 153:20:@8149.4]
  assign RetimeWrapper_1_clock = clock; // @[:@8193.4]
  assign RetimeWrapper_1_reset = reset; // @[:@8194.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@8196.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@8195.4]
  assign RetimeWrapper_2_clock = clock; // @[:@8202.4]
  assign RetimeWrapper_2_reset = reset; // @[:@8203.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@8205.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@8204.4]
  assign RetimeWrapper_3_clock = clock; // @[:@8213.4]
  assign RetimeWrapper_3_reset = reset; // @[:@8214.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@8216.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@8215.4]
endmodule
module RetimeWrapper_56( // @[:@9350.2]
  input   clock, // @[:@9351.4]
  input   reset, // @[:@9352.4]
  input   io_flow, // @[:@9353.4]
  input   io_in, // @[:@9353.4]
  output  io_out // @[:@9353.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@9355.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@9355.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@9355.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@9355.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@9355.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@9355.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(59)) sr ( // @[RetimeShiftRegister.scala 15:20:@9355.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@9368.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@9367.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@9366.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@9365.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@9364.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@9362.4]
endmodule
module RetimeWrapper_60( // @[:@9478.2]
  input   clock, // @[:@9479.4]
  input   reset, // @[:@9480.4]
  input   io_flow, // @[:@9481.4]
  input   io_in, // @[:@9481.4]
  output  io_out // @[:@9481.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@9483.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@9483.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@9483.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@9483.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@9483.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@9483.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(58)) sr ( // @[RetimeShiftRegister.scala 15:20:@9483.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@9496.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@9495.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@9494.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@9493.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@9492.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@9490.4]
endmodule
module x1156_inr_Foreach_SAMPLER_BOX_sm( // @[:@9498.2]
  input   clock, // @[:@9499.4]
  input   reset, // @[:@9500.4]
  input   io_enable, // @[:@9501.4]
  output  io_done, // @[:@9501.4]
  output  io_doneLatch, // @[:@9501.4]
  input   io_ctrDone, // @[:@9501.4]
  output  io_datapathEn, // @[:@9501.4]
  output  io_ctrInc, // @[:@9501.4]
  output  io_ctrRst, // @[:@9501.4]
  input   io_parentAck, // @[:@9501.4]
  input   io_backpressure, // @[:@9501.4]
  input   io_break // @[:@9501.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@9503.4]
  wire  active_reset; // @[Controllers.scala 261:22:@9503.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@9503.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@9503.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@9503.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@9503.4]
  wire  done_clock; // @[Controllers.scala 262:20:@9506.4]
  wire  done_reset; // @[Controllers.scala 262:20:@9506.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@9506.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@9506.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@9506.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@9506.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9540.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9540.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9540.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@9540.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@9540.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@9562.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@9562.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@9562.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@9562.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@9562.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@9574.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@9574.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@9574.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@9574.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@9574.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@9582.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@9582.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@9582.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@9582.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@9582.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@9598.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@9598.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@9598.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@9598.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@9598.4]
  wire  _T_80; // @[Controllers.scala 264:48:@9511.4]
  wire  _T_81; // @[Controllers.scala 264:46:@9512.4]
  wire  _T_82; // @[Controllers.scala 264:62:@9513.4]
  wire  _T_83; // @[Controllers.scala 264:60:@9514.4]
  wire  _T_100; // @[package.scala 100:49:@9531.4]
  reg  _T_103; // @[package.scala 48:56:@9532.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@9545.4 package.scala 96:25:@9546.4]
  wire  _T_110; // @[package.scala 100:49:@9547.4]
  reg  _T_113; // @[package.scala 48:56:@9548.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@9550.4]
  wire  _T_118; // @[Controllers.scala 283:41:@9555.4]
  wire  _T_119; // @[Controllers.scala 283:59:@9556.4]
  wire  _T_121; // @[Controllers.scala 284:37:@9559.4]
  wire  _T_124; // @[package.scala 96:25:@9567.4 package.scala 96:25:@9568.4]
  wire  _T_126; // @[package.scala 100:49:@9569.4]
  reg  _T_129; // @[package.scala 48:56:@9570.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@9592.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@9594.4]
  reg  _T_153; // @[package.scala 48:56:@9595.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@9603.4 package.scala 96:25:@9604.4]
  wire  _T_158; // @[Controllers.scala 292:61:@9605.4]
  wire  _T_159; // @[Controllers.scala 292:24:@9606.4]
  SRFF active ( // @[Controllers.scala 261:22:@9503.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@9506.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_56 RetimeWrapper ( // @[package.scala 93:22:@9540.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_56 RetimeWrapper_1 ( // @[package.scala 93:22:@9562.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@9574.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@9582.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_60 RetimeWrapper_4 ( // @[package.scala 93:22:@9598.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@9511.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@9512.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@9513.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@9514.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@9531.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@9545.4 package.scala 96:25:@9546.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@9547.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@9550.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@9555.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@9556.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@9559.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@9567.4 package.scala 96:25:@9568.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@9569.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@9594.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@9603.4 package.scala 96:25:@9604.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@9605.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@9606.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@9573.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@9608.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@9558.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@9561.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@9553.4]
  assign active_clock = clock; // @[:@9504.4]
  assign active_reset = reset; // @[:@9505.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@9516.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@9520.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@9521.4]
  assign done_clock = clock; // @[:@9507.4]
  assign done_reset = reset; // @[:@9508.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@9536.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@9529.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@9530.4]
  assign RetimeWrapper_clock = clock; // @[:@9541.4]
  assign RetimeWrapper_reset = reset; // @[:@9542.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@9544.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@9543.4]
  assign RetimeWrapper_1_clock = clock; // @[:@9563.4]
  assign RetimeWrapper_1_reset = reset; // @[:@9564.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@9566.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@9565.4]
  assign RetimeWrapper_2_clock = clock; // @[:@9575.4]
  assign RetimeWrapper_2_reset = reset; // @[:@9576.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@9578.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@9577.4]
  assign RetimeWrapper_3_clock = clock; // @[:@9583.4]
  assign RetimeWrapper_3_reset = reset; // @[:@9584.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@9586.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@9585.4]
  assign RetimeWrapper_4_clock = clock; // @[:@9599.4]
  assign RetimeWrapper_4_reset = reset; // @[:@9600.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@9602.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@9601.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_64( // @[:@9809.2]
  input         clock, // @[:@9810.4]
  input         reset, // @[:@9811.4]
  input         io_flow, // @[:@9812.4]
  input  [63:0] io_in, // @[:@9812.4]
  output [63:0] io_out // @[:@9812.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@9814.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@9814.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@9814.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@9814.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@9814.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@9814.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@9814.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@9827.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@9826.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@9825.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@9824.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@9823.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@9821.4]
endmodule
module SRAM_1( // @[:@9845.2]
  input        clock, // @[:@9846.4]
  input  [7:0] io_raddr, // @[:@9848.4]
  input        io_wen, // @[:@9848.4]
  input  [7:0] io_waddr, // @[:@9848.4]
  input  [7:0] io_wdata, // @[:@9848.4]
  output [7:0] io_rdata, // @[:@9848.4]
  input        io_backpressure // @[:@9848.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@9850.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@9850.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@9850.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@9850.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@9850.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@9850.4]
  wire [7:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@9850.4]
  wire [7:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@9850.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@9850.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(192), .AWIDTH(8)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@9850.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@9870.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 190:20:@9864.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@9865.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 188:18:@9862.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@9867.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@9866.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 189:20:@9863.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@9861.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@9860.4]
endmodule
module RetimeWrapper_65( // @[:@9884.2]
  input        clock, // @[:@9885.4]
  input        reset, // @[:@9886.4]
  input        io_flow, // @[:@9887.4]
  input  [7:0] io_in, // @[:@9887.4]
  output [7:0] io_out // @[:@9887.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@9889.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@9889.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@9889.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@9889.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@9889.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@9889.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@9889.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@9902.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@9901.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@9900.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@9899.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@9898.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@9896.4]
endmodule
module Mem1D_5( // @[:@9904.2]
  input        clock, // @[:@9905.4]
  input        reset, // @[:@9906.4]
  input  [7:0] io_r_ofs_0, // @[:@9907.4]
  input        io_r_backpressure, // @[:@9907.4]
  input  [7:0] io_w_ofs_0, // @[:@9907.4]
  input  [7:0] io_w_data_0, // @[:@9907.4]
  input        io_w_en_0, // @[:@9907.4]
  output [7:0] io_output // @[:@9907.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@9911.4]
  wire [7:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@9911.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 705:21:@9911.4]
  wire [7:0] SRAM_io_waddr; // @[MemPrimitives.scala 705:21:@9911.4]
  wire [7:0] SRAM_io_wdata; // @[MemPrimitives.scala 705:21:@9911.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@9911.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@9911.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9914.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9914.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9914.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@9914.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@9914.4]
  wire  wInBound; // @[MemPrimitives.scala 692:32:@9909.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 705:21:@9911.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_65 RetimeWrapper ( // @[package.scala 93:22:@9914.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 8'hc0; // @[MemPrimitives.scala 692:32:@9909.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@9927.4]
  assign SRAM_clock = clock; // @[:@9912.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@9921.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 709:22:@9924.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 708:22:@9922.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 710:22:@9925.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@9926.4]
  assign RetimeWrapper_clock = clock; // @[:@9915.4]
  assign RetimeWrapper_reset = reset; // @[:@9916.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@9918.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@9917.4]
endmodule
module StickySelects_1( // @[:@13829.2]
  input   clock, // @[:@13830.4]
  input   reset, // @[:@13831.4]
  input   io_ins_0, // @[:@13832.4]
  input   io_ins_1, // @[:@13832.4]
  input   io_ins_2, // @[:@13832.4]
  input   io_ins_3, // @[:@13832.4]
  input   io_ins_4, // @[:@13832.4]
  input   io_ins_5, // @[:@13832.4]
  input   io_ins_6, // @[:@13832.4]
  input   io_ins_7, // @[:@13832.4]
  input   io_ins_8, // @[:@13832.4]
  input   io_ins_9, // @[:@13832.4]
  input   io_ins_10, // @[:@13832.4]
  input   io_ins_11, // @[:@13832.4]
  input   io_ins_12, // @[:@13832.4]
  input   io_ins_13, // @[:@13832.4]
  input   io_ins_14, // @[:@13832.4]
  output  io_outs_0, // @[:@13832.4]
  output  io_outs_1, // @[:@13832.4]
  output  io_outs_2, // @[:@13832.4]
  output  io_outs_3, // @[:@13832.4]
  output  io_outs_4, // @[:@13832.4]
  output  io_outs_5, // @[:@13832.4]
  output  io_outs_6, // @[:@13832.4]
  output  io_outs_7, // @[:@13832.4]
  output  io_outs_8, // @[:@13832.4]
  output  io_outs_9, // @[:@13832.4]
  output  io_outs_10, // @[:@13832.4]
  output  io_outs_11, // @[:@13832.4]
  output  io_outs_12, // @[:@13832.4]
  output  io_outs_13, // @[:@13832.4]
  output  io_outs_14 // @[:@13832.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@13834.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@13835.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@13836.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@13837.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@13838.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@13839.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@13840.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@13841.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@13842.4]
  reg [31:0] _RAND_8;
  reg  _T_46; // @[StickySelects.scala 37:46:@13843.4]
  reg [31:0] _RAND_9;
  reg  _T_49; // @[StickySelects.scala 37:46:@13844.4]
  reg [31:0] _RAND_10;
  reg  _T_52; // @[StickySelects.scala 37:46:@13845.4]
  reg [31:0] _RAND_11;
  reg  _T_55; // @[StickySelects.scala 37:46:@13846.4]
  reg [31:0] _RAND_12;
  reg  _T_58; // @[StickySelects.scala 37:46:@13847.4]
  reg [31:0] _RAND_13;
  reg  _T_61; // @[StickySelects.scala 37:46:@13848.4]
  reg [31:0] _RAND_14;
  wire  _T_62; // @[StickySelects.scala 47:46:@13849.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@13850.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@13851.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@13852.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@13853.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@13854.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@13855.4]
  wire  _T_69; // @[StickySelects.scala 47:46:@13856.4]
  wire  _T_70; // @[StickySelects.scala 47:46:@13857.4]
  wire  _T_71; // @[StickySelects.scala 47:46:@13858.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@13859.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@13860.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@13861.4]
  wire  _T_75; // @[StickySelects.scala 49:53:@13862.4]
  wire  _T_76; // @[StickySelects.scala 49:21:@13863.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@13865.4]
  wire  _T_78; // @[StickySelects.scala 47:46:@13866.4]
  wire  _T_79; // @[StickySelects.scala 47:46:@13867.4]
  wire  _T_80; // @[StickySelects.scala 47:46:@13868.4]
  wire  _T_81; // @[StickySelects.scala 47:46:@13869.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@13870.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@13871.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@13872.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@13873.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@13874.4]
  wire  _T_87; // @[StickySelects.scala 47:46:@13875.4]
  wire  _T_88; // @[StickySelects.scala 47:46:@13876.4]
  wire  _T_89; // @[StickySelects.scala 47:46:@13877.4]
  wire  _T_90; // @[StickySelects.scala 49:53:@13878.4]
  wire  _T_91; // @[StickySelects.scala 49:21:@13879.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@13881.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@13882.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@13883.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@13884.4]
  wire  _T_96; // @[StickySelects.scala 47:46:@13885.4]
  wire  _T_97; // @[StickySelects.scala 47:46:@13886.4]
  wire  _T_98; // @[StickySelects.scala 47:46:@13887.4]
  wire  _T_99; // @[StickySelects.scala 47:46:@13888.4]
  wire  _T_100; // @[StickySelects.scala 47:46:@13889.4]
  wire  _T_101; // @[StickySelects.scala 47:46:@13890.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@13891.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@13892.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@13893.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@13894.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@13895.4]
  wire  _T_108; // @[StickySelects.scala 47:46:@13898.4]
  wire  _T_109; // @[StickySelects.scala 47:46:@13899.4]
  wire  _T_110; // @[StickySelects.scala 47:46:@13900.4]
  wire  _T_111; // @[StickySelects.scala 47:46:@13901.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@13902.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@13903.4]
  wire  _T_114; // @[StickySelects.scala 47:46:@13904.4]
  wire  _T_115; // @[StickySelects.scala 47:46:@13905.4]
  wire  _T_116; // @[StickySelects.scala 47:46:@13906.4]
  wire  _T_117; // @[StickySelects.scala 47:46:@13907.4]
  wire  _T_118; // @[StickySelects.scala 47:46:@13908.4]
  wire  _T_119; // @[StickySelects.scala 47:46:@13909.4]
  wire  _T_120; // @[StickySelects.scala 49:53:@13910.4]
  wire  _T_121; // @[StickySelects.scala 49:21:@13911.4]
  wire  _T_124; // @[StickySelects.scala 47:46:@13915.4]
  wire  _T_125; // @[StickySelects.scala 47:46:@13916.4]
  wire  _T_126; // @[StickySelects.scala 47:46:@13917.4]
  wire  _T_127; // @[StickySelects.scala 47:46:@13918.4]
  wire  _T_128; // @[StickySelects.scala 47:46:@13919.4]
  wire  _T_129; // @[StickySelects.scala 47:46:@13920.4]
  wire  _T_130; // @[StickySelects.scala 47:46:@13921.4]
  wire  _T_131; // @[StickySelects.scala 47:46:@13922.4]
  wire  _T_132; // @[StickySelects.scala 47:46:@13923.4]
  wire  _T_133; // @[StickySelects.scala 47:46:@13924.4]
  wire  _T_134; // @[StickySelects.scala 47:46:@13925.4]
  wire  _T_135; // @[StickySelects.scala 49:53:@13926.4]
  wire  _T_136; // @[StickySelects.scala 49:21:@13927.4]
  wire  _T_140; // @[StickySelects.scala 47:46:@13932.4]
  wire  _T_141; // @[StickySelects.scala 47:46:@13933.4]
  wire  _T_142; // @[StickySelects.scala 47:46:@13934.4]
  wire  _T_143; // @[StickySelects.scala 47:46:@13935.4]
  wire  _T_144; // @[StickySelects.scala 47:46:@13936.4]
  wire  _T_145; // @[StickySelects.scala 47:46:@13937.4]
  wire  _T_146; // @[StickySelects.scala 47:46:@13938.4]
  wire  _T_147; // @[StickySelects.scala 47:46:@13939.4]
  wire  _T_148; // @[StickySelects.scala 47:46:@13940.4]
  wire  _T_149; // @[StickySelects.scala 47:46:@13941.4]
  wire  _T_150; // @[StickySelects.scala 49:53:@13942.4]
  wire  _T_151; // @[StickySelects.scala 49:21:@13943.4]
  wire  _T_156; // @[StickySelects.scala 47:46:@13949.4]
  wire  _T_157; // @[StickySelects.scala 47:46:@13950.4]
  wire  _T_158; // @[StickySelects.scala 47:46:@13951.4]
  wire  _T_159; // @[StickySelects.scala 47:46:@13952.4]
  wire  _T_160; // @[StickySelects.scala 47:46:@13953.4]
  wire  _T_161; // @[StickySelects.scala 47:46:@13954.4]
  wire  _T_162; // @[StickySelects.scala 47:46:@13955.4]
  wire  _T_163; // @[StickySelects.scala 47:46:@13956.4]
  wire  _T_164; // @[StickySelects.scala 47:46:@13957.4]
  wire  _T_165; // @[StickySelects.scala 49:53:@13958.4]
  wire  _T_166; // @[StickySelects.scala 49:21:@13959.4]
  wire  _T_172; // @[StickySelects.scala 47:46:@13966.4]
  wire  _T_173; // @[StickySelects.scala 47:46:@13967.4]
  wire  _T_174; // @[StickySelects.scala 47:46:@13968.4]
  wire  _T_175; // @[StickySelects.scala 47:46:@13969.4]
  wire  _T_176; // @[StickySelects.scala 47:46:@13970.4]
  wire  _T_177; // @[StickySelects.scala 47:46:@13971.4]
  wire  _T_178; // @[StickySelects.scala 47:46:@13972.4]
  wire  _T_179; // @[StickySelects.scala 47:46:@13973.4]
  wire  _T_180; // @[StickySelects.scala 49:53:@13974.4]
  wire  _T_181; // @[StickySelects.scala 49:21:@13975.4]
  wire  _T_188; // @[StickySelects.scala 47:46:@13983.4]
  wire  _T_189; // @[StickySelects.scala 47:46:@13984.4]
  wire  _T_190; // @[StickySelects.scala 47:46:@13985.4]
  wire  _T_191; // @[StickySelects.scala 47:46:@13986.4]
  wire  _T_192; // @[StickySelects.scala 47:46:@13987.4]
  wire  _T_193; // @[StickySelects.scala 47:46:@13988.4]
  wire  _T_194; // @[StickySelects.scala 47:46:@13989.4]
  wire  _T_195; // @[StickySelects.scala 49:53:@13990.4]
  wire  _T_196; // @[StickySelects.scala 49:21:@13991.4]
  wire  _T_204; // @[StickySelects.scala 47:46:@14000.4]
  wire  _T_205; // @[StickySelects.scala 47:46:@14001.4]
  wire  _T_206; // @[StickySelects.scala 47:46:@14002.4]
  wire  _T_207; // @[StickySelects.scala 47:46:@14003.4]
  wire  _T_208; // @[StickySelects.scala 47:46:@14004.4]
  wire  _T_209; // @[StickySelects.scala 47:46:@14005.4]
  wire  _T_210; // @[StickySelects.scala 49:53:@14006.4]
  wire  _T_211; // @[StickySelects.scala 49:21:@14007.4]
  wire  _T_220; // @[StickySelects.scala 47:46:@14017.4]
  wire  _T_221; // @[StickySelects.scala 47:46:@14018.4]
  wire  _T_222; // @[StickySelects.scala 47:46:@14019.4]
  wire  _T_223; // @[StickySelects.scala 47:46:@14020.4]
  wire  _T_224; // @[StickySelects.scala 47:46:@14021.4]
  wire  _T_225; // @[StickySelects.scala 49:53:@14022.4]
  wire  _T_226; // @[StickySelects.scala 49:21:@14023.4]
  wire  _T_236; // @[StickySelects.scala 47:46:@14034.4]
  wire  _T_237; // @[StickySelects.scala 47:46:@14035.4]
  wire  _T_238; // @[StickySelects.scala 47:46:@14036.4]
  wire  _T_239; // @[StickySelects.scala 47:46:@14037.4]
  wire  _T_240; // @[StickySelects.scala 49:53:@14038.4]
  wire  _T_241; // @[StickySelects.scala 49:21:@14039.4]
  wire  _T_252; // @[StickySelects.scala 47:46:@14051.4]
  wire  _T_253; // @[StickySelects.scala 47:46:@14052.4]
  wire  _T_254; // @[StickySelects.scala 47:46:@14053.4]
  wire  _T_255; // @[StickySelects.scala 49:53:@14054.4]
  wire  _T_256; // @[StickySelects.scala 49:21:@14055.4]
  wire  _T_268; // @[StickySelects.scala 47:46:@14068.4]
  wire  _T_269; // @[StickySelects.scala 47:46:@14069.4]
  wire  _T_270; // @[StickySelects.scala 49:53:@14070.4]
  wire  _T_271; // @[StickySelects.scala 49:21:@14071.4]
  wire  _T_284; // @[StickySelects.scala 47:46:@14085.4]
  wire  _T_285; // @[StickySelects.scala 49:53:@14086.4]
  wire  _T_286; // @[StickySelects.scala 49:21:@14087.4]
  assign _T_62 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@13849.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@13850.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@13851.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@13852.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@13853.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@13854.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@13855.4]
  assign _T_69 = _T_68 | io_ins_9; // @[StickySelects.scala 47:46:@13856.4]
  assign _T_70 = _T_69 | io_ins_10; // @[StickySelects.scala 47:46:@13857.4]
  assign _T_71 = _T_70 | io_ins_11; // @[StickySelects.scala 47:46:@13858.4]
  assign _T_72 = _T_71 | io_ins_12; // @[StickySelects.scala 47:46:@13859.4]
  assign _T_73 = _T_72 | io_ins_13; // @[StickySelects.scala 47:46:@13860.4]
  assign _T_74 = _T_73 | io_ins_14; // @[StickySelects.scala 47:46:@13861.4]
  assign _T_75 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@13862.4]
  assign _T_76 = _T_74 ? io_ins_0 : _T_75; // @[StickySelects.scala 49:21:@13863.4]
  assign _T_77 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@13865.4]
  assign _T_78 = _T_77 | io_ins_3; // @[StickySelects.scala 47:46:@13866.4]
  assign _T_79 = _T_78 | io_ins_4; // @[StickySelects.scala 47:46:@13867.4]
  assign _T_80 = _T_79 | io_ins_5; // @[StickySelects.scala 47:46:@13868.4]
  assign _T_81 = _T_80 | io_ins_6; // @[StickySelects.scala 47:46:@13869.4]
  assign _T_82 = _T_81 | io_ins_7; // @[StickySelects.scala 47:46:@13870.4]
  assign _T_83 = _T_82 | io_ins_8; // @[StickySelects.scala 47:46:@13871.4]
  assign _T_84 = _T_83 | io_ins_9; // @[StickySelects.scala 47:46:@13872.4]
  assign _T_85 = _T_84 | io_ins_10; // @[StickySelects.scala 47:46:@13873.4]
  assign _T_86 = _T_85 | io_ins_11; // @[StickySelects.scala 47:46:@13874.4]
  assign _T_87 = _T_86 | io_ins_12; // @[StickySelects.scala 47:46:@13875.4]
  assign _T_88 = _T_87 | io_ins_13; // @[StickySelects.scala 47:46:@13876.4]
  assign _T_89 = _T_88 | io_ins_14; // @[StickySelects.scala 47:46:@13877.4]
  assign _T_90 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@13878.4]
  assign _T_91 = _T_89 ? io_ins_1 : _T_90; // @[StickySelects.scala 49:21:@13879.4]
  assign _T_92 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@13881.4]
  assign _T_93 = _T_92 | io_ins_3; // @[StickySelects.scala 47:46:@13882.4]
  assign _T_94 = _T_93 | io_ins_4; // @[StickySelects.scala 47:46:@13883.4]
  assign _T_95 = _T_94 | io_ins_5; // @[StickySelects.scala 47:46:@13884.4]
  assign _T_96 = _T_95 | io_ins_6; // @[StickySelects.scala 47:46:@13885.4]
  assign _T_97 = _T_96 | io_ins_7; // @[StickySelects.scala 47:46:@13886.4]
  assign _T_98 = _T_97 | io_ins_8; // @[StickySelects.scala 47:46:@13887.4]
  assign _T_99 = _T_98 | io_ins_9; // @[StickySelects.scala 47:46:@13888.4]
  assign _T_100 = _T_99 | io_ins_10; // @[StickySelects.scala 47:46:@13889.4]
  assign _T_101 = _T_100 | io_ins_11; // @[StickySelects.scala 47:46:@13890.4]
  assign _T_102 = _T_101 | io_ins_12; // @[StickySelects.scala 47:46:@13891.4]
  assign _T_103 = _T_102 | io_ins_13; // @[StickySelects.scala 47:46:@13892.4]
  assign _T_104 = _T_103 | io_ins_14; // @[StickySelects.scala 47:46:@13893.4]
  assign _T_105 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@13894.4]
  assign _T_106 = _T_104 ? io_ins_2 : _T_105; // @[StickySelects.scala 49:21:@13895.4]
  assign _T_108 = _T_92 | io_ins_2; // @[StickySelects.scala 47:46:@13898.4]
  assign _T_109 = _T_108 | io_ins_4; // @[StickySelects.scala 47:46:@13899.4]
  assign _T_110 = _T_109 | io_ins_5; // @[StickySelects.scala 47:46:@13900.4]
  assign _T_111 = _T_110 | io_ins_6; // @[StickySelects.scala 47:46:@13901.4]
  assign _T_112 = _T_111 | io_ins_7; // @[StickySelects.scala 47:46:@13902.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@13903.4]
  assign _T_114 = _T_113 | io_ins_9; // @[StickySelects.scala 47:46:@13904.4]
  assign _T_115 = _T_114 | io_ins_10; // @[StickySelects.scala 47:46:@13905.4]
  assign _T_116 = _T_115 | io_ins_11; // @[StickySelects.scala 47:46:@13906.4]
  assign _T_117 = _T_116 | io_ins_12; // @[StickySelects.scala 47:46:@13907.4]
  assign _T_118 = _T_117 | io_ins_13; // @[StickySelects.scala 47:46:@13908.4]
  assign _T_119 = _T_118 | io_ins_14; // @[StickySelects.scala 47:46:@13909.4]
  assign _T_120 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@13910.4]
  assign _T_121 = _T_119 ? io_ins_3 : _T_120; // @[StickySelects.scala 49:21:@13911.4]
  assign _T_124 = _T_108 | io_ins_3; // @[StickySelects.scala 47:46:@13915.4]
  assign _T_125 = _T_124 | io_ins_5; // @[StickySelects.scala 47:46:@13916.4]
  assign _T_126 = _T_125 | io_ins_6; // @[StickySelects.scala 47:46:@13917.4]
  assign _T_127 = _T_126 | io_ins_7; // @[StickySelects.scala 47:46:@13918.4]
  assign _T_128 = _T_127 | io_ins_8; // @[StickySelects.scala 47:46:@13919.4]
  assign _T_129 = _T_128 | io_ins_9; // @[StickySelects.scala 47:46:@13920.4]
  assign _T_130 = _T_129 | io_ins_10; // @[StickySelects.scala 47:46:@13921.4]
  assign _T_131 = _T_130 | io_ins_11; // @[StickySelects.scala 47:46:@13922.4]
  assign _T_132 = _T_131 | io_ins_12; // @[StickySelects.scala 47:46:@13923.4]
  assign _T_133 = _T_132 | io_ins_13; // @[StickySelects.scala 47:46:@13924.4]
  assign _T_134 = _T_133 | io_ins_14; // @[StickySelects.scala 47:46:@13925.4]
  assign _T_135 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@13926.4]
  assign _T_136 = _T_134 ? io_ins_4 : _T_135; // @[StickySelects.scala 49:21:@13927.4]
  assign _T_140 = _T_124 | io_ins_4; // @[StickySelects.scala 47:46:@13932.4]
  assign _T_141 = _T_140 | io_ins_6; // @[StickySelects.scala 47:46:@13933.4]
  assign _T_142 = _T_141 | io_ins_7; // @[StickySelects.scala 47:46:@13934.4]
  assign _T_143 = _T_142 | io_ins_8; // @[StickySelects.scala 47:46:@13935.4]
  assign _T_144 = _T_143 | io_ins_9; // @[StickySelects.scala 47:46:@13936.4]
  assign _T_145 = _T_144 | io_ins_10; // @[StickySelects.scala 47:46:@13937.4]
  assign _T_146 = _T_145 | io_ins_11; // @[StickySelects.scala 47:46:@13938.4]
  assign _T_147 = _T_146 | io_ins_12; // @[StickySelects.scala 47:46:@13939.4]
  assign _T_148 = _T_147 | io_ins_13; // @[StickySelects.scala 47:46:@13940.4]
  assign _T_149 = _T_148 | io_ins_14; // @[StickySelects.scala 47:46:@13941.4]
  assign _T_150 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@13942.4]
  assign _T_151 = _T_149 ? io_ins_5 : _T_150; // @[StickySelects.scala 49:21:@13943.4]
  assign _T_156 = _T_140 | io_ins_5; // @[StickySelects.scala 47:46:@13949.4]
  assign _T_157 = _T_156 | io_ins_7; // @[StickySelects.scala 47:46:@13950.4]
  assign _T_158 = _T_157 | io_ins_8; // @[StickySelects.scala 47:46:@13951.4]
  assign _T_159 = _T_158 | io_ins_9; // @[StickySelects.scala 47:46:@13952.4]
  assign _T_160 = _T_159 | io_ins_10; // @[StickySelects.scala 47:46:@13953.4]
  assign _T_161 = _T_160 | io_ins_11; // @[StickySelects.scala 47:46:@13954.4]
  assign _T_162 = _T_161 | io_ins_12; // @[StickySelects.scala 47:46:@13955.4]
  assign _T_163 = _T_162 | io_ins_13; // @[StickySelects.scala 47:46:@13956.4]
  assign _T_164 = _T_163 | io_ins_14; // @[StickySelects.scala 47:46:@13957.4]
  assign _T_165 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@13958.4]
  assign _T_166 = _T_164 ? io_ins_6 : _T_165; // @[StickySelects.scala 49:21:@13959.4]
  assign _T_172 = _T_156 | io_ins_6; // @[StickySelects.scala 47:46:@13966.4]
  assign _T_173 = _T_172 | io_ins_8; // @[StickySelects.scala 47:46:@13967.4]
  assign _T_174 = _T_173 | io_ins_9; // @[StickySelects.scala 47:46:@13968.4]
  assign _T_175 = _T_174 | io_ins_10; // @[StickySelects.scala 47:46:@13969.4]
  assign _T_176 = _T_175 | io_ins_11; // @[StickySelects.scala 47:46:@13970.4]
  assign _T_177 = _T_176 | io_ins_12; // @[StickySelects.scala 47:46:@13971.4]
  assign _T_178 = _T_177 | io_ins_13; // @[StickySelects.scala 47:46:@13972.4]
  assign _T_179 = _T_178 | io_ins_14; // @[StickySelects.scala 47:46:@13973.4]
  assign _T_180 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@13974.4]
  assign _T_181 = _T_179 ? io_ins_7 : _T_180; // @[StickySelects.scala 49:21:@13975.4]
  assign _T_188 = _T_172 | io_ins_7; // @[StickySelects.scala 47:46:@13983.4]
  assign _T_189 = _T_188 | io_ins_9; // @[StickySelects.scala 47:46:@13984.4]
  assign _T_190 = _T_189 | io_ins_10; // @[StickySelects.scala 47:46:@13985.4]
  assign _T_191 = _T_190 | io_ins_11; // @[StickySelects.scala 47:46:@13986.4]
  assign _T_192 = _T_191 | io_ins_12; // @[StickySelects.scala 47:46:@13987.4]
  assign _T_193 = _T_192 | io_ins_13; // @[StickySelects.scala 47:46:@13988.4]
  assign _T_194 = _T_193 | io_ins_14; // @[StickySelects.scala 47:46:@13989.4]
  assign _T_195 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@13990.4]
  assign _T_196 = _T_194 ? io_ins_8 : _T_195; // @[StickySelects.scala 49:21:@13991.4]
  assign _T_204 = _T_188 | io_ins_8; // @[StickySelects.scala 47:46:@14000.4]
  assign _T_205 = _T_204 | io_ins_10; // @[StickySelects.scala 47:46:@14001.4]
  assign _T_206 = _T_205 | io_ins_11; // @[StickySelects.scala 47:46:@14002.4]
  assign _T_207 = _T_206 | io_ins_12; // @[StickySelects.scala 47:46:@14003.4]
  assign _T_208 = _T_207 | io_ins_13; // @[StickySelects.scala 47:46:@14004.4]
  assign _T_209 = _T_208 | io_ins_14; // @[StickySelects.scala 47:46:@14005.4]
  assign _T_210 = io_ins_9 | _T_46; // @[StickySelects.scala 49:53:@14006.4]
  assign _T_211 = _T_209 ? io_ins_9 : _T_210; // @[StickySelects.scala 49:21:@14007.4]
  assign _T_220 = _T_204 | io_ins_9; // @[StickySelects.scala 47:46:@14017.4]
  assign _T_221 = _T_220 | io_ins_11; // @[StickySelects.scala 47:46:@14018.4]
  assign _T_222 = _T_221 | io_ins_12; // @[StickySelects.scala 47:46:@14019.4]
  assign _T_223 = _T_222 | io_ins_13; // @[StickySelects.scala 47:46:@14020.4]
  assign _T_224 = _T_223 | io_ins_14; // @[StickySelects.scala 47:46:@14021.4]
  assign _T_225 = io_ins_10 | _T_49; // @[StickySelects.scala 49:53:@14022.4]
  assign _T_226 = _T_224 ? io_ins_10 : _T_225; // @[StickySelects.scala 49:21:@14023.4]
  assign _T_236 = _T_220 | io_ins_10; // @[StickySelects.scala 47:46:@14034.4]
  assign _T_237 = _T_236 | io_ins_12; // @[StickySelects.scala 47:46:@14035.4]
  assign _T_238 = _T_237 | io_ins_13; // @[StickySelects.scala 47:46:@14036.4]
  assign _T_239 = _T_238 | io_ins_14; // @[StickySelects.scala 47:46:@14037.4]
  assign _T_240 = io_ins_11 | _T_52; // @[StickySelects.scala 49:53:@14038.4]
  assign _T_241 = _T_239 ? io_ins_11 : _T_240; // @[StickySelects.scala 49:21:@14039.4]
  assign _T_252 = _T_236 | io_ins_11; // @[StickySelects.scala 47:46:@14051.4]
  assign _T_253 = _T_252 | io_ins_13; // @[StickySelects.scala 47:46:@14052.4]
  assign _T_254 = _T_253 | io_ins_14; // @[StickySelects.scala 47:46:@14053.4]
  assign _T_255 = io_ins_12 | _T_55; // @[StickySelects.scala 49:53:@14054.4]
  assign _T_256 = _T_254 ? io_ins_12 : _T_255; // @[StickySelects.scala 49:21:@14055.4]
  assign _T_268 = _T_252 | io_ins_12; // @[StickySelects.scala 47:46:@14068.4]
  assign _T_269 = _T_268 | io_ins_14; // @[StickySelects.scala 47:46:@14069.4]
  assign _T_270 = io_ins_13 | _T_58; // @[StickySelects.scala 49:53:@14070.4]
  assign _T_271 = _T_269 ? io_ins_13 : _T_270; // @[StickySelects.scala 49:21:@14071.4]
  assign _T_284 = _T_268 | io_ins_13; // @[StickySelects.scala 47:46:@14085.4]
  assign _T_285 = io_ins_14 | _T_61; // @[StickySelects.scala 49:53:@14086.4]
  assign _T_286 = _T_284 ? io_ins_14 : _T_285; // @[StickySelects.scala 49:21:@14087.4]
  assign io_outs_0 = _T_74 ? io_ins_0 : _T_75; // @[StickySelects.scala 53:57:@14089.4]
  assign io_outs_1 = _T_89 ? io_ins_1 : _T_90; // @[StickySelects.scala 53:57:@14090.4]
  assign io_outs_2 = _T_104 ? io_ins_2 : _T_105; // @[StickySelects.scala 53:57:@14091.4]
  assign io_outs_3 = _T_119 ? io_ins_3 : _T_120; // @[StickySelects.scala 53:57:@14092.4]
  assign io_outs_4 = _T_134 ? io_ins_4 : _T_135; // @[StickySelects.scala 53:57:@14093.4]
  assign io_outs_5 = _T_149 ? io_ins_5 : _T_150; // @[StickySelects.scala 53:57:@14094.4]
  assign io_outs_6 = _T_164 ? io_ins_6 : _T_165; // @[StickySelects.scala 53:57:@14095.4]
  assign io_outs_7 = _T_179 ? io_ins_7 : _T_180; // @[StickySelects.scala 53:57:@14096.4]
  assign io_outs_8 = _T_194 ? io_ins_8 : _T_195; // @[StickySelects.scala 53:57:@14097.4]
  assign io_outs_9 = _T_209 ? io_ins_9 : _T_210; // @[StickySelects.scala 53:57:@14098.4]
  assign io_outs_10 = _T_224 ? io_ins_10 : _T_225; // @[StickySelects.scala 53:57:@14099.4]
  assign io_outs_11 = _T_239 ? io_ins_11 : _T_240; // @[StickySelects.scala 53:57:@14100.4]
  assign io_outs_12 = _T_254 ? io_ins_12 : _T_255; // @[StickySelects.scala 53:57:@14101.4]
  assign io_outs_13 = _T_269 ? io_ins_13 : _T_270; // @[StickySelects.scala 53:57:@14102.4]
  assign io_outs_14 = _T_284 ? io_ins_14 : _T_285; // @[StickySelects.scala 53:57:@14103.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_46 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_49 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_52 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_55 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_58 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_61 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_74) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_75;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_89) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_90;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_105;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_119) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_120;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_134) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_135;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_149) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_150;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_164) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_165;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_179) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_180;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_194) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_195;
      end
    end
    if (reset) begin
      _T_46 <= 1'h0;
    end else begin
      if (_T_209) begin
        _T_46 <= io_ins_9;
      end else begin
        _T_46 <= _T_210;
      end
    end
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_224) begin
        _T_49 <= io_ins_10;
      end else begin
        _T_49 <= _T_225;
      end
    end
    if (reset) begin
      _T_52 <= 1'h0;
    end else begin
      if (_T_239) begin
        _T_52 <= io_ins_11;
      end else begin
        _T_52 <= _T_240;
      end
    end
    if (reset) begin
      _T_55 <= 1'h0;
    end else begin
      if (_T_254) begin
        _T_55 <= io_ins_12;
      end else begin
        _T_55 <= _T_255;
      end
    end
    if (reset) begin
      _T_58 <= 1'h0;
    end else begin
      if (_T_269) begin
        _T_58 <= io_ins_13;
      end else begin
        _T_58 <= _T_270;
      end
    end
    if (reset) begin
      _T_61 <= 1'h0;
    end else begin
      if (_T_284) begin
        _T_61 <= io_ins_14;
      end else begin
        _T_61 <= _T_285;
      end
    end
  end
endmodule
module x805_lb_0( // @[:@44069.2]
  input        clock, // @[:@44070.4]
  input        reset, // @[:@44071.4]
  input  [3:0] io_rPort_29_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_29_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_29_ofs_0, // @[:@44072.4]
  input        io_rPort_29_en_0, // @[:@44072.4]
  input        io_rPort_29_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_29_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_28_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_28_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_28_ofs_0, // @[:@44072.4]
  input        io_rPort_28_en_0, // @[:@44072.4]
  input        io_rPort_28_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_28_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_27_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_27_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_27_ofs_0, // @[:@44072.4]
  input        io_rPort_27_en_0, // @[:@44072.4]
  input        io_rPort_27_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_27_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_26_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_26_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_26_ofs_0, // @[:@44072.4]
  input        io_rPort_26_en_0, // @[:@44072.4]
  input        io_rPort_26_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_26_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_25_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_25_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_25_ofs_0, // @[:@44072.4]
  input        io_rPort_25_en_0, // @[:@44072.4]
  input        io_rPort_25_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_25_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_24_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_24_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_24_ofs_0, // @[:@44072.4]
  input        io_rPort_24_en_0, // @[:@44072.4]
  input        io_rPort_24_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_24_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_23_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_23_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_23_ofs_0, // @[:@44072.4]
  input        io_rPort_23_en_0, // @[:@44072.4]
  input        io_rPort_23_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_23_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_22_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_22_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_22_ofs_0, // @[:@44072.4]
  input        io_rPort_22_en_0, // @[:@44072.4]
  input        io_rPort_22_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_22_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_21_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_21_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_21_ofs_0, // @[:@44072.4]
  input        io_rPort_21_en_0, // @[:@44072.4]
  input        io_rPort_21_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_21_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_20_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_20_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_20_ofs_0, // @[:@44072.4]
  input        io_rPort_20_en_0, // @[:@44072.4]
  input        io_rPort_20_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_20_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_19_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_19_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_19_ofs_0, // @[:@44072.4]
  input        io_rPort_19_en_0, // @[:@44072.4]
  input        io_rPort_19_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_19_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_18_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_18_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_18_ofs_0, // @[:@44072.4]
  input        io_rPort_18_en_0, // @[:@44072.4]
  input        io_rPort_18_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_18_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_17_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_17_ofs_0, // @[:@44072.4]
  input        io_rPort_17_en_0, // @[:@44072.4]
  input        io_rPort_17_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_17_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_16_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_16_ofs_0, // @[:@44072.4]
  input        io_rPort_16_en_0, // @[:@44072.4]
  input        io_rPort_16_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_16_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_15_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_15_ofs_0, // @[:@44072.4]
  input        io_rPort_15_en_0, // @[:@44072.4]
  input        io_rPort_15_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_15_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_14_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_14_ofs_0, // @[:@44072.4]
  input        io_rPort_14_en_0, // @[:@44072.4]
  input        io_rPort_14_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_14_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_13_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_13_ofs_0, // @[:@44072.4]
  input        io_rPort_13_en_0, // @[:@44072.4]
  input        io_rPort_13_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_13_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_12_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_12_ofs_0, // @[:@44072.4]
  input        io_rPort_12_en_0, // @[:@44072.4]
  input        io_rPort_12_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_12_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_11_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_11_ofs_0, // @[:@44072.4]
  input        io_rPort_11_en_0, // @[:@44072.4]
  input        io_rPort_11_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_11_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_10_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_10_ofs_0, // @[:@44072.4]
  input        io_rPort_10_en_0, // @[:@44072.4]
  input        io_rPort_10_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_10_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_9_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_9_ofs_0, // @[:@44072.4]
  input        io_rPort_9_en_0, // @[:@44072.4]
  input        io_rPort_9_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_9_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_8_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_8_ofs_0, // @[:@44072.4]
  input        io_rPort_8_en_0, // @[:@44072.4]
  input        io_rPort_8_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_8_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_7_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_7_ofs_0, // @[:@44072.4]
  input        io_rPort_7_en_0, // @[:@44072.4]
  input        io_rPort_7_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_7_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_6_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_6_ofs_0, // @[:@44072.4]
  input        io_rPort_6_en_0, // @[:@44072.4]
  input        io_rPort_6_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_6_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_5_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_5_ofs_0, // @[:@44072.4]
  input        io_rPort_5_en_0, // @[:@44072.4]
  input        io_rPort_5_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_5_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_4_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_4_ofs_0, // @[:@44072.4]
  input        io_rPort_4_en_0, // @[:@44072.4]
  input        io_rPort_4_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_4_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_3_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_3_ofs_0, // @[:@44072.4]
  input        io_rPort_3_en_0, // @[:@44072.4]
  input        io_rPort_3_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_3_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_2_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_2_ofs_0, // @[:@44072.4]
  input        io_rPort_2_en_0, // @[:@44072.4]
  input        io_rPort_2_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_2_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_1_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_1_ofs_0, // @[:@44072.4]
  input        io_rPort_1_en_0, // @[:@44072.4]
  input        io_rPort_1_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_1_output_0, // @[:@44072.4]
  input  [3:0] io_rPort_0_banks_1, // @[:@44072.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@44072.4]
  input  [7:0] io_rPort_0_ofs_0, // @[:@44072.4]
  input        io_rPort_0_en_0, // @[:@44072.4]
  input        io_rPort_0_backpressure, // @[:@44072.4]
  output [7:0] io_rPort_0_output_0, // @[:@44072.4]
  input  [3:0] io_wPort_7_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_7_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_7_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_7_data_0, // @[:@44072.4]
  input        io_wPort_7_en_0, // @[:@44072.4]
  input  [3:0] io_wPort_6_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_6_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_6_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_6_data_0, // @[:@44072.4]
  input        io_wPort_6_en_0, // @[:@44072.4]
  input  [3:0] io_wPort_5_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_5_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_5_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_5_data_0, // @[:@44072.4]
  input        io_wPort_5_en_0, // @[:@44072.4]
  input  [3:0] io_wPort_4_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_4_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_4_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_4_data_0, // @[:@44072.4]
  input        io_wPort_4_en_0, // @[:@44072.4]
  input  [3:0] io_wPort_3_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_3_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_3_data_0, // @[:@44072.4]
  input        io_wPort_3_en_0, // @[:@44072.4]
  input  [3:0] io_wPort_2_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_2_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_2_data_0, // @[:@44072.4]
  input        io_wPort_2_en_0, // @[:@44072.4]
  input  [3:0] io_wPort_1_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_1_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_1_data_0, // @[:@44072.4]
  input        io_wPort_1_en_0, // @[:@44072.4]
  input  [3:0] io_wPort_0_banks_1, // @[:@44072.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@44072.4]
  input  [7:0] io_wPort_0_ofs_0, // @[:@44072.4]
  input  [7:0] io_wPort_0_data_0, // @[:@44072.4]
  input        io_wPort_0_en_0 // @[:@44072.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@44319.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@44319.4]
  wire [7:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44319.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44319.4]
  wire [7:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44319.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@44319.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@44319.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@44319.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@44335.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@44335.4]
  wire [7:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44335.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44335.4]
  wire [7:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44335.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@44335.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@44335.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@44335.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@44351.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@44351.4]
  wire [7:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44351.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44351.4]
  wire [7:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44351.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@44351.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@44351.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@44351.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@44367.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@44367.4]
  wire [7:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44367.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44367.4]
  wire [7:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44367.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@44367.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@44367.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@44367.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@44383.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@44383.4]
  wire [7:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44383.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44383.4]
  wire [7:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44383.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@44383.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@44383.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@44383.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@44399.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@44399.4]
  wire [7:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44399.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44399.4]
  wire [7:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44399.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@44399.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@44399.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@44399.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@44415.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@44415.4]
  wire [7:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44415.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44415.4]
  wire [7:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44415.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@44415.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@44415.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@44415.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@44431.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@44431.4]
  wire [7:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44431.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44431.4]
  wire [7:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44431.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@44431.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@44431.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@44431.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@44447.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@44447.4]
  wire [7:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44447.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44447.4]
  wire [7:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44447.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@44447.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@44447.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@44447.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@44463.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@44463.4]
  wire [7:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44463.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44463.4]
  wire [7:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44463.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@44463.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@44463.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@44463.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@44479.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@44479.4]
  wire [7:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44479.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44479.4]
  wire [7:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44479.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@44479.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@44479.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@44479.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@44495.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@44495.4]
  wire [7:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44495.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44495.4]
  wire [7:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44495.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@44495.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@44495.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@44495.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@44511.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@44511.4]
  wire [7:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44511.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44511.4]
  wire [7:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44511.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@44511.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@44511.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@44511.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@44527.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@44527.4]
  wire [7:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44527.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44527.4]
  wire [7:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44527.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@44527.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@44527.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@44527.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@44543.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@44543.4]
  wire [7:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44543.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44543.4]
  wire [7:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44543.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@44543.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@44543.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@44543.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@44559.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@44559.4]
  wire [7:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44559.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44559.4]
  wire [7:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44559.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@44559.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@44559.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@44559.4]
  wire  Mem1D_16_clock; // @[MemPrimitives.scala 64:21:@44575.4]
  wire  Mem1D_16_reset; // @[MemPrimitives.scala 64:21:@44575.4]
  wire [7:0] Mem1D_16_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44575.4]
  wire  Mem1D_16_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44575.4]
  wire [7:0] Mem1D_16_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44575.4]
  wire [7:0] Mem1D_16_io_w_data_0; // @[MemPrimitives.scala 64:21:@44575.4]
  wire  Mem1D_16_io_w_en_0; // @[MemPrimitives.scala 64:21:@44575.4]
  wire [7:0] Mem1D_16_io_output; // @[MemPrimitives.scala 64:21:@44575.4]
  wire  Mem1D_17_clock; // @[MemPrimitives.scala 64:21:@44591.4]
  wire  Mem1D_17_reset; // @[MemPrimitives.scala 64:21:@44591.4]
  wire [7:0] Mem1D_17_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44591.4]
  wire  Mem1D_17_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44591.4]
  wire [7:0] Mem1D_17_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44591.4]
  wire [7:0] Mem1D_17_io_w_data_0; // @[MemPrimitives.scala 64:21:@44591.4]
  wire  Mem1D_17_io_w_en_0; // @[MemPrimitives.scala 64:21:@44591.4]
  wire [7:0] Mem1D_17_io_output; // @[MemPrimitives.scala 64:21:@44591.4]
  wire  Mem1D_18_clock; // @[MemPrimitives.scala 64:21:@44607.4]
  wire  Mem1D_18_reset; // @[MemPrimitives.scala 64:21:@44607.4]
  wire [7:0] Mem1D_18_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44607.4]
  wire  Mem1D_18_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44607.4]
  wire [7:0] Mem1D_18_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44607.4]
  wire [7:0] Mem1D_18_io_w_data_0; // @[MemPrimitives.scala 64:21:@44607.4]
  wire  Mem1D_18_io_w_en_0; // @[MemPrimitives.scala 64:21:@44607.4]
  wire [7:0] Mem1D_18_io_output; // @[MemPrimitives.scala 64:21:@44607.4]
  wire  Mem1D_19_clock; // @[MemPrimitives.scala 64:21:@44623.4]
  wire  Mem1D_19_reset; // @[MemPrimitives.scala 64:21:@44623.4]
  wire [7:0] Mem1D_19_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44623.4]
  wire  Mem1D_19_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44623.4]
  wire [7:0] Mem1D_19_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44623.4]
  wire [7:0] Mem1D_19_io_w_data_0; // @[MemPrimitives.scala 64:21:@44623.4]
  wire  Mem1D_19_io_w_en_0; // @[MemPrimitives.scala 64:21:@44623.4]
  wire [7:0] Mem1D_19_io_output; // @[MemPrimitives.scala 64:21:@44623.4]
  wire  Mem1D_20_clock; // @[MemPrimitives.scala 64:21:@44639.4]
  wire  Mem1D_20_reset; // @[MemPrimitives.scala 64:21:@44639.4]
  wire [7:0] Mem1D_20_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44639.4]
  wire  Mem1D_20_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44639.4]
  wire [7:0] Mem1D_20_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44639.4]
  wire [7:0] Mem1D_20_io_w_data_0; // @[MemPrimitives.scala 64:21:@44639.4]
  wire  Mem1D_20_io_w_en_0; // @[MemPrimitives.scala 64:21:@44639.4]
  wire [7:0] Mem1D_20_io_output; // @[MemPrimitives.scala 64:21:@44639.4]
  wire  Mem1D_21_clock; // @[MemPrimitives.scala 64:21:@44655.4]
  wire  Mem1D_21_reset; // @[MemPrimitives.scala 64:21:@44655.4]
  wire [7:0] Mem1D_21_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44655.4]
  wire  Mem1D_21_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44655.4]
  wire [7:0] Mem1D_21_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44655.4]
  wire [7:0] Mem1D_21_io_w_data_0; // @[MemPrimitives.scala 64:21:@44655.4]
  wire  Mem1D_21_io_w_en_0; // @[MemPrimitives.scala 64:21:@44655.4]
  wire [7:0] Mem1D_21_io_output; // @[MemPrimitives.scala 64:21:@44655.4]
  wire  Mem1D_22_clock; // @[MemPrimitives.scala 64:21:@44671.4]
  wire  Mem1D_22_reset; // @[MemPrimitives.scala 64:21:@44671.4]
  wire [7:0] Mem1D_22_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44671.4]
  wire  Mem1D_22_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44671.4]
  wire [7:0] Mem1D_22_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44671.4]
  wire [7:0] Mem1D_22_io_w_data_0; // @[MemPrimitives.scala 64:21:@44671.4]
  wire  Mem1D_22_io_w_en_0; // @[MemPrimitives.scala 64:21:@44671.4]
  wire [7:0] Mem1D_22_io_output; // @[MemPrimitives.scala 64:21:@44671.4]
  wire  Mem1D_23_clock; // @[MemPrimitives.scala 64:21:@44687.4]
  wire  Mem1D_23_reset; // @[MemPrimitives.scala 64:21:@44687.4]
  wire [7:0] Mem1D_23_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44687.4]
  wire  Mem1D_23_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44687.4]
  wire [7:0] Mem1D_23_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44687.4]
  wire [7:0] Mem1D_23_io_w_data_0; // @[MemPrimitives.scala 64:21:@44687.4]
  wire  Mem1D_23_io_w_en_0; // @[MemPrimitives.scala 64:21:@44687.4]
  wire [7:0] Mem1D_23_io_output; // @[MemPrimitives.scala 64:21:@44687.4]
  wire  Mem1D_24_clock; // @[MemPrimitives.scala 64:21:@44703.4]
  wire  Mem1D_24_reset; // @[MemPrimitives.scala 64:21:@44703.4]
  wire [7:0] Mem1D_24_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44703.4]
  wire  Mem1D_24_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44703.4]
  wire [7:0] Mem1D_24_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44703.4]
  wire [7:0] Mem1D_24_io_w_data_0; // @[MemPrimitives.scala 64:21:@44703.4]
  wire  Mem1D_24_io_w_en_0; // @[MemPrimitives.scala 64:21:@44703.4]
  wire [7:0] Mem1D_24_io_output; // @[MemPrimitives.scala 64:21:@44703.4]
  wire  Mem1D_25_clock; // @[MemPrimitives.scala 64:21:@44719.4]
  wire  Mem1D_25_reset; // @[MemPrimitives.scala 64:21:@44719.4]
  wire [7:0] Mem1D_25_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44719.4]
  wire  Mem1D_25_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44719.4]
  wire [7:0] Mem1D_25_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44719.4]
  wire [7:0] Mem1D_25_io_w_data_0; // @[MemPrimitives.scala 64:21:@44719.4]
  wire  Mem1D_25_io_w_en_0; // @[MemPrimitives.scala 64:21:@44719.4]
  wire [7:0] Mem1D_25_io_output; // @[MemPrimitives.scala 64:21:@44719.4]
  wire  Mem1D_26_clock; // @[MemPrimitives.scala 64:21:@44735.4]
  wire  Mem1D_26_reset; // @[MemPrimitives.scala 64:21:@44735.4]
  wire [7:0] Mem1D_26_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44735.4]
  wire  Mem1D_26_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44735.4]
  wire [7:0] Mem1D_26_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44735.4]
  wire [7:0] Mem1D_26_io_w_data_0; // @[MemPrimitives.scala 64:21:@44735.4]
  wire  Mem1D_26_io_w_en_0; // @[MemPrimitives.scala 64:21:@44735.4]
  wire [7:0] Mem1D_26_io_output; // @[MemPrimitives.scala 64:21:@44735.4]
  wire  Mem1D_27_clock; // @[MemPrimitives.scala 64:21:@44751.4]
  wire  Mem1D_27_reset; // @[MemPrimitives.scala 64:21:@44751.4]
  wire [7:0] Mem1D_27_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44751.4]
  wire  Mem1D_27_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44751.4]
  wire [7:0] Mem1D_27_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44751.4]
  wire [7:0] Mem1D_27_io_w_data_0; // @[MemPrimitives.scala 64:21:@44751.4]
  wire  Mem1D_27_io_w_en_0; // @[MemPrimitives.scala 64:21:@44751.4]
  wire [7:0] Mem1D_27_io_output; // @[MemPrimitives.scala 64:21:@44751.4]
  wire  Mem1D_28_clock; // @[MemPrimitives.scala 64:21:@44767.4]
  wire  Mem1D_28_reset; // @[MemPrimitives.scala 64:21:@44767.4]
  wire [7:0] Mem1D_28_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44767.4]
  wire  Mem1D_28_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44767.4]
  wire [7:0] Mem1D_28_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44767.4]
  wire [7:0] Mem1D_28_io_w_data_0; // @[MemPrimitives.scala 64:21:@44767.4]
  wire  Mem1D_28_io_w_en_0; // @[MemPrimitives.scala 64:21:@44767.4]
  wire [7:0] Mem1D_28_io_output; // @[MemPrimitives.scala 64:21:@44767.4]
  wire  Mem1D_29_clock; // @[MemPrimitives.scala 64:21:@44783.4]
  wire  Mem1D_29_reset; // @[MemPrimitives.scala 64:21:@44783.4]
  wire [7:0] Mem1D_29_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44783.4]
  wire  Mem1D_29_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44783.4]
  wire [7:0] Mem1D_29_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44783.4]
  wire [7:0] Mem1D_29_io_w_data_0; // @[MemPrimitives.scala 64:21:@44783.4]
  wire  Mem1D_29_io_w_en_0; // @[MemPrimitives.scala 64:21:@44783.4]
  wire [7:0] Mem1D_29_io_output; // @[MemPrimitives.scala 64:21:@44783.4]
  wire  Mem1D_30_clock; // @[MemPrimitives.scala 64:21:@44799.4]
  wire  Mem1D_30_reset; // @[MemPrimitives.scala 64:21:@44799.4]
  wire [7:0] Mem1D_30_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44799.4]
  wire  Mem1D_30_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44799.4]
  wire [7:0] Mem1D_30_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44799.4]
  wire [7:0] Mem1D_30_io_w_data_0; // @[MemPrimitives.scala 64:21:@44799.4]
  wire  Mem1D_30_io_w_en_0; // @[MemPrimitives.scala 64:21:@44799.4]
  wire [7:0] Mem1D_30_io_output; // @[MemPrimitives.scala 64:21:@44799.4]
  wire  Mem1D_31_clock; // @[MemPrimitives.scala 64:21:@44815.4]
  wire  Mem1D_31_reset; // @[MemPrimitives.scala 64:21:@44815.4]
  wire [7:0] Mem1D_31_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44815.4]
  wire  Mem1D_31_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44815.4]
  wire [7:0] Mem1D_31_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44815.4]
  wire [7:0] Mem1D_31_io_w_data_0; // @[MemPrimitives.scala 64:21:@44815.4]
  wire  Mem1D_31_io_w_en_0; // @[MemPrimitives.scala 64:21:@44815.4]
  wire [7:0] Mem1D_31_io_output; // @[MemPrimitives.scala 64:21:@44815.4]
  wire  Mem1D_32_clock; // @[MemPrimitives.scala 64:21:@44831.4]
  wire  Mem1D_32_reset; // @[MemPrimitives.scala 64:21:@44831.4]
  wire [7:0] Mem1D_32_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44831.4]
  wire  Mem1D_32_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44831.4]
  wire [7:0] Mem1D_32_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44831.4]
  wire [7:0] Mem1D_32_io_w_data_0; // @[MemPrimitives.scala 64:21:@44831.4]
  wire  Mem1D_32_io_w_en_0; // @[MemPrimitives.scala 64:21:@44831.4]
  wire [7:0] Mem1D_32_io_output; // @[MemPrimitives.scala 64:21:@44831.4]
  wire  Mem1D_33_clock; // @[MemPrimitives.scala 64:21:@44847.4]
  wire  Mem1D_33_reset; // @[MemPrimitives.scala 64:21:@44847.4]
  wire [7:0] Mem1D_33_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44847.4]
  wire  Mem1D_33_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44847.4]
  wire [7:0] Mem1D_33_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44847.4]
  wire [7:0] Mem1D_33_io_w_data_0; // @[MemPrimitives.scala 64:21:@44847.4]
  wire  Mem1D_33_io_w_en_0; // @[MemPrimitives.scala 64:21:@44847.4]
  wire [7:0] Mem1D_33_io_output; // @[MemPrimitives.scala 64:21:@44847.4]
  wire  Mem1D_34_clock; // @[MemPrimitives.scala 64:21:@44863.4]
  wire  Mem1D_34_reset; // @[MemPrimitives.scala 64:21:@44863.4]
  wire [7:0] Mem1D_34_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44863.4]
  wire  Mem1D_34_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44863.4]
  wire [7:0] Mem1D_34_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44863.4]
  wire [7:0] Mem1D_34_io_w_data_0; // @[MemPrimitives.scala 64:21:@44863.4]
  wire  Mem1D_34_io_w_en_0; // @[MemPrimitives.scala 64:21:@44863.4]
  wire [7:0] Mem1D_34_io_output; // @[MemPrimitives.scala 64:21:@44863.4]
  wire  Mem1D_35_clock; // @[MemPrimitives.scala 64:21:@44879.4]
  wire  Mem1D_35_reset; // @[MemPrimitives.scala 64:21:@44879.4]
  wire [7:0] Mem1D_35_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44879.4]
  wire  Mem1D_35_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44879.4]
  wire [7:0] Mem1D_35_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44879.4]
  wire [7:0] Mem1D_35_io_w_data_0; // @[MemPrimitives.scala 64:21:@44879.4]
  wire  Mem1D_35_io_w_en_0; // @[MemPrimitives.scala 64:21:@44879.4]
  wire [7:0] Mem1D_35_io_output; // @[MemPrimitives.scala 64:21:@44879.4]
  wire  Mem1D_36_clock; // @[MemPrimitives.scala 64:21:@44895.4]
  wire  Mem1D_36_reset; // @[MemPrimitives.scala 64:21:@44895.4]
  wire [7:0] Mem1D_36_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44895.4]
  wire  Mem1D_36_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44895.4]
  wire [7:0] Mem1D_36_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44895.4]
  wire [7:0] Mem1D_36_io_w_data_0; // @[MemPrimitives.scala 64:21:@44895.4]
  wire  Mem1D_36_io_w_en_0; // @[MemPrimitives.scala 64:21:@44895.4]
  wire [7:0] Mem1D_36_io_output; // @[MemPrimitives.scala 64:21:@44895.4]
  wire  Mem1D_37_clock; // @[MemPrimitives.scala 64:21:@44911.4]
  wire  Mem1D_37_reset; // @[MemPrimitives.scala 64:21:@44911.4]
  wire [7:0] Mem1D_37_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44911.4]
  wire  Mem1D_37_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44911.4]
  wire [7:0] Mem1D_37_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44911.4]
  wire [7:0] Mem1D_37_io_w_data_0; // @[MemPrimitives.scala 64:21:@44911.4]
  wire  Mem1D_37_io_w_en_0; // @[MemPrimitives.scala 64:21:@44911.4]
  wire [7:0] Mem1D_37_io_output; // @[MemPrimitives.scala 64:21:@44911.4]
  wire  Mem1D_38_clock; // @[MemPrimitives.scala 64:21:@44927.4]
  wire  Mem1D_38_reset; // @[MemPrimitives.scala 64:21:@44927.4]
  wire [7:0] Mem1D_38_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44927.4]
  wire  Mem1D_38_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44927.4]
  wire [7:0] Mem1D_38_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44927.4]
  wire [7:0] Mem1D_38_io_w_data_0; // @[MemPrimitives.scala 64:21:@44927.4]
  wire  Mem1D_38_io_w_en_0; // @[MemPrimitives.scala 64:21:@44927.4]
  wire [7:0] Mem1D_38_io_output; // @[MemPrimitives.scala 64:21:@44927.4]
  wire  Mem1D_39_clock; // @[MemPrimitives.scala 64:21:@44943.4]
  wire  Mem1D_39_reset; // @[MemPrimitives.scala 64:21:@44943.4]
  wire [7:0] Mem1D_39_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@44943.4]
  wire  Mem1D_39_io_r_backpressure; // @[MemPrimitives.scala 64:21:@44943.4]
  wire [7:0] Mem1D_39_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@44943.4]
  wire [7:0] Mem1D_39_io_w_data_0; // @[MemPrimitives.scala 64:21:@44943.4]
  wire  Mem1D_39_io_w_en_0; // @[MemPrimitives.scala 64:21:@44943.4]
  wire [7:0] Mem1D_39_io_output; // @[MemPrimitives.scala 64:21:@44943.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_9; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_10; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_11; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_12; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_13; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_ins_14; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_9; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_10; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_11; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_12; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_13; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_io_outs_14; // @[MemPrimitives.scala 121:29:@46339.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_9; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_10; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_11; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_12; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_13; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_ins_14; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_9; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_10; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_11; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_12; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_13; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_1_io_outs_14; // @[MemPrimitives.scala 121:29:@46482.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_9; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_10; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_11; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_12; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_13; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_ins_14; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_9; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_10; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_11; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_12; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_13; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_2_io_outs_14; // @[MemPrimitives.scala 121:29:@46625.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_9; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_10; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_11; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_12; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_13; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_ins_14; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_9; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_10; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_11; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_12; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_13; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_3_io_outs_14; // @[MemPrimitives.scala 121:29:@46768.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_9; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_10; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_11; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_12; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_13; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_ins_14; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_9; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_10; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_11; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_12; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_13; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_4_io_outs_14; // @[MemPrimitives.scala 121:29:@46911.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_9; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_10; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_11; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_12; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_13; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_ins_14; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_9; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_10; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_11; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_12; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_13; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_5_io_outs_14; // @[MemPrimitives.scala 121:29:@47054.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_9; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_10; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_11; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_12; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_13; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_ins_14; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_9; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_10; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_11; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_12; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_13; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_6_io_outs_14; // @[MemPrimitives.scala 121:29:@47197.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_9; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_10; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_11; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_12; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_13; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_ins_14; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_9; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_10; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_11; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_12; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_13; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_7_io_outs_14; // @[MemPrimitives.scala 121:29:@47340.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_9; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_10; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_11; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_12; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_13; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_ins_14; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_9; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_10; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_11; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_12; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_13; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_8_io_outs_14; // @[MemPrimitives.scala 121:29:@47483.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_9; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_10; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_11; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_12; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_13; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_ins_14; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_9; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_10; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_11; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_12; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_13; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_9_io_outs_14; // @[MemPrimitives.scala 121:29:@47626.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_9; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_10; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_11; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_12; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_13; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_ins_14; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_9; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_10; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_11; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_12; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_13; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_10_io_outs_14; // @[MemPrimitives.scala 121:29:@47769.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_9; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_10; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_11; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_12; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_13; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_ins_14; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_9; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_10; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_11; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_12; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_13; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_11_io_outs_14; // @[MemPrimitives.scala 121:29:@47912.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_6; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_7; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_8; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_9; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_10; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_11; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_12; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_13; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_ins_14; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_6; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_7; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_8; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_9; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_10; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_11; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_12; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_13; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_12_io_outs_14; // @[MemPrimitives.scala 121:29:@48055.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_6; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_7; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_8; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_9; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_10; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_11; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_12; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_13; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_ins_14; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_6; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_7; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_8; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_9; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_10; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_11; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_12; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_13; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_13_io_outs_14; // @[MemPrimitives.scala 121:29:@48198.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_8; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_9; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_10; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_11; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_12; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_13; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_ins_14; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_8; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_9; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_10; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_11; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_12; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_13; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_14_io_outs_14; // @[MemPrimitives.scala 121:29:@48341.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_8; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_9; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_10; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_11; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_12; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_13; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_ins_14; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_8; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_9; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_10; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_11; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_12; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_13; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_15_io_outs_14; // @[MemPrimitives.scala 121:29:@48484.4]
  wire  StickySelects_16_clock; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_reset; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_0; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_1; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_2; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_3; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_4; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_5; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_6; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_7; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_8; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_9; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_10; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_11; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_12; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_13; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_ins_14; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_0; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_1; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_2; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_3; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_4; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_5; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_6; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_7; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_8; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_9; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_10; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_11; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_12; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_13; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_16_io_outs_14; // @[MemPrimitives.scala 121:29:@48627.4]
  wire  StickySelects_17_clock; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_reset; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_0; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_1; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_2; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_3; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_4; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_5; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_6; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_7; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_8; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_9; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_10; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_11; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_12; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_13; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_ins_14; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_0; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_1; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_2; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_3; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_4; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_5; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_6; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_7; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_8; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_9; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_10; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_11; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_12; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_13; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_17_io_outs_14; // @[MemPrimitives.scala 121:29:@48770.4]
  wire  StickySelects_18_clock; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_reset; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_0; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_1; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_2; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_3; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_4; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_5; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_6; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_7; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_8; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_9; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_10; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_11; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_12; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_13; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_ins_14; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_0; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_1; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_2; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_3; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_4; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_5; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_6; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_7; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_8; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_9; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_10; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_11; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_12; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_13; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_18_io_outs_14; // @[MemPrimitives.scala 121:29:@48913.4]
  wire  StickySelects_19_clock; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_reset; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_0; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_1; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_2; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_3; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_4; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_5; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_6; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_7; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_8; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_9; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_10; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_11; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_12; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_13; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_ins_14; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_0; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_1; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_2; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_3; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_4; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_5; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_6; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_7; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_8; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_9; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_10; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_11; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_12; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_13; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_19_io_outs_14; // @[MemPrimitives.scala 121:29:@49056.4]
  wire  StickySelects_20_clock; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_reset; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_0; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_1; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_2; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_3; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_4; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_5; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_6; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_7; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_8; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_9; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_10; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_11; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_12; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_13; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_ins_14; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_0; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_1; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_2; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_3; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_4; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_5; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_6; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_7; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_8; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_9; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_10; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_11; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_12; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_13; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_20_io_outs_14; // @[MemPrimitives.scala 121:29:@49199.4]
  wire  StickySelects_21_clock; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_reset; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_0; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_1; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_2; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_3; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_4; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_5; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_6; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_7; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_8; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_9; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_10; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_11; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_12; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_13; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_ins_14; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_0; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_1; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_2; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_3; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_4; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_5; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_6; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_7; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_8; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_9; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_10; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_11; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_12; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_13; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_21_io_outs_14; // @[MemPrimitives.scala 121:29:@49342.4]
  wire  StickySelects_22_clock; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_reset; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_0; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_1; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_2; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_3; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_4; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_5; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_6; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_7; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_8; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_9; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_10; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_11; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_12; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_13; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_ins_14; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_0; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_1; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_2; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_3; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_4; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_5; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_6; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_7; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_8; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_9; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_10; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_11; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_12; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_13; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_22_io_outs_14; // @[MemPrimitives.scala 121:29:@49485.4]
  wire  StickySelects_23_clock; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_reset; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_0; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_1; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_2; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_3; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_4; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_5; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_6; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_7; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_8; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_9; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_10; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_11; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_12; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_13; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_ins_14; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_0; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_1; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_2; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_3; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_4; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_5; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_6; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_7; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_8; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_9; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_10; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_11; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_12; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_13; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_23_io_outs_14; // @[MemPrimitives.scala 121:29:@49628.4]
  wire  StickySelects_24_clock; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_reset; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_0; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_1; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_2; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_3; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_4; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_5; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_6; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_7; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_8; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_9; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_10; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_11; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_12; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_13; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_ins_14; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_0; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_1; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_2; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_3; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_4; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_5; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_6; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_7; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_8; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_9; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_10; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_11; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_12; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_13; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_24_io_outs_14; // @[MemPrimitives.scala 121:29:@49771.4]
  wire  StickySelects_25_clock; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_reset; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_0; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_1; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_2; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_3; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_4; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_5; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_6; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_7; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_8; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_9; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_10; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_11; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_12; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_13; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_ins_14; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_0; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_1; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_2; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_3; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_4; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_5; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_6; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_7; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_8; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_9; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_10; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_11; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_12; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_13; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_25_io_outs_14; // @[MemPrimitives.scala 121:29:@49914.4]
  wire  StickySelects_26_clock; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_reset; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_0; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_1; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_2; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_3; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_4; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_5; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_6; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_7; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_8; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_9; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_10; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_11; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_12; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_13; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_ins_14; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_0; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_1; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_2; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_3; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_4; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_5; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_6; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_7; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_8; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_9; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_10; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_11; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_12; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_13; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_26_io_outs_14; // @[MemPrimitives.scala 121:29:@50057.4]
  wire  StickySelects_27_clock; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_reset; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_0; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_1; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_2; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_3; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_4; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_5; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_6; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_7; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_8; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_9; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_10; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_11; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_12; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_13; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_ins_14; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_0; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_1; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_2; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_3; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_4; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_5; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_6; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_7; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_8; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_9; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_10; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_11; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_12; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_13; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_27_io_outs_14; // @[MemPrimitives.scala 121:29:@50200.4]
  wire  StickySelects_28_clock; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_reset; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_0; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_1; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_2; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_3; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_4; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_5; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_6; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_7; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_8; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_9; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_10; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_11; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_12; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_13; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_ins_14; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_0; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_1; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_2; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_3; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_4; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_5; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_6; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_7; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_8; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_9; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_10; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_11; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_12; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_13; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_28_io_outs_14; // @[MemPrimitives.scala 121:29:@50343.4]
  wire  StickySelects_29_clock; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_reset; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_0; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_1; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_2; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_3; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_4; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_5; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_6; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_7; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_8; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_9; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_10; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_11; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_12; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_13; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_ins_14; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_0; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_1; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_2; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_3; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_4; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_5; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_6; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_7; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_8; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_9; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_10; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_11; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_12; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_13; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_29_io_outs_14; // @[MemPrimitives.scala 121:29:@50486.4]
  wire  StickySelects_30_clock; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_reset; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_0; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_1; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_2; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_3; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_4; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_5; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_6; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_7; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_8; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_9; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_10; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_11; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_12; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_13; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_ins_14; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_0; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_1; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_2; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_3; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_4; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_5; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_6; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_7; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_8; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_9; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_10; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_11; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_12; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_13; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_30_io_outs_14; // @[MemPrimitives.scala 121:29:@50629.4]
  wire  StickySelects_31_clock; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_reset; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_0; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_1; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_2; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_3; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_4; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_5; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_6; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_7; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_8; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_9; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_10; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_11; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_12; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_13; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_ins_14; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_0; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_1; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_2; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_3; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_4; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_5; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_6; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_7; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_8; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_9; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_10; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_11; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_12; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_13; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_31_io_outs_14; // @[MemPrimitives.scala 121:29:@50772.4]
  wire  StickySelects_32_clock; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_reset; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_0; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_1; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_2; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_3; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_4; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_5; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_6; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_7; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_8; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_9; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_10; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_11; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_12; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_13; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_ins_14; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_0; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_1; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_2; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_3; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_4; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_5; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_6; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_7; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_8; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_9; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_10; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_11; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_12; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_13; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_32_io_outs_14; // @[MemPrimitives.scala 121:29:@50915.4]
  wire  StickySelects_33_clock; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_reset; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_0; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_1; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_2; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_3; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_4; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_5; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_6; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_7; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_8; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_9; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_10; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_11; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_12; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_13; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_ins_14; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_0; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_1; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_2; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_3; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_4; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_5; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_6; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_7; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_8; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_9; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_10; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_11; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_12; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_13; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_33_io_outs_14; // @[MemPrimitives.scala 121:29:@51058.4]
  wire  StickySelects_34_clock; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_reset; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_0; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_1; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_2; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_3; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_4; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_5; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_6; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_7; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_8; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_9; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_10; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_11; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_12; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_13; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_ins_14; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_0; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_1; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_2; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_3; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_4; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_5; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_6; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_7; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_8; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_9; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_10; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_11; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_12; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_13; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_34_io_outs_14; // @[MemPrimitives.scala 121:29:@51201.4]
  wire  StickySelects_35_clock; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_reset; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_0; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_1; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_2; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_3; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_4; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_5; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_6; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_7; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_8; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_9; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_10; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_11; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_12; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_13; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_ins_14; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_0; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_1; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_2; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_3; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_4; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_5; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_6; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_7; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_8; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_9; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_10; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_11; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_12; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_13; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_35_io_outs_14; // @[MemPrimitives.scala 121:29:@51344.4]
  wire  StickySelects_36_clock; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_reset; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_0; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_1; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_2; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_3; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_4; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_5; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_6; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_7; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_8; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_9; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_10; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_11; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_12; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_13; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_ins_14; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_0; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_1; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_2; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_3; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_4; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_5; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_6; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_7; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_8; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_9; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_10; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_11; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_12; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_13; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_36_io_outs_14; // @[MemPrimitives.scala 121:29:@51487.4]
  wire  StickySelects_37_clock; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_reset; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_0; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_1; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_2; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_3; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_4; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_5; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_6; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_7; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_8; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_9; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_10; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_11; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_12; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_13; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_ins_14; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_0; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_1; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_2; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_3; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_4; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_5; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_6; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_7; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_8; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_9; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_10; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_11; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_12; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_13; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_37_io_outs_14; // @[MemPrimitives.scala 121:29:@51630.4]
  wire  StickySelects_38_clock; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_reset; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_0; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_1; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_2; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_3; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_4; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_5; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_6; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_7; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_8; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_9; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_10; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_11; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_12; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_13; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_ins_14; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_0; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_1; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_2; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_3; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_4; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_5; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_6; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_7; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_8; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_9; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_10; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_11; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_12; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_13; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_38_io_outs_14; // @[MemPrimitives.scala 121:29:@51773.4]
  wire  StickySelects_39_clock; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_reset; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_0; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_1; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_2; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_3; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_4; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_5; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_6; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_7; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_8; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_9; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_10; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_11; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_12; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_13; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_ins_14; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_0; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_1; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_2; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_3; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_4; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_5; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_6; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_7; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_8; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_9; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_10; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_11; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_12; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_13; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  StickySelects_39_io_outs_14; // @[MemPrimitives.scala 121:29:@51916.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@52060.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@52060.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@52060.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@52060.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@52060.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@52068.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@52068.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@52068.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@52068.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@52068.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@52076.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@52076.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@52076.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@52076.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@52076.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@52084.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@52084.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@52084.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@52084.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@52084.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@52092.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@52092.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@52092.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@52092.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@52092.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@52100.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@52100.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@52100.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@52100.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@52100.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@52108.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@52108.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@52108.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@52108.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@52108.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@52116.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@52116.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@52116.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@52116.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@52116.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@52124.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@52124.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@52124.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@52124.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@52124.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@52132.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@52132.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@52132.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@52132.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@52132.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@52140.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@52140.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@52140.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@52140.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@52140.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@52148.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@52148.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@52148.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@52148.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@52148.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@52156.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@52156.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@52156.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@52156.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@52156.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@52164.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@52164.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@52164.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@52164.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@52164.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@52172.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@52172.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@52172.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@52172.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@52172.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@52180.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@52180.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@52180.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@52180.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@52180.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@52188.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@52188.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@52188.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@52188.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@52188.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@52196.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@52196.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@52196.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@52196.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@52196.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@52204.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@52204.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@52204.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@52204.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@52204.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@52212.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@52212.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@52212.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@52212.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@52212.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@52300.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@52300.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@52300.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@52300.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@52300.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@52308.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@52308.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@52308.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@52308.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@52308.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@52316.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@52316.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@52316.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@52316.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@52316.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@52324.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@52324.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@52324.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@52324.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@52324.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@52332.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@52332.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@52332.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@52332.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@52332.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@52340.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@52340.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@52340.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@52340.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@52340.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@52348.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@52348.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@52348.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@52348.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@52348.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@52356.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@52356.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@52356.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@52356.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@52356.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@52364.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@52364.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@52364.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@52364.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@52364.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@52372.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@52372.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@52372.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@52372.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@52372.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@52380.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@52380.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@52380.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@52380.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@52380.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@52388.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@52388.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@52388.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@52388.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@52388.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@52396.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@52396.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@52396.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@52396.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@52396.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@52412.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@52412.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@52412.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@52412.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@52412.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@52420.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@52420.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@52420.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@52420.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@52420.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@52428.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@52428.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@52428.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@52428.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@52428.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@52436.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@52436.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@52436.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@52436.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@52436.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@52444.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@52444.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@52444.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@52444.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@52444.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@52452.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@52452.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@52452.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@52452.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@52452.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@52540.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@52540.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@52540.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@52540.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@52540.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@52548.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@52548.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@52548.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@52548.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@52548.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@52556.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@52556.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@52556.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@52556.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@52556.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@52564.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@52564.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@52564.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@52564.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@52564.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@52572.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@52572.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@52572.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@52572.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@52572.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@52580.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@52580.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@52580.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@52580.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@52580.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@52588.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@52588.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@52588.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@52588.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@52588.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@52596.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@52596.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@52596.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@52596.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@52596.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@52604.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@52604.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@52604.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@52604.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@52604.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@52612.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@52612.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@52612.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@52612.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@52612.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@52620.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@52620.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@52620.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@52620.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@52620.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@52628.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@52628.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@52628.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@52628.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@52628.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@52636.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@52636.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@52636.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@52636.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@52636.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@52644.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@52644.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@52644.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@52644.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@52644.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@52652.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@52652.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@52652.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@52652.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@52652.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@52660.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@52660.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@52660.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@52660.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@52660.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@52668.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@52668.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@52668.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@52668.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@52668.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@52676.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@52676.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@52676.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@52676.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@52676.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@52684.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@52684.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@52684.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@52684.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@52684.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@52692.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@52692.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@52692.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@52692.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@52692.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@52780.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@52780.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@52780.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@52780.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@52780.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@52788.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@52788.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@52788.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@52788.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@52788.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@52796.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@52796.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@52796.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@52796.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@52796.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@52804.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@52804.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@52804.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@52804.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@52804.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@52812.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@52812.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@52812.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@52812.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@52812.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@52820.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@52820.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@52820.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@52820.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@52820.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@52828.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@52828.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@52828.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@52828.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@52828.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@52836.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@52836.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@52836.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@52836.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@52836.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@52844.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@52844.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@52844.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@52844.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@52844.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@52852.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@52852.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@52852.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@52852.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@52852.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@52860.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@52860.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@52860.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@52860.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@52860.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@52868.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@52868.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@52868.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@52868.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@52868.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@52876.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@52876.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@52876.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@52876.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@52876.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@52884.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@52884.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@52884.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@52884.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@52884.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@52892.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@52892.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@52892.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@52892.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@52892.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@52900.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@52900.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@52900.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@52900.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@52900.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@52908.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@52908.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@52908.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@52908.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@52908.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@52916.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@52916.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@52916.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@52916.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@52916.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@52924.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@52924.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@52924.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@52924.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@52924.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@52932.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@52932.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@52932.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@52932.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@52932.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@53020.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@53020.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@53020.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@53020.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@53020.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@53028.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@53028.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@53028.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@53028.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@53028.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@53036.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@53036.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@53036.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@53036.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@53036.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@53044.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@53044.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@53044.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@53044.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@53044.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@53052.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@53052.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@53052.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@53052.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@53052.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@53060.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@53060.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@53060.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@53060.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@53060.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@53068.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@53068.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@53068.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@53068.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@53068.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@53076.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@53076.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@53076.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@53076.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@53076.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@53084.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@53084.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@53084.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@53084.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@53084.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@53092.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@53092.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@53092.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@53092.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@53092.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@53100.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@53100.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@53100.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@53100.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@53100.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@53108.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@53108.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@53108.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@53108.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@53108.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@53116.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@53116.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@53116.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@53116.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@53116.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@53124.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@53124.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@53124.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@53124.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@53124.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@53132.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@53132.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@53132.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@53132.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@53132.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@53140.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@53140.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@53140.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@53140.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@53140.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@53148.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@53148.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@53148.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@53148.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@53148.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@53156.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@53156.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@53156.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@53156.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@53156.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@53164.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@53164.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@53164.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@53164.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@53164.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@53172.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@53172.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@53172.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@53172.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@53172.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@53260.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@53260.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@53260.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@53260.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@53260.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@53268.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@53268.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@53268.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@53268.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@53268.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@53276.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@53276.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@53276.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@53276.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@53276.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@53284.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@53284.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@53284.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@53284.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@53284.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@53292.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@53292.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@53292.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@53292.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@53292.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@53300.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@53300.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@53300.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@53300.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@53300.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@53308.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@53308.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@53308.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@53308.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@53308.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@53316.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@53316.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@53316.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@53316.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@53316.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@53324.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@53324.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@53324.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@53324.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@53324.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@53332.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@53332.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@53332.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@53332.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@53332.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@53340.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@53340.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@53340.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@53340.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@53340.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@53348.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@53348.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@53348.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@53348.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@53348.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@53356.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@53356.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@53356.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@53356.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@53356.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@53364.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@53364.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@53364.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@53364.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@53364.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@53372.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@53372.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@53372.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@53372.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@53372.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@53380.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@53380.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@53380.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@53380.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@53380.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@53388.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@53388.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@53388.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@53388.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@53388.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@53396.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@53396.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@53396.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@53396.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@53396.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@53404.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@53404.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@53404.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@53404.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@53404.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@53412.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@53412.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@53412.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@53412.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@53412.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@53500.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@53500.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@53500.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@53500.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@53500.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@53508.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@53508.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@53508.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@53508.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@53508.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@53516.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@53516.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@53516.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@53516.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@53516.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@53524.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@53524.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@53524.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@53524.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@53524.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@53532.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@53532.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@53532.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@53532.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@53532.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@53540.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@53540.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@53540.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@53540.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@53540.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@53548.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@53548.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@53548.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@53548.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@53548.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@53564.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@53564.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@53564.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@53564.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@53564.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@53572.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@53572.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@53572.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@53572.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@53572.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@53580.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@53580.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@53580.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@53580.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@53580.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@53588.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@53588.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@53588.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@53588.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@53588.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@53596.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@53596.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@53596.4]
  wire  RetimeWrapper_132_io_in; // @[package.scala 93:22:@53596.4]
  wire  RetimeWrapper_132_io_out; // @[package.scala 93:22:@53596.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@53604.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@53604.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@53604.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@53604.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@53604.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@53612.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@53612.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@53612.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@53612.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@53612.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@53620.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@53620.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@53620.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@53620.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@53620.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@53628.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@53628.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@53628.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@53628.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@53628.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@53636.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@53636.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@53636.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@53636.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@53636.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@53644.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@53644.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@53644.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@53644.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@53644.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@53652.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@53652.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@53652.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@53652.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@53652.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@53740.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@53740.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@53740.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@53740.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@53740.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@53748.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@53748.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@53748.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@53748.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@53748.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@53756.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@53756.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@53756.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@53756.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@53756.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@53764.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@53764.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@53764.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@53764.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@53764.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@53772.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@53772.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@53772.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@53772.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@53772.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@53780.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@53780.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@53780.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@53780.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@53780.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@53788.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@53788.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@53788.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@53788.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@53788.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@53796.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@53796.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@53796.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@53796.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@53796.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@53804.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@53804.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@53804.4]
  wire  RetimeWrapper_148_io_in; // @[package.scala 93:22:@53804.4]
  wire  RetimeWrapper_148_io_out; // @[package.scala 93:22:@53804.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@53812.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@53812.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@53812.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@53812.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@53812.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@53820.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@53820.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@53820.4]
  wire  RetimeWrapper_150_io_in; // @[package.scala 93:22:@53820.4]
  wire  RetimeWrapper_150_io_out; // @[package.scala 93:22:@53820.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@53828.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@53828.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@53828.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@53828.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@53828.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@53836.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@53836.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@53836.4]
  wire  RetimeWrapper_152_io_in; // @[package.scala 93:22:@53836.4]
  wire  RetimeWrapper_152_io_out; // @[package.scala 93:22:@53836.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@53844.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@53844.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@53844.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@53844.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@53844.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@53852.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@53852.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@53852.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@53852.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@53852.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@53860.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@53860.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@53860.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@53860.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@53860.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@53868.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@53868.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@53868.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@53868.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@53868.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@53876.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@53876.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@53876.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@53876.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@53876.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@53884.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@53884.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@53884.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@53884.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@53884.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@53892.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@53892.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@53892.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@53892.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@53892.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@53980.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@53980.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@53980.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@53980.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@53980.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@53988.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@53988.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@53988.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@53988.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@53988.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@53996.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@53996.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@53996.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@53996.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@53996.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@54004.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@54004.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@54004.4]
  wire  RetimeWrapper_163_io_in; // @[package.scala 93:22:@54004.4]
  wire  RetimeWrapper_163_io_out; // @[package.scala 93:22:@54004.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@54012.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@54012.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@54012.4]
  wire  RetimeWrapper_164_io_in; // @[package.scala 93:22:@54012.4]
  wire  RetimeWrapper_164_io_out; // @[package.scala 93:22:@54012.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@54020.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@54020.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@54020.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@54020.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@54020.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@54028.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@54028.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@54028.4]
  wire  RetimeWrapper_166_io_in; // @[package.scala 93:22:@54028.4]
  wire  RetimeWrapper_166_io_out; // @[package.scala 93:22:@54028.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@54036.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@54036.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@54036.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@54036.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@54036.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@54044.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@54044.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@54044.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@54044.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@54044.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@54052.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@54052.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@54052.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@54052.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@54052.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@54060.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@54060.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@54060.4]
  wire  RetimeWrapper_170_io_in; // @[package.scala 93:22:@54060.4]
  wire  RetimeWrapper_170_io_out; // @[package.scala 93:22:@54060.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@54068.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@54068.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@54068.4]
  wire  RetimeWrapper_171_io_in; // @[package.scala 93:22:@54068.4]
  wire  RetimeWrapper_171_io_out; // @[package.scala 93:22:@54068.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@54076.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@54076.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@54076.4]
  wire  RetimeWrapper_172_io_in; // @[package.scala 93:22:@54076.4]
  wire  RetimeWrapper_172_io_out; // @[package.scala 93:22:@54076.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@54084.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@54084.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@54084.4]
  wire  RetimeWrapper_173_io_in; // @[package.scala 93:22:@54084.4]
  wire  RetimeWrapper_173_io_out; // @[package.scala 93:22:@54084.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@54092.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@54092.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@54092.4]
  wire  RetimeWrapper_174_io_in; // @[package.scala 93:22:@54092.4]
  wire  RetimeWrapper_174_io_out; // @[package.scala 93:22:@54092.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@54100.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@54100.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@54100.4]
  wire  RetimeWrapper_175_io_in; // @[package.scala 93:22:@54100.4]
  wire  RetimeWrapper_175_io_out; // @[package.scala 93:22:@54100.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@54108.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@54108.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@54108.4]
  wire  RetimeWrapper_176_io_in; // @[package.scala 93:22:@54108.4]
  wire  RetimeWrapper_176_io_out; // @[package.scala 93:22:@54108.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_177_io_in; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_177_io_out; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@54124.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@54124.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@54124.4]
  wire  RetimeWrapper_178_io_in; // @[package.scala 93:22:@54124.4]
  wire  RetimeWrapper_178_io_out; // @[package.scala 93:22:@54124.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@54132.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@54132.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@54132.4]
  wire  RetimeWrapper_179_io_in; // @[package.scala 93:22:@54132.4]
  wire  RetimeWrapper_179_io_out; // @[package.scala 93:22:@54132.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@54220.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@54220.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@54220.4]
  wire  RetimeWrapper_180_io_in; // @[package.scala 93:22:@54220.4]
  wire  RetimeWrapper_180_io_out; // @[package.scala 93:22:@54220.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@54228.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@54228.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@54228.4]
  wire  RetimeWrapper_181_io_in; // @[package.scala 93:22:@54228.4]
  wire  RetimeWrapper_181_io_out; // @[package.scala 93:22:@54228.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@54236.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@54236.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@54236.4]
  wire  RetimeWrapper_182_io_in; // @[package.scala 93:22:@54236.4]
  wire  RetimeWrapper_182_io_out; // @[package.scala 93:22:@54236.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@54244.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@54244.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@54244.4]
  wire  RetimeWrapper_183_io_in; // @[package.scala 93:22:@54244.4]
  wire  RetimeWrapper_183_io_out; // @[package.scala 93:22:@54244.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@54252.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@54252.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@54252.4]
  wire  RetimeWrapper_184_io_in; // @[package.scala 93:22:@54252.4]
  wire  RetimeWrapper_184_io_out; // @[package.scala 93:22:@54252.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@54260.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@54260.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@54260.4]
  wire  RetimeWrapper_185_io_in; // @[package.scala 93:22:@54260.4]
  wire  RetimeWrapper_185_io_out; // @[package.scala 93:22:@54260.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@54268.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@54268.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@54268.4]
  wire  RetimeWrapper_186_io_in; // @[package.scala 93:22:@54268.4]
  wire  RetimeWrapper_186_io_out; // @[package.scala 93:22:@54268.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@54276.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@54276.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@54276.4]
  wire  RetimeWrapper_187_io_in; // @[package.scala 93:22:@54276.4]
  wire  RetimeWrapper_187_io_out; // @[package.scala 93:22:@54276.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@54284.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@54284.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@54284.4]
  wire  RetimeWrapper_188_io_in; // @[package.scala 93:22:@54284.4]
  wire  RetimeWrapper_188_io_out; // @[package.scala 93:22:@54284.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@54292.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@54292.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@54292.4]
  wire  RetimeWrapper_189_io_in; // @[package.scala 93:22:@54292.4]
  wire  RetimeWrapper_189_io_out; // @[package.scala 93:22:@54292.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@54300.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@54300.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@54300.4]
  wire  RetimeWrapper_190_io_in; // @[package.scala 93:22:@54300.4]
  wire  RetimeWrapper_190_io_out; // @[package.scala 93:22:@54300.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@54308.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@54308.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@54308.4]
  wire  RetimeWrapper_191_io_in; // @[package.scala 93:22:@54308.4]
  wire  RetimeWrapper_191_io_out; // @[package.scala 93:22:@54308.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@54316.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@54316.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@54316.4]
  wire  RetimeWrapper_192_io_in; // @[package.scala 93:22:@54316.4]
  wire  RetimeWrapper_192_io_out; // @[package.scala 93:22:@54316.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@54324.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@54324.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@54324.4]
  wire  RetimeWrapper_193_io_in; // @[package.scala 93:22:@54324.4]
  wire  RetimeWrapper_193_io_out; // @[package.scala 93:22:@54324.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@54332.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@54332.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@54332.4]
  wire  RetimeWrapper_194_io_in; // @[package.scala 93:22:@54332.4]
  wire  RetimeWrapper_194_io_out; // @[package.scala 93:22:@54332.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@54340.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@54340.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@54340.4]
  wire  RetimeWrapper_195_io_in; // @[package.scala 93:22:@54340.4]
  wire  RetimeWrapper_195_io_out; // @[package.scala 93:22:@54340.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@54348.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@54348.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@54348.4]
  wire  RetimeWrapper_196_io_in; // @[package.scala 93:22:@54348.4]
  wire  RetimeWrapper_196_io_out; // @[package.scala 93:22:@54348.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@54356.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@54356.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@54356.4]
  wire  RetimeWrapper_197_io_in; // @[package.scala 93:22:@54356.4]
  wire  RetimeWrapper_197_io_out; // @[package.scala 93:22:@54356.4]
  wire  RetimeWrapper_198_clock; // @[package.scala 93:22:@54364.4]
  wire  RetimeWrapper_198_reset; // @[package.scala 93:22:@54364.4]
  wire  RetimeWrapper_198_io_flow; // @[package.scala 93:22:@54364.4]
  wire  RetimeWrapper_198_io_in; // @[package.scala 93:22:@54364.4]
  wire  RetimeWrapper_198_io_out; // @[package.scala 93:22:@54364.4]
  wire  RetimeWrapper_199_clock; // @[package.scala 93:22:@54372.4]
  wire  RetimeWrapper_199_reset; // @[package.scala 93:22:@54372.4]
  wire  RetimeWrapper_199_io_flow; // @[package.scala 93:22:@54372.4]
  wire  RetimeWrapper_199_io_in; // @[package.scala 93:22:@54372.4]
  wire  RetimeWrapper_199_io_out; // @[package.scala 93:22:@54372.4]
  wire  RetimeWrapper_200_clock; // @[package.scala 93:22:@54460.4]
  wire  RetimeWrapper_200_reset; // @[package.scala 93:22:@54460.4]
  wire  RetimeWrapper_200_io_flow; // @[package.scala 93:22:@54460.4]
  wire  RetimeWrapper_200_io_in; // @[package.scala 93:22:@54460.4]
  wire  RetimeWrapper_200_io_out; // @[package.scala 93:22:@54460.4]
  wire  RetimeWrapper_201_clock; // @[package.scala 93:22:@54468.4]
  wire  RetimeWrapper_201_reset; // @[package.scala 93:22:@54468.4]
  wire  RetimeWrapper_201_io_flow; // @[package.scala 93:22:@54468.4]
  wire  RetimeWrapper_201_io_in; // @[package.scala 93:22:@54468.4]
  wire  RetimeWrapper_201_io_out; // @[package.scala 93:22:@54468.4]
  wire  RetimeWrapper_202_clock; // @[package.scala 93:22:@54476.4]
  wire  RetimeWrapper_202_reset; // @[package.scala 93:22:@54476.4]
  wire  RetimeWrapper_202_io_flow; // @[package.scala 93:22:@54476.4]
  wire  RetimeWrapper_202_io_in; // @[package.scala 93:22:@54476.4]
  wire  RetimeWrapper_202_io_out; // @[package.scala 93:22:@54476.4]
  wire  RetimeWrapper_203_clock; // @[package.scala 93:22:@54484.4]
  wire  RetimeWrapper_203_reset; // @[package.scala 93:22:@54484.4]
  wire  RetimeWrapper_203_io_flow; // @[package.scala 93:22:@54484.4]
  wire  RetimeWrapper_203_io_in; // @[package.scala 93:22:@54484.4]
  wire  RetimeWrapper_203_io_out; // @[package.scala 93:22:@54484.4]
  wire  RetimeWrapper_204_clock; // @[package.scala 93:22:@54492.4]
  wire  RetimeWrapper_204_reset; // @[package.scala 93:22:@54492.4]
  wire  RetimeWrapper_204_io_flow; // @[package.scala 93:22:@54492.4]
  wire  RetimeWrapper_204_io_in; // @[package.scala 93:22:@54492.4]
  wire  RetimeWrapper_204_io_out; // @[package.scala 93:22:@54492.4]
  wire  RetimeWrapper_205_clock; // @[package.scala 93:22:@54500.4]
  wire  RetimeWrapper_205_reset; // @[package.scala 93:22:@54500.4]
  wire  RetimeWrapper_205_io_flow; // @[package.scala 93:22:@54500.4]
  wire  RetimeWrapper_205_io_in; // @[package.scala 93:22:@54500.4]
  wire  RetimeWrapper_205_io_out; // @[package.scala 93:22:@54500.4]
  wire  RetimeWrapper_206_clock; // @[package.scala 93:22:@54508.4]
  wire  RetimeWrapper_206_reset; // @[package.scala 93:22:@54508.4]
  wire  RetimeWrapper_206_io_flow; // @[package.scala 93:22:@54508.4]
  wire  RetimeWrapper_206_io_in; // @[package.scala 93:22:@54508.4]
  wire  RetimeWrapper_206_io_out; // @[package.scala 93:22:@54508.4]
  wire  RetimeWrapper_207_clock; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_207_reset; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_207_io_flow; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_207_io_in; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_207_io_out; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_208_clock; // @[package.scala 93:22:@54524.4]
  wire  RetimeWrapper_208_reset; // @[package.scala 93:22:@54524.4]
  wire  RetimeWrapper_208_io_flow; // @[package.scala 93:22:@54524.4]
  wire  RetimeWrapper_208_io_in; // @[package.scala 93:22:@54524.4]
  wire  RetimeWrapper_208_io_out; // @[package.scala 93:22:@54524.4]
  wire  RetimeWrapper_209_clock; // @[package.scala 93:22:@54532.4]
  wire  RetimeWrapper_209_reset; // @[package.scala 93:22:@54532.4]
  wire  RetimeWrapper_209_io_flow; // @[package.scala 93:22:@54532.4]
  wire  RetimeWrapper_209_io_in; // @[package.scala 93:22:@54532.4]
  wire  RetimeWrapper_209_io_out; // @[package.scala 93:22:@54532.4]
  wire  RetimeWrapper_210_clock; // @[package.scala 93:22:@54540.4]
  wire  RetimeWrapper_210_reset; // @[package.scala 93:22:@54540.4]
  wire  RetimeWrapper_210_io_flow; // @[package.scala 93:22:@54540.4]
  wire  RetimeWrapper_210_io_in; // @[package.scala 93:22:@54540.4]
  wire  RetimeWrapper_210_io_out; // @[package.scala 93:22:@54540.4]
  wire  RetimeWrapper_211_clock; // @[package.scala 93:22:@54548.4]
  wire  RetimeWrapper_211_reset; // @[package.scala 93:22:@54548.4]
  wire  RetimeWrapper_211_io_flow; // @[package.scala 93:22:@54548.4]
  wire  RetimeWrapper_211_io_in; // @[package.scala 93:22:@54548.4]
  wire  RetimeWrapper_211_io_out; // @[package.scala 93:22:@54548.4]
  wire  RetimeWrapper_212_clock; // @[package.scala 93:22:@54556.4]
  wire  RetimeWrapper_212_reset; // @[package.scala 93:22:@54556.4]
  wire  RetimeWrapper_212_io_flow; // @[package.scala 93:22:@54556.4]
  wire  RetimeWrapper_212_io_in; // @[package.scala 93:22:@54556.4]
  wire  RetimeWrapper_212_io_out; // @[package.scala 93:22:@54556.4]
  wire  RetimeWrapper_213_clock; // @[package.scala 93:22:@54564.4]
  wire  RetimeWrapper_213_reset; // @[package.scala 93:22:@54564.4]
  wire  RetimeWrapper_213_io_flow; // @[package.scala 93:22:@54564.4]
  wire  RetimeWrapper_213_io_in; // @[package.scala 93:22:@54564.4]
  wire  RetimeWrapper_213_io_out; // @[package.scala 93:22:@54564.4]
  wire  RetimeWrapper_214_clock; // @[package.scala 93:22:@54572.4]
  wire  RetimeWrapper_214_reset; // @[package.scala 93:22:@54572.4]
  wire  RetimeWrapper_214_io_flow; // @[package.scala 93:22:@54572.4]
  wire  RetimeWrapper_214_io_in; // @[package.scala 93:22:@54572.4]
  wire  RetimeWrapper_214_io_out; // @[package.scala 93:22:@54572.4]
  wire  RetimeWrapper_215_clock; // @[package.scala 93:22:@54580.4]
  wire  RetimeWrapper_215_reset; // @[package.scala 93:22:@54580.4]
  wire  RetimeWrapper_215_io_flow; // @[package.scala 93:22:@54580.4]
  wire  RetimeWrapper_215_io_in; // @[package.scala 93:22:@54580.4]
  wire  RetimeWrapper_215_io_out; // @[package.scala 93:22:@54580.4]
  wire  RetimeWrapper_216_clock; // @[package.scala 93:22:@54588.4]
  wire  RetimeWrapper_216_reset; // @[package.scala 93:22:@54588.4]
  wire  RetimeWrapper_216_io_flow; // @[package.scala 93:22:@54588.4]
  wire  RetimeWrapper_216_io_in; // @[package.scala 93:22:@54588.4]
  wire  RetimeWrapper_216_io_out; // @[package.scala 93:22:@54588.4]
  wire  RetimeWrapper_217_clock; // @[package.scala 93:22:@54596.4]
  wire  RetimeWrapper_217_reset; // @[package.scala 93:22:@54596.4]
  wire  RetimeWrapper_217_io_flow; // @[package.scala 93:22:@54596.4]
  wire  RetimeWrapper_217_io_in; // @[package.scala 93:22:@54596.4]
  wire  RetimeWrapper_217_io_out; // @[package.scala 93:22:@54596.4]
  wire  RetimeWrapper_218_clock; // @[package.scala 93:22:@54604.4]
  wire  RetimeWrapper_218_reset; // @[package.scala 93:22:@54604.4]
  wire  RetimeWrapper_218_io_flow; // @[package.scala 93:22:@54604.4]
  wire  RetimeWrapper_218_io_in; // @[package.scala 93:22:@54604.4]
  wire  RetimeWrapper_218_io_out; // @[package.scala 93:22:@54604.4]
  wire  RetimeWrapper_219_clock; // @[package.scala 93:22:@54612.4]
  wire  RetimeWrapper_219_reset; // @[package.scala 93:22:@54612.4]
  wire  RetimeWrapper_219_io_flow; // @[package.scala 93:22:@54612.4]
  wire  RetimeWrapper_219_io_in; // @[package.scala 93:22:@54612.4]
  wire  RetimeWrapper_219_io_out; // @[package.scala 93:22:@54612.4]
  wire  RetimeWrapper_220_clock; // @[package.scala 93:22:@54700.4]
  wire  RetimeWrapper_220_reset; // @[package.scala 93:22:@54700.4]
  wire  RetimeWrapper_220_io_flow; // @[package.scala 93:22:@54700.4]
  wire  RetimeWrapper_220_io_in; // @[package.scala 93:22:@54700.4]
  wire  RetimeWrapper_220_io_out; // @[package.scala 93:22:@54700.4]
  wire  RetimeWrapper_221_clock; // @[package.scala 93:22:@54708.4]
  wire  RetimeWrapper_221_reset; // @[package.scala 93:22:@54708.4]
  wire  RetimeWrapper_221_io_flow; // @[package.scala 93:22:@54708.4]
  wire  RetimeWrapper_221_io_in; // @[package.scala 93:22:@54708.4]
  wire  RetimeWrapper_221_io_out; // @[package.scala 93:22:@54708.4]
  wire  RetimeWrapper_222_clock; // @[package.scala 93:22:@54716.4]
  wire  RetimeWrapper_222_reset; // @[package.scala 93:22:@54716.4]
  wire  RetimeWrapper_222_io_flow; // @[package.scala 93:22:@54716.4]
  wire  RetimeWrapper_222_io_in; // @[package.scala 93:22:@54716.4]
  wire  RetimeWrapper_222_io_out; // @[package.scala 93:22:@54716.4]
  wire  RetimeWrapper_223_clock; // @[package.scala 93:22:@54724.4]
  wire  RetimeWrapper_223_reset; // @[package.scala 93:22:@54724.4]
  wire  RetimeWrapper_223_io_flow; // @[package.scala 93:22:@54724.4]
  wire  RetimeWrapper_223_io_in; // @[package.scala 93:22:@54724.4]
  wire  RetimeWrapper_223_io_out; // @[package.scala 93:22:@54724.4]
  wire  RetimeWrapper_224_clock; // @[package.scala 93:22:@54732.4]
  wire  RetimeWrapper_224_reset; // @[package.scala 93:22:@54732.4]
  wire  RetimeWrapper_224_io_flow; // @[package.scala 93:22:@54732.4]
  wire  RetimeWrapper_224_io_in; // @[package.scala 93:22:@54732.4]
  wire  RetimeWrapper_224_io_out; // @[package.scala 93:22:@54732.4]
  wire  RetimeWrapper_225_clock; // @[package.scala 93:22:@54740.4]
  wire  RetimeWrapper_225_reset; // @[package.scala 93:22:@54740.4]
  wire  RetimeWrapper_225_io_flow; // @[package.scala 93:22:@54740.4]
  wire  RetimeWrapper_225_io_in; // @[package.scala 93:22:@54740.4]
  wire  RetimeWrapper_225_io_out; // @[package.scala 93:22:@54740.4]
  wire  RetimeWrapper_226_clock; // @[package.scala 93:22:@54748.4]
  wire  RetimeWrapper_226_reset; // @[package.scala 93:22:@54748.4]
  wire  RetimeWrapper_226_io_flow; // @[package.scala 93:22:@54748.4]
  wire  RetimeWrapper_226_io_in; // @[package.scala 93:22:@54748.4]
  wire  RetimeWrapper_226_io_out; // @[package.scala 93:22:@54748.4]
  wire  RetimeWrapper_227_clock; // @[package.scala 93:22:@54756.4]
  wire  RetimeWrapper_227_reset; // @[package.scala 93:22:@54756.4]
  wire  RetimeWrapper_227_io_flow; // @[package.scala 93:22:@54756.4]
  wire  RetimeWrapper_227_io_in; // @[package.scala 93:22:@54756.4]
  wire  RetimeWrapper_227_io_out; // @[package.scala 93:22:@54756.4]
  wire  RetimeWrapper_228_clock; // @[package.scala 93:22:@54764.4]
  wire  RetimeWrapper_228_reset; // @[package.scala 93:22:@54764.4]
  wire  RetimeWrapper_228_io_flow; // @[package.scala 93:22:@54764.4]
  wire  RetimeWrapper_228_io_in; // @[package.scala 93:22:@54764.4]
  wire  RetimeWrapper_228_io_out; // @[package.scala 93:22:@54764.4]
  wire  RetimeWrapper_229_clock; // @[package.scala 93:22:@54772.4]
  wire  RetimeWrapper_229_reset; // @[package.scala 93:22:@54772.4]
  wire  RetimeWrapper_229_io_flow; // @[package.scala 93:22:@54772.4]
  wire  RetimeWrapper_229_io_in; // @[package.scala 93:22:@54772.4]
  wire  RetimeWrapper_229_io_out; // @[package.scala 93:22:@54772.4]
  wire  RetimeWrapper_230_clock; // @[package.scala 93:22:@54780.4]
  wire  RetimeWrapper_230_reset; // @[package.scala 93:22:@54780.4]
  wire  RetimeWrapper_230_io_flow; // @[package.scala 93:22:@54780.4]
  wire  RetimeWrapper_230_io_in; // @[package.scala 93:22:@54780.4]
  wire  RetimeWrapper_230_io_out; // @[package.scala 93:22:@54780.4]
  wire  RetimeWrapper_231_clock; // @[package.scala 93:22:@54788.4]
  wire  RetimeWrapper_231_reset; // @[package.scala 93:22:@54788.4]
  wire  RetimeWrapper_231_io_flow; // @[package.scala 93:22:@54788.4]
  wire  RetimeWrapper_231_io_in; // @[package.scala 93:22:@54788.4]
  wire  RetimeWrapper_231_io_out; // @[package.scala 93:22:@54788.4]
  wire  RetimeWrapper_232_clock; // @[package.scala 93:22:@54796.4]
  wire  RetimeWrapper_232_reset; // @[package.scala 93:22:@54796.4]
  wire  RetimeWrapper_232_io_flow; // @[package.scala 93:22:@54796.4]
  wire  RetimeWrapper_232_io_in; // @[package.scala 93:22:@54796.4]
  wire  RetimeWrapper_232_io_out; // @[package.scala 93:22:@54796.4]
  wire  RetimeWrapper_233_clock; // @[package.scala 93:22:@54804.4]
  wire  RetimeWrapper_233_reset; // @[package.scala 93:22:@54804.4]
  wire  RetimeWrapper_233_io_flow; // @[package.scala 93:22:@54804.4]
  wire  RetimeWrapper_233_io_in; // @[package.scala 93:22:@54804.4]
  wire  RetimeWrapper_233_io_out; // @[package.scala 93:22:@54804.4]
  wire  RetimeWrapper_234_clock; // @[package.scala 93:22:@54812.4]
  wire  RetimeWrapper_234_reset; // @[package.scala 93:22:@54812.4]
  wire  RetimeWrapper_234_io_flow; // @[package.scala 93:22:@54812.4]
  wire  RetimeWrapper_234_io_in; // @[package.scala 93:22:@54812.4]
  wire  RetimeWrapper_234_io_out; // @[package.scala 93:22:@54812.4]
  wire  RetimeWrapper_235_clock; // @[package.scala 93:22:@54820.4]
  wire  RetimeWrapper_235_reset; // @[package.scala 93:22:@54820.4]
  wire  RetimeWrapper_235_io_flow; // @[package.scala 93:22:@54820.4]
  wire  RetimeWrapper_235_io_in; // @[package.scala 93:22:@54820.4]
  wire  RetimeWrapper_235_io_out; // @[package.scala 93:22:@54820.4]
  wire  RetimeWrapper_236_clock; // @[package.scala 93:22:@54828.4]
  wire  RetimeWrapper_236_reset; // @[package.scala 93:22:@54828.4]
  wire  RetimeWrapper_236_io_flow; // @[package.scala 93:22:@54828.4]
  wire  RetimeWrapper_236_io_in; // @[package.scala 93:22:@54828.4]
  wire  RetimeWrapper_236_io_out; // @[package.scala 93:22:@54828.4]
  wire  RetimeWrapper_237_clock; // @[package.scala 93:22:@54836.4]
  wire  RetimeWrapper_237_reset; // @[package.scala 93:22:@54836.4]
  wire  RetimeWrapper_237_io_flow; // @[package.scala 93:22:@54836.4]
  wire  RetimeWrapper_237_io_in; // @[package.scala 93:22:@54836.4]
  wire  RetimeWrapper_237_io_out; // @[package.scala 93:22:@54836.4]
  wire  RetimeWrapper_238_clock; // @[package.scala 93:22:@54844.4]
  wire  RetimeWrapper_238_reset; // @[package.scala 93:22:@54844.4]
  wire  RetimeWrapper_238_io_flow; // @[package.scala 93:22:@54844.4]
  wire  RetimeWrapper_238_io_in; // @[package.scala 93:22:@54844.4]
  wire  RetimeWrapper_238_io_out; // @[package.scala 93:22:@54844.4]
  wire  RetimeWrapper_239_clock; // @[package.scala 93:22:@54852.4]
  wire  RetimeWrapper_239_reset; // @[package.scala 93:22:@54852.4]
  wire  RetimeWrapper_239_io_flow; // @[package.scala 93:22:@54852.4]
  wire  RetimeWrapper_239_io_in; // @[package.scala 93:22:@54852.4]
  wire  RetimeWrapper_239_io_out; // @[package.scala 93:22:@54852.4]
  wire  RetimeWrapper_240_clock; // @[package.scala 93:22:@54940.4]
  wire  RetimeWrapper_240_reset; // @[package.scala 93:22:@54940.4]
  wire  RetimeWrapper_240_io_flow; // @[package.scala 93:22:@54940.4]
  wire  RetimeWrapper_240_io_in; // @[package.scala 93:22:@54940.4]
  wire  RetimeWrapper_240_io_out; // @[package.scala 93:22:@54940.4]
  wire  RetimeWrapper_241_clock; // @[package.scala 93:22:@54948.4]
  wire  RetimeWrapper_241_reset; // @[package.scala 93:22:@54948.4]
  wire  RetimeWrapper_241_io_flow; // @[package.scala 93:22:@54948.4]
  wire  RetimeWrapper_241_io_in; // @[package.scala 93:22:@54948.4]
  wire  RetimeWrapper_241_io_out; // @[package.scala 93:22:@54948.4]
  wire  RetimeWrapper_242_clock; // @[package.scala 93:22:@54956.4]
  wire  RetimeWrapper_242_reset; // @[package.scala 93:22:@54956.4]
  wire  RetimeWrapper_242_io_flow; // @[package.scala 93:22:@54956.4]
  wire  RetimeWrapper_242_io_in; // @[package.scala 93:22:@54956.4]
  wire  RetimeWrapper_242_io_out; // @[package.scala 93:22:@54956.4]
  wire  RetimeWrapper_243_clock; // @[package.scala 93:22:@54964.4]
  wire  RetimeWrapper_243_reset; // @[package.scala 93:22:@54964.4]
  wire  RetimeWrapper_243_io_flow; // @[package.scala 93:22:@54964.4]
  wire  RetimeWrapper_243_io_in; // @[package.scala 93:22:@54964.4]
  wire  RetimeWrapper_243_io_out; // @[package.scala 93:22:@54964.4]
  wire  RetimeWrapper_244_clock; // @[package.scala 93:22:@54972.4]
  wire  RetimeWrapper_244_reset; // @[package.scala 93:22:@54972.4]
  wire  RetimeWrapper_244_io_flow; // @[package.scala 93:22:@54972.4]
  wire  RetimeWrapper_244_io_in; // @[package.scala 93:22:@54972.4]
  wire  RetimeWrapper_244_io_out; // @[package.scala 93:22:@54972.4]
  wire  RetimeWrapper_245_clock; // @[package.scala 93:22:@54980.4]
  wire  RetimeWrapper_245_reset; // @[package.scala 93:22:@54980.4]
  wire  RetimeWrapper_245_io_flow; // @[package.scala 93:22:@54980.4]
  wire  RetimeWrapper_245_io_in; // @[package.scala 93:22:@54980.4]
  wire  RetimeWrapper_245_io_out; // @[package.scala 93:22:@54980.4]
  wire  RetimeWrapper_246_clock; // @[package.scala 93:22:@54988.4]
  wire  RetimeWrapper_246_reset; // @[package.scala 93:22:@54988.4]
  wire  RetimeWrapper_246_io_flow; // @[package.scala 93:22:@54988.4]
  wire  RetimeWrapper_246_io_in; // @[package.scala 93:22:@54988.4]
  wire  RetimeWrapper_246_io_out; // @[package.scala 93:22:@54988.4]
  wire  RetimeWrapper_247_clock; // @[package.scala 93:22:@54996.4]
  wire  RetimeWrapper_247_reset; // @[package.scala 93:22:@54996.4]
  wire  RetimeWrapper_247_io_flow; // @[package.scala 93:22:@54996.4]
  wire  RetimeWrapper_247_io_in; // @[package.scala 93:22:@54996.4]
  wire  RetimeWrapper_247_io_out; // @[package.scala 93:22:@54996.4]
  wire  RetimeWrapper_248_clock; // @[package.scala 93:22:@55004.4]
  wire  RetimeWrapper_248_reset; // @[package.scala 93:22:@55004.4]
  wire  RetimeWrapper_248_io_flow; // @[package.scala 93:22:@55004.4]
  wire  RetimeWrapper_248_io_in; // @[package.scala 93:22:@55004.4]
  wire  RetimeWrapper_248_io_out; // @[package.scala 93:22:@55004.4]
  wire  RetimeWrapper_249_clock; // @[package.scala 93:22:@55012.4]
  wire  RetimeWrapper_249_reset; // @[package.scala 93:22:@55012.4]
  wire  RetimeWrapper_249_io_flow; // @[package.scala 93:22:@55012.4]
  wire  RetimeWrapper_249_io_in; // @[package.scala 93:22:@55012.4]
  wire  RetimeWrapper_249_io_out; // @[package.scala 93:22:@55012.4]
  wire  RetimeWrapper_250_clock; // @[package.scala 93:22:@55020.4]
  wire  RetimeWrapper_250_reset; // @[package.scala 93:22:@55020.4]
  wire  RetimeWrapper_250_io_flow; // @[package.scala 93:22:@55020.4]
  wire  RetimeWrapper_250_io_in; // @[package.scala 93:22:@55020.4]
  wire  RetimeWrapper_250_io_out; // @[package.scala 93:22:@55020.4]
  wire  RetimeWrapper_251_clock; // @[package.scala 93:22:@55028.4]
  wire  RetimeWrapper_251_reset; // @[package.scala 93:22:@55028.4]
  wire  RetimeWrapper_251_io_flow; // @[package.scala 93:22:@55028.4]
  wire  RetimeWrapper_251_io_in; // @[package.scala 93:22:@55028.4]
  wire  RetimeWrapper_251_io_out; // @[package.scala 93:22:@55028.4]
  wire  RetimeWrapper_252_clock; // @[package.scala 93:22:@55036.4]
  wire  RetimeWrapper_252_reset; // @[package.scala 93:22:@55036.4]
  wire  RetimeWrapper_252_io_flow; // @[package.scala 93:22:@55036.4]
  wire  RetimeWrapper_252_io_in; // @[package.scala 93:22:@55036.4]
  wire  RetimeWrapper_252_io_out; // @[package.scala 93:22:@55036.4]
  wire  RetimeWrapper_253_clock; // @[package.scala 93:22:@55044.4]
  wire  RetimeWrapper_253_reset; // @[package.scala 93:22:@55044.4]
  wire  RetimeWrapper_253_io_flow; // @[package.scala 93:22:@55044.4]
  wire  RetimeWrapper_253_io_in; // @[package.scala 93:22:@55044.4]
  wire  RetimeWrapper_253_io_out; // @[package.scala 93:22:@55044.4]
  wire  RetimeWrapper_254_clock; // @[package.scala 93:22:@55052.4]
  wire  RetimeWrapper_254_reset; // @[package.scala 93:22:@55052.4]
  wire  RetimeWrapper_254_io_flow; // @[package.scala 93:22:@55052.4]
  wire  RetimeWrapper_254_io_in; // @[package.scala 93:22:@55052.4]
  wire  RetimeWrapper_254_io_out; // @[package.scala 93:22:@55052.4]
  wire  RetimeWrapper_255_clock; // @[package.scala 93:22:@55060.4]
  wire  RetimeWrapper_255_reset; // @[package.scala 93:22:@55060.4]
  wire  RetimeWrapper_255_io_flow; // @[package.scala 93:22:@55060.4]
  wire  RetimeWrapper_255_io_in; // @[package.scala 93:22:@55060.4]
  wire  RetimeWrapper_255_io_out; // @[package.scala 93:22:@55060.4]
  wire  RetimeWrapper_256_clock; // @[package.scala 93:22:@55068.4]
  wire  RetimeWrapper_256_reset; // @[package.scala 93:22:@55068.4]
  wire  RetimeWrapper_256_io_flow; // @[package.scala 93:22:@55068.4]
  wire  RetimeWrapper_256_io_in; // @[package.scala 93:22:@55068.4]
  wire  RetimeWrapper_256_io_out; // @[package.scala 93:22:@55068.4]
  wire  RetimeWrapper_257_clock; // @[package.scala 93:22:@55076.4]
  wire  RetimeWrapper_257_reset; // @[package.scala 93:22:@55076.4]
  wire  RetimeWrapper_257_io_flow; // @[package.scala 93:22:@55076.4]
  wire  RetimeWrapper_257_io_in; // @[package.scala 93:22:@55076.4]
  wire  RetimeWrapper_257_io_out; // @[package.scala 93:22:@55076.4]
  wire  RetimeWrapper_258_clock; // @[package.scala 93:22:@55084.4]
  wire  RetimeWrapper_258_reset; // @[package.scala 93:22:@55084.4]
  wire  RetimeWrapper_258_io_flow; // @[package.scala 93:22:@55084.4]
  wire  RetimeWrapper_258_io_in; // @[package.scala 93:22:@55084.4]
  wire  RetimeWrapper_258_io_out; // @[package.scala 93:22:@55084.4]
  wire  RetimeWrapper_259_clock; // @[package.scala 93:22:@55092.4]
  wire  RetimeWrapper_259_reset; // @[package.scala 93:22:@55092.4]
  wire  RetimeWrapper_259_io_flow; // @[package.scala 93:22:@55092.4]
  wire  RetimeWrapper_259_io_in; // @[package.scala 93:22:@55092.4]
  wire  RetimeWrapper_259_io_out; // @[package.scala 93:22:@55092.4]
  wire  RetimeWrapper_260_clock; // @[package.scala 93:22:@55180.4]
  wire  RetimeWrapper_260_reset; // @[package.scala 93:22:@55180.4]
  wire  RetimeWrapper_260_io_flow; // @[package.scala 93:22:@55180.4]
  wire  RetimeWrapper_260_io_in; // @[package.scala 93:22:@55180.4]
  wire  RetimeWrapper_260_io_out; // @[package.scala 93:22:@55180.4]
  wire  RetimeWrapper_261_clock; // @[package.scala 93:22:@55188.4]
  wire  RetimeWrapper_261_reset; // @[package.scala 93:22:@55188.4]
  wire  RetimeWrapper_261_io_flow; // @[package.scala 93:22:@55188.4]
  wire  RetimeWrapper_261_io_in; // @[package.scala 93:22:@55188.4]
  wire  RetimeWrapper_261_io_out; // @[package.scala 93:22:@55188.4]
  wire  RetimeWrapper_262_clock; // @[package.scala 93:22:@55196.4]
  wire  RetimeWrapper_262_reset; // @[package.scala 93:22:@55196.4]
  wire  RetimeWrapper_262_io_flow; // @[package.scala 93:22:@55196.4]
  wire  RetimeWrapper_262_io_in; // @[package.scala 93:22:@55196.4]
  wire  RetimeWrapper_262_io_out; // @[package.scala 93:22:@55196.4]
  wire  RetimeWrapper_263_clock; // @[package.scala 93:22:@55204.4]
  wire  RetimeWrapper_263_reset; // @[package.scala 93:22:@55204.4]
  wire  RetimeWrapper_263_io_flow; // @[package.scala 93:22:@55204.4]
  wire  RetimeWrapper_263_io_in; // @[package.scala 93:22:@55204.4]
  wire  RetimeWrapper_263_io_out; // @[package.scala 93:22:@55204.4]
  wire  RetimeWrapper_264_clock; // @[package.scala 93:22:@55212.4]
  wire  RetimeWrapper_264_reset; // @[package.scala 93:22:@55212.4]
  wire  RetimeWrapper_264_io_flow; // @[package.scala 93:22:@55212.4]
  wire  RetimeWrapper_264_io_in; // @[package.scala 93:22:@55212.4]
  wire  RetimeWrapper_264_io_out; // @[package.scala 93:22:@55212.4]
  wire  RetimeWrapper_265_clock; // @[package.scala 93:22:@55220.4]
  wire  RetimeWrapper_265_reset; // @[package.scala 93:22:@55220.4]
  wire  RetimeWrapper_265_io_flow; // @[package.scala 93:22:@55220.4]
  wire  RetimeWrapper_265_io_in; // @[package.scala 93:22:@55220.4]
  wire  RetimeWrapper_265_io_out; // @[package.scala 93:22:@55220.4]
  wire  RetimeWrapper_266_clock; // @[package.scala 93:22:@55228.4]
  wire  RetimeWrapper_266_reset; // @[package.scala 93:22:@55228.4]
  wire  RetimeWrapper_266_io_flow; // @[package.scala 93:22:@55228.4]
  wire  RetimeWrapper_266_io_in; // @[package.scala 93:22:@55228.4]
  wire  RetimeWrapper_266_io_out; // @[package.scala 93:22:@55228.4]
  wire  RetimeWrapper_267_clock; // @[package.scala 93:22:@55236.4]
  wire  RetimeWrapper_267_reset; // @[package.scala 93:22:@55236.4]
  wire  RetimeWrapper_267_io_flow; // @[package.scala 93:22:@55236.4]
  wire  RetimeWrapper_267_io_in; // @[package.scala 93:22:@55236.4]
  wire  RetimeWrapper_267_io_out; // @[package.scala 93:22:@55236.4]
  wire  RetimeWrapper_268_clock; // @[package.scala 93:22:@55244.4]
  wire  RetimeWrapper_268_reset; // @[package.scala 93:22:@55244.4]
  wire  RetimeWrapper_268_io_flow; // @[package.scala 93:22:@55244.4]
  wire  RetimeWrapper_268_io_in; // @[package.scala 93:22:@55244.4]
  wire  RetimeWrapper_268_io_out; // @[package.scala 93:22:@55244.4]
  wire  RetimeWrapper_269_clock; // @[package.scala 93:22:@55252.4]
  wire  RetimeWrapper_269_reset; // @[package.scala 93:22:@55252.4]
  wire  RetimeWrapper_269_io_flow; // @[package.scala 93:22:@55252.4]
  wire  RetimeWrapper_269_io_in; // @[package.scala 93:22:@55252.4]
  wire  RetimeWrapper_269_io_out; // @[package.scala 93:22:@55252.4]
  wire  RetimeWrapper_270_clock; // @[package.scala 93:22:@55260.4]
  wire  RetimeWrapper_270_reset; // @[package.scala 93:22:@55260.4]
  wire  RetimeWrapper_270_io_flow; // @[package.scala 93:22:@55260.4]
  wire  RetimeWrapper_270_io_in; // @[package.scala 93:22:@55260.4]
  wire  RetimeWrapper_270_io_out; // @[package.scala 93:22:@55260.4]
  wire  RetimeWrapper_271_clock; // @[package.scala 93:22:@55268.4]
  wire  RetimeWrapper_271_reset; // @[package.scala 93:22:@55268.4]
  wire  RetimeWrapper_271_io_flow; // @[package.scala 93:22:@55268.4]
  wire  RetimeWrapper_271_io_in; // @[package.scala 93:22:@55268.4]
  wire  RetimeWrapper_271_io_out; // @[package.scala 93:22:@55268.4]
  wire  RetimeWrapper_272_clock; // @[package.scala 93:22:@55276.4]
  wire  RetimeWrapper_272_reset; // @[package.scala 93:22:@55276.4]
  wire  RetimeWrapper_272_io_flow; // @[package.scala 93:22:@55276.4]
  wire  RetimeWrapper_272_io_in; // @[package.scala 93:22:@55276.4]
  wire  RetimeWrapper_272_io_out; // @[package.scala 93:22:@55276.4]
  wire  RetimeWrapper_273_clock; // @[package.scala 93:22:@55284.4]
  wire  RetimeWrapper_273_reset; // @[package.scala 93:22:@55284.4]
  wire  RetimeWrapper_273_io_flow; // @[package.scala 93:22:@55284.4]
  wire  RetimeWrapper_273_io_in; // @[package.scala 93:22:@55284.4]
  wire  RetimeWrapper_273_io_out; // @[package.scala 93:22:@55284.4]
  wire  RetimeWrapper_274_clock; // @[package.scala 93:22:@55292.4]
  wire  RetimeWrapper_274_reset; // @[package.scala 93:22:@55292.4]
  wire  RetimeWrapper_274_io_flow; // @[package.scala 93:22:@55292.4]
  wire  RetimeWrapper_274_io_in; // @[package.scala 93:22:@55292.4]
  wire  RetimeWrapper_274_io_out; // @[package.scala 93:22:@55292.4]
  wire  RetimeWrapper_275_clock; // @[package.scala 93:22:@55300.4]
  wire  RetimeWrapper_275_reset; // @[package.scala 93:22:@55300.4]
  wire  RetimeWrapper_275_io_flow; // @[package.scala 93:22:@55300.4]
  wire  RetimeWrapper_275_io_in; // @[package.scala 93:22:@55300.4]
  wire  RetimeWrapper_275_io_out; // @[package.scala 93:22:@55300.4]
  wire  RetimeWrapper_276_clock; // @[package.scala 93:22:@55308.4]
  wire  RetimeWrapper_276_reset; // @[package.scala 93:22:@55308.4]
  wire  RetimeWrapper_276_io_flow; // @[package.scala 93:22:@55308.4]
  wire  RetimeWrapper_276_io_in; // @[package.scala 93:22:@55308.4]
  wire  RetimeWrapper_276_io_out; // @[package.scala 93:22:@55308.4]
  wire  RetimeWrapper_277_clock; // @[package.scala 93:22:@55316.4]
  wire  RetimeWrapper_277_reset; // @[package.scala 93:22:@55316.4]
  wire  RetimeWrapper_277_io_flow; // @[package.scala 93:22:@55316.4]
  wire  RetimeWrapper_277_io_in; // @[package.scala 93:22:@55316.4]
  wire  RetimeWrapper_277_io_out; // @[package.scala 93:22:@55316.4]
  wire  RetimeWrapper_278_clock; // @[package.scala 93:22:@55324.4]
  wire  RetimeWrapper_278_reset; // @[package.scala 93:22:@55324.4]
  wire  RetimeWrapper_278_io_flow; // @[package.scala 93:22:@55324.4]
  wire  RetimeWrapper_278_io_in; // @[package.scala 93:22:@55324.4]
  wire  RetimeWrapper_278_io_out; // @[package.scala 93:22:@55324.4]
  wire  RetimeWrapper_279_clock; // @[package.scala 93:22:@55332.4]
  wire  RetimeWrapper_279_reset; // @[package.scala 93:22:@55332.4]
  wire  RetimeWrapper_279_io_flow; // @[package.scala 93:22:@55332.4]
  wire  RetimeWrapper_279_io_in; // @[package.scala 93:22:@55332.4]
  wire  RetimeWrapper_279_io_out; // @[package.scala 93:22:@55332.4]
  wire  RetimeWrapper_280_clock; // @[package.scala 93:22:@55420.4]
  wire  RetimeWrapper_280_reset; // @[package.scala 93:22:@55420.4]
  wire  RetimeWrapper_280_io_flow; // @[package.scala 93:22:@55420.4]
  wire  RetimeWrapper_280_io_in; // @[package.scala 93:22:@55420.4]
  wire  RetimeWrapper_280_io_out; // @[package.scala 93:22:@55420.4]
  wire  RetimeWrapper_281_clock; // @[package.scala 93:22:@55428.4]
  wire  RetimeWrapper_281_reset; // @[package.scala 93:22:@55428.4]
  wire  RetimeWrapper_281_io_flow; // @[package.scala 93:22:@55428.4]
  wire  RetimeWrapper_281_io_in; // @[package.scala 93:22:@55428.4]
  wire  RetimeWrapper_281_io_out; // @[package.scala 93:22:@55428.4]
  wire  RetimeWrapper_282_clock; // @[package.scala 93:22:@55436.4]
  wire  RetimeWrapper_282_reset; // @[package.scala 93:22:@55436.4]
  wire  RetimeWrapper_282_io_flow; // @[package.scala 93:22:@55436.4]
  wire  RetimeWrapper_282_io_in; // @[package.scala 93:22:@55436.4]
  wire  RetimeWrapper_282_io_out; // @[package.scala 93:22:@55436.4]
  wire  RetimeWrapper_283_clock; // @[package.scala 93:22:@55444.4]
  wire  RetimeWrapper_283_reset; // @[package.scala 93:22:@55444.4]
  wire  RetimeWrapper_283_io_flow; // @[package.scala 93:22:@55444.4]
  wire  RetimeWrapper_283_io_in; // @[package.scala 93:22:@55444.4]
  wire  RetimeWrapper_283_io_out; // @[package.scala 93:22:@55444.4]
  wire  RetimeWrapper_284_clock; // @[package.scala 93:22:@55452.4]
  wire  RetimeWrapper_284_reset; // @[package.scala 93:22:@55452.4]
  wire  RetimeWrapper_284_io_flow; // @[package.scala 93:22:@55452.4]
  wire  RetimeWrapper_284_io_in; // @[package.scala 93:22:@55452.4]
  wire  RetimeWrapper_284_io_out; // @[package.scala 93:22:@55452.4]
  wire  RetimeWrapper_285_clock; // @[package.scala 93:22:@55460.4]
  wire  RetimeWrapper_285_reset; // @[package.scala 93:22:@55460.4]
  wire  RetimeWrapper_285_io_flow; // @[package.scala 93:22:@55460.4]
  wire  RetimeWrapper_285_io_in; // @[package.scala 93:22:@55460.4]
  wire  RetimeWrapper_285_io_out; // @[package.scala 93:22:@55460.4]
  wire  RetimeWrapper_286_clock; // @[package.scala 93:22:@55468.4]
  wire  RetimeWrapper_286_reset; // @[package.scala 93:22:@55468.4]
  wire  RetimeWrapper_286_io_flow; // @[package.scala 93:22:@55468.4]
  wire  RetimeWrapper_286_io_in; // @[package.scala 93:22:@55468.4]
  wire  RetimeWrapper_286_io_out; // @[package.scala 93:22:@55468.4]
  wire  RetimeWrapper_287_clock; // @[package.scala 93:22:@55476.4]
  wire  RetimeWrapper_287_reset; // @[package.scala 93:22:@55476.4]
  wire  RetimeWrapper_287_io_flow; // @[package.scala 93:22:@55476.4]
  wire  RetimeWrapper_287_io_in; // @[package.scala 93:22:@55476.4]
  wire  RetimeWrapper_287_io_out; // @[package.scala 93:22:@55476.4]
  wire  RetimeWrapper_288_clock; // @[package.scala 93:22:@55484.4]
  wire  RetimeWrapper_288_reset; // @[package.scala 93:22:@55484.4]
  wire  RetimeWrapper_288_io_flow; // @[package.scala 93:22:@55484.4]
  wire  RetimeWrapper_288_io_in; // @[package.scala 93:22:@55484.4]
  wire  RetimeWrapper_288_io_out; // @[package.scala 93:22:@55484.4]
  wire  RetimeWrapper_289_clock; // @[package.scala 93:22:@55492.4]
  wire  RetimeWrapper_289_reset; // @[package.scala 93:22:@55492.4]
  wire  RetimeWrapper_289_io_flow; // @[package.scala 93:22:@55492.4]
  wire  RetimeWrapper_289_io_in; // @[package.scala 93:22:@55492.4]
  wire  RetimeWrapper_289_io_out; // @[package.scala 93:22:@55492.4]
  wire  RetimeWrapper_290_clock; // @[package.scala 93:22:@55500.4]
  wire  RetimeWrapper_290_reset; // @[package.scala 93:22:@55500.4]
  wire  RetimeWrapper_290_io_flow; // @[package.scala 93:22:@55500.4]
  wire  RetimeWrapper_290_io_in; // @[package.scala 93:22:@55500.4]
  wire  RetimeWrapper_290_io_out; // @[package.scala 93:22:@55500.4]
  wire  RetimeWrapper_291_clock; // @[package.scala 93:22:@55508.4]
  wire  RetimeWrapper_291_reset; // @[package.scala 93:22:@55508.4]
  wire  RetimeWrapper_291_io_flow; // @[package.scala 93:22:@55508.4]
  wire  RetimeWrapper_291_io_in; // @[package.scala 93:22:@55508.4]
  wire  RetimeWrapper_291_io_out; // @[package.scala 93:22:@55508.4]
  wire  RetimeWrapper_292_clock; // @[package.scala 93:22:@55516.4]
  wire  RetimeWrapper_292_reset; // @[package.scala 93:22:@55516.4]
  wire  RetimeWrapper_292_io_flow; // @[package.scala 93:22:@55516.4]
  wire  RetimeWrapper_292_io_in; // @[package.scala 93:22:@55516.4]
  wire  RetimeWrapper_292_io_out; // @[package.scala 93:22:@55516.4]
  wire  RetimeWrapper_293_clock; // @[package.scala 93:22:@55524.4]
  wire  RetimeWrapper_293_reset; // @[package.scala 93:22:@55524.4]
  wire  RetimeWrapper_293_io_flow; // @[package.scala 93:22:@55524.4]
  wire  RetimeWrapper_293_io_in; // @[package.scala 93:22:@55524.4]
  wire  RetimeWrapper_293_io_out; // @[package.scala 93:22:@55524.4]
  wire  RetimeWrapper_294_clock; // @[package.scala 93:22:@55532.4]
  wire  RetimeWrapper_294_reset; // @[package.scala 93:22:@55532.4]
  wire  RetimeWrapper_294_io_flow; // @[package.scala 93:22:@55532.4]
  wire  RetimeWrapper_294_io_in; // @[package.scala 93:22:@55532.4]
  wire  RetimeWrapper_294_io_out; // @[package.scala 93:22:@55532.4]
  wire  RetimeWrapper_295_clock; // @[package.scala 93:22:@55540.4]
  wire  RetimeWrapper_295_reset; // @[package.scala 93:22:@55540.4]
  wire  RetimeWrapper_295_io_flow; // @[package.scala 93:22:@55540.4]
  wire  RetimeWrapper_295_io_in; // @[package.scala 93:22:@55540.4]
  wire  RetimeWrapper_295_io_out; // @[package.scala 93:22:@55540.4]
  wire  RetimeWrapper_296_clock; // @[package.scala 93:22:@55548.4]
  wire  RetimeWrapper_296_reset; // @[package.scala 93:22:@55548.4]
  wire  RetimeWrapper_296_io_flow; // @[package.scala 93:22:@55548.4]
  wire  RetimeWrapper_296_io_in; // @[package.scala 93:22:@55548.4]
  wire  RetimeWrapper_296_io_out; // @[package.scala 93:22:@55548.4]
  wire  RetimeWrapper_297_clock; // @[package.scala 93:22:@55556.4]
  wire  RetimeWrapper_297_reset; // @[package.scala 93:22:@55556.4]
  wire  RetimeWrapper_297_io_flow; // @[package.scala 93:22:@55556.4]
  wire  RetimeWrapper_297_io_in; // @[package.scala 93:22:@55556.4]
  wire  RetimeWrapper_297_io_out; // @[package.scala 93:22:@55556.4]
  wire  RetimeWrapper_298_clock; // @[package.scala 93:22:@55564.4]
  wire  RetimeWrapper_298_reset; // @[package.scala 93:22:@55564.4]
  wire  RetimeWrapper_298_io_flow; // @[package.scala 93:22:@55564.4]
  wire  RetimeWrapper_298_io_in; // @[package.scala 93:22:@55564.4]
  wire  RetimeWrapper_298_io_out; // @[package.scala 93:22:@55564.4]
  wire  RetimeWrapper_299_clock; // @[package.scala 93:22:@55572.4]
  wire  RetimeWrapper_299_reset; // @[package.scala 93:22:@55572.4]
  wire  RetimeWrapper_299_io_flow; // @[package.scala 93:22:@55572.4]
  wire  RetimeWrapper_299_io_in; // @[package.scala 93:22:@55572.4]
  wire  RetimeWrapper_299_io_out; // @[package.scala 93:22:@55572.4]
  wire  RetimeWrapper_300_clock; // @[package.scala 93:22:@55660.4]
  wire  RetimeWrapper_300_reset; // @[package.scala 93:22:@55660.4]
  wire  RetimeWrapper_300_io_flow; // @[package.scala 93:22:@55660.4]
  wire  RetimeWrapper_300_io_in; // @[package.scala 93:22:@55660.4]
  wire  RetimeWrapper_300_io_out; // @[package.scala 93:22:@55660.4]
  wire  RetimeWrapper_301_clock; // @[package.scala 93:22:@55668.4]
  wire  RetimeWrapper_301_reset; // @[package.scala 93:22:@55668.4]
  wire  RetimeWrapper_301_io_flow; // @[package.scala 93:22:@55668.4]
  wire  RetimeWrapper_301_io_in; // @[package.scala 93:22:@55668.4]
  wire  RetimeWrapper_301_io_out; // @[package.scala 93:22:@55668.4]
  wire  RetimeWrapper_302_clock; // @[package.scala 93:22:@55676.4]
  wire  RetimeWrapper_302_reset; // @[package.scala 93:22:@55676.4]
  wire  RetimeWrapper_302_io_flow; // @[package.scala 93:22:@55676.4]
  wire  RetimeWrapper_302_io_in; // @[package.scala 93:22:@55676.4]
  wire  RetimeWrapper_302_io_out; // @[package.scala 93:22:@55676.4]
  wire  RetimeWrapper_303_clock; // @[package.scala 93:22:@55684.4]
  wire  RetimeWrapper_303_reset; // @[package.scala 93:22:@55684.4]
  wire  RetimeWrapper_303_io_flow; // @[package.scala 93:22:@55684.4]
  wire  RetimeWrapper_303_io_in; // @[package.scala 93:22:@55684.4]
  wire  RetimeWrapper_303_io_out; // @[package.scala 93:22:@55684.4]
  wire  RetimeWrapper_304_clock; // @[package.scala 93:22:@55692.4]
  wire  RetimeWrapper_304_reset; // @[package.scala 93:22:@55692.4]
  wire  RetimeWrapper_304_io_flow; // @[package.scala 93:22:@55692.4]
  wire  RetimeWrapper_304_io_in; // @[package.scala 93:22:@55692.4]
  wire  RetimeWrapper_304_io_out; // @[package.scala 93:22:@55692.4]
  wire  RetimeWrapper_305_clock; // @[package.scala 93:22:@55700.4]
  wire  RetimeWrapper_305_reset; // @[package.scala 93:22:@55700.4]
  wire  RetimeWrapper_305_io_flow; // @[package.scala 93:22:@55700.4]
  wire  RetimeWrapper_305_io_in; // @[package.scala 93:22:@55700.4]
  wire  RetimeWrapper_305_io_out; // @[package.scala 93:22:@55700.4]
  wire  RetimeWrapper_306_clock; // @[package.scala 93:22:@55708.4]
  wire  RetimeWrapper_306_reset; // @[package.scala 93:22:@55708.4]
  wire  RetimeWrapper_306_io_flow; // @[package.scala 93:22:@55708.4]
  wire  RetimeWrapper_306_io_in; // @[package.scala 93:22:@55708.4]
  wire  RetimeWrapper_306_io_out; // @[package.scala 93:22:@55708.4]
  wire  RetimeWrapper_307_clock; // @[package.scala 93:22:@55716.4]
  wire  RetimeWrapper_307_reset; // @[package.scala 93:22:@55716.4]
  wire  RetimeWrapper_307_io_flow; // @[package.scala 93:22:@55716.4]
  wire  RetimeWrapper_307_io_in; // @[package.scala 93:22:@55716.4]
  wire  RetimeWrapper_307_io_out; // @[package.scala 93:22:@55716.4]
  wire  RetimeWrapper_308_clock; // @[package.scala 93:22:@55724.4]
  wire  RetimeWrapper_308_reset; // @[package.scala 93:22:@55724.4]
  wire  RetimeWrapper_308_io_flow; // @[package.scala 93:22:@55724.4]
  wire  RetimeWrapper_308_io_in; // @[package.scala 93:22:@55724.4]
  wire  RetimeWrapper_308_io_out; // @[package.scala 93:22:@55724.4]
  wire  RetimeWrapper_309_clock; // @[package.scala 93:22:@55732.4]
  wire  RetimeWrapper_309_reset; // @[package.scala 93:22:@55732.4]
  wire  RetimeWrapper_309_io_flow; // @[package.scala 93:22:@55732.4]
  wire  RetimeWrapper_309_io_in; // @[package.scala 93:22:@55732.4]
  wire  RetimeWrapper_309_io_out; // @[package.scala 93:22:@55732.4]
  wire  RetimeWrapper_310_clock; // @[package.scala 93:22:@55740.4]
  wire  RetimeWrapper_310_reset; // @[package.scala 93:22:@55740.4]
  wire  RetimeWrapper_310_io_flow; // @[package.scala 93:22:@55740.4]
  wire  RetimeWrapper_310_io_in; // @[package.scala 93:22:@55740.4]
  wire  RetimeWrapper_310_io_out; // @[package.scala 93:22:@55740.4]
  wire  RetimeWrapper_311_clock; // @[package.scala 93:22:@55748.4]
  wire  RetimeWrapper_311_reset; // @[package.scala 93:22:@55748.4]
  wire  RetimeWrapper_311_io_flow; // @[package.scala 93:22:@55748.4]
  wire  RetimeWrapper_311_io_in; // @[package.scala 93:22:@55748.4]
  wire  RetimeWrapper_311_io_out; // @[package.scala 93:22:@55748.4]
  wire  RetimeWrapper_312_clock; // @[package.scala 93:22:@55756.4]
  wire  RetimeWrapper_312_reset; // @[package.scala 93:22:@55756.4]
  wire  RetimeWrapper_312_io_flow; // @[package.scala 93:22:@55756.4]
  wire  RetimeWrapper_312_io_in; // @[package.scala 93:22:@55756.4]
  wire  RetimeWrapper_312_io_out; // @[package.scala 93:22:@55756.4]
  wire  RetimeWrapper_313_clock; // @[package.scala 93:22:@55764.4]
  wire  RetimeWrapper_313_reset; // @[package.scala 93:22:@55764.4]
  wire  RetimeWrapper_313_io_flow; // @[package.scala 93:22:@55764.4]
  wire  RetimeWrapper_313_io_in; // @[package.scala 93:22:@55764.4]
  wire  RetimeWrapper_313_io_out; // @[package.scala 93:22:@55764.4]
  wire  RetimeWrapper_314_clock; // @[package.scala 93:22:@55772.4]
  wire  RetimeWrapper_314_reset; // @[package.scala 93:22:@55772.4]
  wire  RetimeWrapper_314_io_flow; // @[package.scala 93:22:@55772.4]
  wire  RetimeWrapper_314_io_in; // @[package.scala 93:22:@55772.4]
  wire  RetimeWrapper_314_io_out; // @[package.scala 93:22:@55772.4]
  wire  RetimeWrapper_315_clock; // @[package.scala 93:22:@55780.4]
  wire  RetimeWrapper_315_reset; // @[package.scala 93:22:@55780.4]
  wire  RetimeWrapper_315_io_flow; // @[package.scala 93:22:@55780.4]
  wire  RetimeWrapper_315_io_in; // @[package.scala 93:22:@55780.4]
  wire  RetimeWrapper_315_io_out; // @[package.scala 93:22:@55780.4]
  wire  RetimeWrapper_316_clock; // @[package.scala 93:22:@55788.4]
  wire  RetimeWrapper_316_reset; // @[package.scala 93:22:@55788.4]
  wire  RetimeWrapper_316_io_flow; // @[package.scala 93:22:@55788.4]
  wire  RetimeWrapper_316_io_in; // @[package.scala 93:22:@55788.4]
  wire  RetimeWrapper_316_io_out; // @[package.scala 93:22:@55788.4]
  wire  RetimeWrapper_317_clock; // @[package.scala 93:22:@55796.4]
  wire  RetimeWrapper_317_reset; // @[package.scala 93:22:@55796.4]
  wire  RetimeWrapper_317_io_flow; // @[package.scala 93:22:@55796.4]
  wire  RetimeWrapper_317_io_in; // @[package.scala 93:22:@55796.4]
  wire  RetimeWrapper_317_io_out; // @[package.scala 93:22:@55796.4]
  wire  RetimeWrapper_318_clock; // @[package.scala 93:22:@55804.4]
  wire  RetimeWrapper_318_reset; // @[package.scala 93:22:@55804.4]
  wire  RetimeWrapper_318_io_flow; // @[package.scala 93:22:@55804.4]
  wire  RetimeWrapper_318_io_in; // @[package.scala 93:22:@55804.4]
  wire  RetimeWrapper_318_io_out; // @[package.scala 93:22:@55804.4]
  wire  RetimeWrapper_319_clock; // @[package.scala 93:22:@55812.4]
  wire  RetimeWrapper_319_reset; // @[package.scala 93:22:@55812.4]
  wire  RetimeWrapper_319_io_flow; // @[package.scala 93:22:@55812.4]
  wire  RetimeWrapper_319_io_in; // @[package.scala 93:22:@55812.4]
  wire  RetimeWrapper_319_io_out; // @[package.scala 93:22:@55812.4]
  wire  RetimeWrapper_320_clock; // @[package.scala 93:22:@55900.4]
  wire  RetimeWrapper_320_reset; // @[package.scala 93:22:@55900.4]
  wire  RetimeWrapper_320_io_flow; // @[package.scala 93:22:@55900.4]
  wire  RetimeWrapper_320_io_in; // @[package.scala 93:22:@55900.4]
  wire  RetimeWrapper_320_io_out; // @[package.scala 93:22:@55900.4]
  wire  RetimeWrapper_321_clock; // @[package.scala 93:22:@55908.4]
  wire  RetimeWrapper_321_reset; // @[package.scala 93:22:@55908.4]
  wire  RetimeWrapper_321_io_flow; // @[package.scala 93:22:@55908.4]
  wire  RetimeWrapper_321_io_in; // @[package.scala 93:22:@55908.4]
  wire  RetimeWrapper_321_io_out; // @[package.scala 93:22:@55908.4]
  wire  RetimeWrapper_322_clock; // @[package.scala 93:22:@55916.4]
  wire  RetimeWrapper_322_reset; // @[package.scala 93:22:@55916.4]
  wire  RetimeWrapper_322_io_flow; // @[package.scala 93:22:@55916.4]
  wire  RetimeWrapper_322_io_in; // @[package.scala 93:22:@55916.4]
  wire  RetimeWrapper_322_io_out; // @[package.scala 93:22:@55916.4]
  wire  RetimeWrapper_323_clock; // @[package.scala 93:22:@55924.4]
  wire  RetimeWrapper_323_reset; // @[package.scala 93:22:@55924.4]
  wire  RetimeWrapper_323_io_flow; // @[package.scala 93:22:@55924.4]
  wire  RetimeWrapper_323_io_in; // @[package.scala 93:22:@55924.4]
  wire  RetimeWrapper_323_io_out; // @[package.scala 93:22:@55924.4]
  wire  RetimeWrapper_324_clock; // @[package.scala 93:22:@55932.4]
  wire  RetimeWrapper_324_reset; // @[package.scala 93:22:@55932.4]
  wire  RetimeWrapper_324_io_flow; // @[package.scala 93:22:@55932.4]
  wire  RetimeWrapper_324_io_in; // @[package.scala 93:22:@55932.4]
  wire  RetimeWrapper_324_io_out; // @[package.scala 93:22:@55932.4]
  wire  RetimeWrapper_325_clock; // @[package.scala 93:22:@55940.4]
  wire  RetimeWrapper_325_reset; // @[package.scala 93:22:@55940.4]
  wire  RetimeWrapper_325_io_flow; // @[package.scala 93:22:@55940.4]
  wire  RetimeWrapper_325_io_in; // @[package.scala 93:22:@55940.4]
  wire  RetimeWrapper_325_io_out; // @[package.scala 93:22:@55940.4]
  wire  RetimeWrapper_326_clock; // @[package.scala 93:22:@55948.4]
  wire  RetimeWrapper_326_reset; // @[package.scala 93:22:@55948.4]
  wire  RetimeWrapper_326_io_flow; // @[package.scala 93:22:@55948.4]
  wire  RetimeWrapper_326_io_in; // @[package.scala 93:22:@55948.4]
  wire  RetimeWrapper_326_io_out; // @[package.scala 93:22:@55948.4]
  wire  RetimeWrapper_327_clock; // @[package.scala 93:22:@55956.4]
  wire  RetimeWrapper_327_reset; // @[package.scala 93:22:@55956.4]
  wire  RetimeWrapper_327_io_flow; // @[package.scala 93:22:@55956.4]
  wire  RetimeWrapper_327_io_in; // @[package.scala 93:22:@55956.4]
  wire  RetimeWrapper_327_io_out; // @[package.scala 93:22:@55956.4]
  wire  RetimeWrapper_328_clock; // @[package.scala 93:22:@55964.4]
  wire  RetimeWrapper_328_reset; // @[package.scala 93:22:@55964.4]
  wire  RetimeWrapper_328_io_flow; // @[package.scala 93:22:@55964.4]
  wire  RetimeWrapper_328_io_in; // @[package.scala 93:22:@55964.4]
  wire  RetimeWrapper_328_io_out; // @[package.scala 93:22:@55964.4]
  wire  RetimeWrapper_329_clock; // @[package.scala 93:22:@55972.4]
  wire  RetimeWrapper_329_reset; // @[package.scala 93:22:@55972.4]
  wire  RetimeWrapper_329_io_flow; // @[package.scala 93:22:@55972.4]
  wire  RetimeWrapper_329_io_in; // @[package.scala 93:22:@55972.4]
  wire  RetimeWrapper_329_io_out; // @[package.scala 93:22:@55972.4]
  wire  RetimeWrapper_330_clock; // @[package.scala 93:22:@55980.4]
  wire  RetimeWrapper_330_reset; // @[package.scala 93:22:@55980.4]
  wire  RetimeWrapper_330_io_flow; // @[package.scala 93:22:@55980.4]
  wire  RetimeWrapper_330_io_in; // @[package.scala 93:22:@55980.4]
  wire  RetimeWrapper_330_io_out; // @[package.scala 93:22:@55980.4]
  wire  RetimeWrapper_331_clock; // @[package.scala 93:22:@55988.4]
  wire  RetimeWrapper_331_reset; // @[package.scala 93:22:@55988.4]
  wire  RetimeWrapper_331_io_flow; // @[package.scala 93:22:@55988.4]
  wire  RetimeWrapper_331_io_in; // @[package.scala 93:22:@55988.4]
  wire  RetimeWrapper_331_io_out; // @[package.scala 93:22:@55988.4]
  wire  RetimeWrapper_332_clock; // @[package.scala 93:22:@55996.4]
  wire  RetimeWrapper_332_reset; // @[package.scala 93:22:@55996.4]
  wire  RetimeWrapper_332_io_flow; // @[package.scala 93:22:@55996.4]
  wire  RetimeWrapper_332_io_in; // @[package.scala 93:22:@55996.4]
  wire  RetimeWrapper_332_io_out; // @[package.scala 93:22:@55996.4]
  wire  RetimeWrapper_333_clock; // @[package.scala 93:22:@56004.4]
  wire  RetimeWrapper_333_reset; // @[package.scala 93:22:@56004.4]
  wire  RetimeWrapper_333_io_flow; // @[package.scala 93:22:@56004.4]
  wire  RetimeWrapper_333_io_in; // @[package.scala 93:22:@56004.4]
  wire  RetimeWrapper_333_io_out; // @[package.scala 93:22:@56004.4]
  wire  RetimeWrapper_334_clock; // @[package.scala 93:22:@56012.4]
  wire  RetimeWrapper_334_reset; // @[package.scala 93:22:@56012.4]
  wire  RetimeWrapper_334_io_flow; // @[package.scala 93:22:@56012.4]
  wire  RetimeWrapper_334_io_in; // @[package.scala 93:22:@56012.4]
  wire  RetimeWrapper_334_io_out; // @[package.scala 93:22:@56012.4]
  wire  RetimeWrapper_335_clock; // @[package.scala 93:22:@56020.4]
  wire  RetimeWrapper_335_reset; // @[package.scala 93:22:@56020.4]
  wire  RetimeWrapper_335_io_flow; // @[package.scala 93:22:@56020.4]
  wire  RetimeWrapper_335_io_in; // @[package.scala 93:22:@56020.4]
  wire  RetimeWrapper_335_io_out; // @[package.scala 93:22:@56020.4]
  wire  RetimeWrapper_336_clock; // @[package.scala 93:22:@56028.4]
  wire  RetimeWrapper_336_reset; // @[package.scala 93:22:@56028.4]
  wire  RetimeWrapper_336_io_flow; // @[package.scala 93:22:@56028.4]
  wire  RetimeWrapper_336_io_in; // @[package.scala 93:22:@56028.4]
  wire  RetimeWrapper_336_io_out; // @[package.scala 93:22:@56028.4]
  wire  RetimeWrapper_337_clock; // @[package.scala 93:22:@56036.4]
  wire  RetimeWrapper_337_reset; // @[package.scala 93:22:@56036.4]
  wire  RetimeWrapper_337_io_flow; // @[package.scala 93:22:@56036.4]
  wire  RetimeWrapper_337_io_in; // @[package.scala 93:22:@56036.4]
  wire  RetimeWrapper_337_io_out; // @[package.scala 93:22:@56036.4]
  wire  RetimeWrapper_338_clock; // @[package.scala 93:22:@56044.4]
  wire  RetimeWrapper_338_reset; // @[package.scala 93:22:@56044.4]
  wire  RetimeWrapper_338_io_flow; // @[package.scala 93:22:@56044.4]
  wire  RetimeWrapper_338_io_in; // @[package.scala 93:22:@56044.4]
  wire  RetimeWrapper_338_io_out; // @[package.scala 93:22:@56044.4]
  wire  RetimeWrapper_339_clock; // @[package.scala 93:22:@56052.4]
  wire  RetimeWrapper_339_reset; // @[package.scala 93:22:@56052.4]
  wire  RetimeWrapper_339_io_flow; // @[package.scala 93:22:@56052.4]
  wire  RetimeWrapper_339_io_in; // @[package.scala 93:22:@56052.4]
  wire  RetimeWrapper_339_io_out; // @[package.scala 93:22:@56052.4]
  wire  RetimeWrapper_340_clock; // @[package.scala 93:22:@56140.4]
  wire  RetimeWrapper_340_reset; // @[package.scala 93:22:@56140.4]
  wire  RetimeWrapper_340_io_flow; // @[package.scala 93:22:@56140.4]
  wire  RetimeWrapper_340_io_in; // @[package.scala 93:22:@56140.4]
  wire  RetimeWrapper_340_io_out; // @[package.scala 93:22:@56140.4]
  wire  RetimeWrapper_341_clock; // @[package.scala 93:22:@56148.4]
  wire  RetimeWrapper_341_reset; // @[package.scala 93:22:@56148.4]
  wire  RetimeWrapper_341_io_flow; // @[package.scala 93:22:@56148.4]
  wire  RetimeWrapper_341_io_in; // @[package.scala 93:22:@56148.4]
  wire  RetimeWrapper_341_io_out; // @[package.scala 93:22:@56148.4]
  wire  RetimeWrapper_342_clock; // @[package.scala 93:22:@56156.4]
  wire  RetimeWrapper_342_reset; // @[package.scala 93:22:@56156.4]
  wire  RetimeWrapper_342_io_flow; // @[package.scala 93:22:@56156.4]
  wire  RetimeWrapper_342_io_in; // @[package.scala 93:22:@56156.4]
  wire  RetimeWrapper_342_io_out; // @[package.scala 93:22:@56156.4]
  wire  RetimeWrapper_343_clock; // @[package.scala 93:22:@56164.4]
  wire  RetimeWrapper_343_reset; // @[package.scala 93:22:@56164.4]
  wire  RetimeWrapper_343_io_flow; // @[package.scala 93:22:@56164.4]
  wire  RetimeWrapper_343_io_in; // @[package.scala 93:22:@56164.4]
  wire  RetimeWrapper_343_io_out; // @[package.scala 93:22:@56164.4]
  wire  RetimeWrapper_344_clock; // @[package.scala 93:22:@56172.4]
  wire  RetimeWrapper_344_reset; // @[package.scala 93:22:@56172.4]
  wire  RetimeWrapper_344_io_flow; // @[package.scala 93:22:@56172.4]
  wire  RetimeWrapper_344_io_in; // @[package.scala 93:22:@56172.4]
  wire  RetimeWrapper_344_io_out; // @[package.scala 93:22:@56172.4]
  wire  RetimeWrapper_345_clock; // @[package.scala 93:22:@56180.4]
  wire  RetimeWrapper_345_reset; // @[package.scala 93:22:@56180.4]
  wire  RetimeWrapper_345_io_flow; // @[package.scala 93:22:@56180.4]
  wire  RetimeWrapper_345_io_in; // @[package.scala 93:22:@56180.4]
  wire  RetimeWrapper_345_io_out; // @[package.scala 93:22:@56180.4]
  wire  RetimeWrapper_346_clock; // @[package.scala 93:22:@56188.4]
  wire  RetimeWrapper_346_reset; // @[package.scala 93:22:@56188.4]
  wire  RetimeWrapper_346_io_flow; // @[package.scala 93:22:@56188.4]
  wire  RetimeWrapper_346_io_in; // @[package.scala 93:22:@56188.4]
  wire  RetimeWrapper_346_io_out; // @[package.scala 93:22:@56188.4]
  wire  RetimeWrapper_347_clock; // @[package.scala 93:22:@56196.4]
  wire  RetimeWrapper_347_reset; // @[package.scala 93:22:@56196.4]
  wire  RetimeWrapper_347_io_flow; // @[package.scala 93:22:@56196.4]
  wire  RetimeWrapper_347_io_in; // @[package.scala 93:22:@56196.4]
  wire  RetimeWrapper_347_io_out; // @[package.scala 93:22:@56196.4]
  wire  RetimeWrapper_348_clock; // @[package.scala 93:22:@56204.4]
  wire  RetimeWrapper_348_reset; // @[package.scala 93:22:@56204.4]
  wire  RetimeWrapper_348_io_flow; // @[package.scala 93:22:@56204.4]
  wire  RetimeWrapper_348_io_in; // @[package.scala 93:22:@56204.4]
  wire  RetimeWrapper_348_io_out; // @[package.scala 93:22:@56204.4]
  wire  RetimeWrapper_349_clock; // @[package.scala 93:22:@56212.4]
  wire  RetimeWrapper_349_reset; // @[package.scala 93:22:@56212.4]
  wire  RetimeWrapper_349_io_flow; // @[package.scala 93:22:@56212.4]
  wire  RetimeWrapper_349_io_in; // @[package.scala 93:22:@56212.4]
  wire  RetimeWrapper_349_io_out; // @[package.scala 93:22:@56212.4]
  wire  RetimeWrapper_350_clock; // @[package.scala 93:22:@56220.4]
  wire  RetimeWrapper_350_reset; // @[package.scala 93:22:@56220.4]
  wire  RetimeWrapper_350_io_flow; // @[package.scala 93:22:@56220.4]
  wire  RetimeWrapper_350_io_in; // @[package.scala 93:22:@56220.4]
  wire  RetimeWrapper_350_io_out; // @[package.scala 93:22:@56220.4]
  wire  RetimeWrapper_351_clock; // @[package.scala 93:22:@56228.4]
  wire  RetimeWrapper_351_reset; // @[package.scala 93:22:@56228.4]
  wire  RetimeWrapper_351_io_flow; // @[package.scala 93:22:@56228.4]
  wire  RetimeWrapper_351_io_in; // @[package.scala 93:22:@56228.4]
  wire  RetimeWrapper_351_io_out; // @[package.scala 93:22:@56228.4]
  wire  RetimeWrapper_352_clock; // @[package.scala 93:22:@56236.4]
  wire  RetimeWrapper_352_reset; // @[package.scala 93:22:@56236.4]
  wire  RetimeWrapper_352_io_flow; // @[package.scala 93:22:@56236.4]
  wire  RetimeWrapper_352_io_in; // @[package.scala 93:22:@56236.4]
  wire  RetimeWrapper_352_io_out; // @[package.scala 93:22:@56236.4]
  wire  RetimeWrapper_353_clock; // @[package.scala 93:22:@56244.4]
  wire  RetimeWrapper_353_reset; // @[package.scala 93:22:@56244.4]
  wire  RetimeWrapper_353_io_flow; // @[package.scala 93:22:@56244.4]
  wire  RetimeWrapper_353_io_in; // @[package.scala 93:22:@56244.4]
  wire  RetimeWrapper_353_io_out; // @[package.scala 93:22:@56244.4]
  wire  RetimeWrapper_354_clock; // @[package.scala 93:22:@56252.4]
  wire  RetimeWrapper_354_reset; // @[package.scala 93:22:@56252.4]
  wire  RetimeWrapper_354_io_flow; // @[package.scala 93:22:@56252.4]
  wire  RetimeWrapper_354_io_in; // @[package.scala 93:22:@56252.4]
  wire  RetimeWrapper_354_io_out; // @[package.scala 93:22:@56252.4]
  wire  RetimeWrapper_355_clock; // @[package.scala 93:22:@56260.4]
  wire  RetimeWrapper_355_reset; // @[package.scala 93:22:@56260.4]
  wire  RetimeWrapper_355_io_flow; // @[package.scala 93:22:@56260.4]
  wire  RetimeWrapper_355_io_in; // @[package.scala 93:22:@56260.4]
  wire  RetimeWrapper_355_io_out; // @[package.scala 93:22:@56260.4]
  wire  RetimeWrapper_356_clock; // @[package.scala 93:22:@56268.4]
  wire  RetimeWrapper_356_reset; // @[package.scala 93:22:@56268.4]
  wire  RetimeWrapper_356_io_flow; // @[package.scala 93:22:@56268.4]
  wire  RetimeWrapper_356_io_in; // @[package.scala 93:22:@56268.4]
  wire  RetimeWrapper_356_io_out; // @[package.scala 93:22:@56268.4]
  wire  RetimeWrapper_357_clock; // @[package.scala 93:22:@56276.4]
  wire  RetimeWrapper_357_reset; // @[package.scala 93:22:@56276.4]
  wire  RetimeWrapper_357_io_flow; // @[package.scala 93:22:@56276.4]
  wire  RetimeWrapper_357_io_in; // @[package.scala 93:22:@56276.4]
  wire  RetimeWrapper_357_io_out; // @[package.scala 93:22:@56276.4]
  wire  RetimeWrapper_358_clock; // @[package.scala 93:22:@56284.4]
  wire  RetimeWrapper_358_reset; // @[package.scala 93:22:@56284.4]
  wire  RetimeWrapper_358_io_flow; // @[package.scala 93:22:@56284.4]
  wire  RetimeWrapper_358_io_in; // @[package.scala 93:22:@56284.4]
  wire  RetimeWrapper_358_io_out; // @[package.scala 93:22:@56284.4]
  wire  RetimeWrapper_359_clock; // @[package.scala 93:22:@56292.4]
  wire  RetimeWrapper_359_reset; // @[package.scala 93:22:@56292.4]
  wire  RetimeWrapper_359_io_flow; // @[package.scala 93:22:@56292.4]
  wire  RetimeWrapper_359_io_in; // @[package.scala 93:22:@56292.4]
  wire  RetimeWrapper_359_io_out; // @[package.scala 93:22:@56292.4]
  wire  RetimeWrapper_360_clock; // @[package.scala 93:22:@56380.4]
  wire  RetimeWrapper_360_reset; // @[package.scala 93:22:@56380.4]
  wire  RetimeWrapper_360_io_flow; // @[package.scala 93:22:@56380.4]
  wire  RetimeWrapper_360_io_in; // @[package.scala 93:22:@56380.4]
  wire  RetimeWrapper_360_io_out; // @[package.scala 93:22:@56380.4]
  wire  RetimeWrapper_361_clock; // @[package.scala 93:22:@56388.4]
  wire  RetimeWrapper_361_reset; // @[package.scala 93:22:@56388.4]
  wire  RetimeWrapper_361_io_flow; // @[package.scala 93:22:@56388.4]
  wire  RetimeWrapper_361_io_in; // @[package.scala 93:22:@56388.4]
  wire  RetimeWrapper_361_io_out; // @[package.scala 93:22:@56388.4]
  wire  RetimeWrapper_362_clock; // @[package.scala 93:22:@56396.4]
  wire  RetimeWrapper_362_reset; // @[package.scala 93:22:@56396.4]
  wire  RetimeWrapper_362_io_flow; // @[package.scala 93:22:@56396.4]
  wire  RetimeWrapper_362_io_in; // @[package.scala 93:22:@56396.4]
  wire  RetimeWrapper_362_io_out; // @[package.scala 93:22:@56396.4]
  wire  RetimeWrapper_363_clock; // @[package.scala 93:22:@56404.4]
  wire  RetimeWrapper_363_reset; // @[package.scala 93:22:@56404.4]
  wire  RetimeWrapper_363_io_flow; // @[package.scala 93:22:@56404.4]
  wire  RetimeWrapper_363_io_in; // @[package.scala 93:22:@56404.4]
  wire  RetimeWrapper_363_io_out; // @[package.scala 93:22:@56404.4]
  wire  RetimeWrapper_364_clock; // @[package.scala 93:22:@56412.4]
  wire  RetimeWrapper_364_reset; // @[package.scala 93:22:@56412.4]
  wire  RetimeWrapper_364_io_flow; // @[package.scala 93:22:@56412.4]
  wire  RetimeWrapper_364_io_in; // @[package.scala 93:22:@56412.4]
  wire  RetimeWrapper_364_io_out; // @[package.scala 93:22:@56412.4]
  wire  RetimeWrapper_365_clock; // @[package.scala 93:22:@56420.4]
  wire  RetimeWrapper_365_reset; // @[package.scala 93:22:@56420.4]
  wire  RetimeWrapper_365_io_flow; // @[package.scala 93:22:@56420.4]
  wire  RetimeWrapper_365_io_in; // @[package.scala 93:22:@56420.4]
  wire  RetimeWrapper_365_io_out; // @[package.scala 93:22:@56420.4]
  wire  RetimeWrapper_366_clock; // @[package.scala 93:22:@56428.4]
  wire  RetimeWrapper_366_reset; // @[package.scala 93:22:@56428.4]
  wire  RetimeWrapper_366_io_flow; // @[package.scala 93:22:@56428.4]
  wire  RetimeWrapper_366_io_in; // @[package.scala 93:22:@56428.4]
  wire  RetimeWrapper_366_io_out; // @[package.scala 93:22:@56428.4]
  wire  RetimeWrapper_367_clock; // @[package.scala 93:22:@56436.4]
  wire  RetimeWrapper_367_reset; // @[package.scala 93:22:@56436.4]
  wire  RetimeWrapper_367_io_flow; // @[package.scala 93:22:@56436.4]
  wire  RetimeWrapper_367_io_in; // @[package.scala 93:22:@56436.4]
  wire  RetimeWrapper_367_io_out; // @[package.scala 93:22:@56436.4]
  wire  RetimeWrapper_368_clock; // @[package.scala 93:22:@56444.4]
  wire  RetimeWrapper_368_reset; // @[package.scala 93:22:@56444.4]
  wire  RetimeWrapper_368_io_flow; // @[package.scala 93:22:@56444.4]
  wire  RetimeWrapper_368_io_in; // @[package.scala 93:22:@56444.4]
  wire  RetimeWrapper_368_io_out; // @[package.scala 93:22:@56444.4]
  wire  RetimeWrapper_369_clock; // @[package.scala 93:22:@56452.4]
  wire  RetimeWrapper_369_reset; // @[package.scala 93:22:@56452.4]
  wire  RetimeWrapper_369_io_flow; // @[package.scala 93:22:@56452.4]
  wire  RetimeWrapper_369_io_in; // @[package.scala 93:22:@56452.4]
  wire  RetimeWrapper_369_io_out; // @[package.scala 93:22:@56452.4]
  wire  RetimeWrapper_370_clock; // @[package.scala 93:22:@56460.4]
  wire  RetimeWrapper_370_reset; // @[package.scala 93:22:@56460.4]
  wire  RetimeWrapper_370_io_flow; // @[package.scala 93:22:@56460.4]
  wire  RetimeWrapper_370_io_in; // @[package.scala 93:22:@56460.4]
  wire  RetimeWrapper_370_io_out; // @[package.scala 93:22:@56460.4]
  wire  RetimeWrapper_371_clock; // @[package.scala 93:22:@56468.4]
  wire  RetimeWrapper_371_reset; // @[package.scala 93:22:@56468.4]
  wire  RetimeWrapper_371_io_flow; // @[package.scala 93:22:@56468.4]
  wire  RetimeWrapper_371_io_in; // @[package.scala 93:22:@56468.4]
  wire  RetimeWrapper_371_io_out; // @[package.scala 93:22:@56468.4]
  wire  RetimeWrapper_372_clock; // @[package.scala 93:22:@56476.4]
  wire  RetimeWrapper_372_reset; // @[package.scala 93:22:@56476.4]
  wire  RetimeWrapper_372_io_flow; // @[package.scala 93:22:@56476.4]
  wire  RetimeWrapper_372_io_in; // @[package.scala 93:22:@56476.4]
  wire  RetimeWrapper_372_io_out; // @[package.scala 93:22:@56476.4]
  wire  RetimeWrapper_373_clock; // @[package.scala 93:22:@56484.4]
  wire  RetimeWrapper_373_reset; // @[package.scala 93:22:@56484.4]
  wire  RetimeWrapper_373_io_flow; // @[package.scala 93:22:@56484.4]
  wire  RetimeWrapper_373_io_in; // @[package.scala 93:22:@56484.4]
  wire  RetimeWrapper_373_io_out; // @[package.scala 93:22:@56484.4]
  wire  RetimeWrapper_374_clock; // @[package.scala 93:22:@56492.4]
  wire  RetimeWrapper_374_reset; // @[package.scala 93:22:@56492.4]
  wire  RetimeWrapper_374_io_flow; // @[package.scala 93:22:@56492.4]
  wire  RetimeWrapper_374_io_in; // @[package.scala 93:22:@56492.4]
  wire  RetimeWrapper_374_io_out; // @[package.scala 93:22:@56492.4]
  wire  RetimeWrapper_375_clock; // @[package.scala 93:22:@56500.4]
  wire  RetimeWrapper_375_reset; // @[package.scala 93:22:@56500.4]
  wire  RetimeWrapper_375_io_flow; // @[package.scala 93:22:@56500.4]
  wire  RetimeWrapper_375_io_in; // @[package.scala 93:22:@56500.4]
  wire  RetimeWrapper_375_io_out; // @[package.scala 93:22:@56500.4]
  wire  RetimeWrapper_376_clock; // @[package.scala 93:22:@56508.4]
  wire  RetimeWrapper_376_reset; // @[package.scala 93:22:@56508.4]
  wire  RetimeWrapper_376_io_flow; // @[package.scala 93:22:@56508.4]
  wire  RetimeWrapper_376_io_in; // @[package.scala 93:22:@56508.4]
  wire  RetimeWrapper_376_io_out; // @[package.scala 93:22:@56508.4]
  wire  RetimeWrapper_377_clock; // @[package.scala 93:22:@56516.4]
  wire  RetimeWrapper_377_reset; // @[package.scala 93:22:@56516.4]
  wire  RetimeWrapper_377_io_flow; // @[package.scala 93:22:@56516.4]
  wire  RetimeWrapper_377_io_in; // @[package.scala 93:22:@56516.4]
  wire  RetimeWrapper_377_io_out; // @[package.scala 93:22:@56516.4]
  wire  RetimeWrapper_378_clock; // @[package.scala 93:22:@56524.4]
  wire  RetimeWrapper_378_reset; // @[package.scala 93:22:@56524.4]
  wire  RetimeWrapper_378_io_flow; // @[package.scala 93:22:@56524.4]
  wire  RetimeWrapper_378_io_in; // @[package.scala 93:22:@56524.4]
  wire  RetimeWrapper_378_io_out; // @[package.scala 93:22:@56524.4]
  wire  RetimeWrapper_379_clock; // @[package.scala 93:22:@56532.4]
  wire  RetimeWrapper_379_reset; // @[package.scala 93:22:@56532.4]
  wire  RetimeWrapper_379_io_flow; // @[package.scala 93:22:@56532.4]
  wire  RetimeWrapper_379_io_in; // @[package.scala 93:22:@56532.4]
  wire  RetimeWrapper_379_io_out; // @[package.scala 93:22:@56532.4]
  wire  RetimeWrapper_380_clock; // @[package.scala 93:22:@56620.4]
  wire  RetimeWrapper_380_reset; // @[package.scala 93:22:@56620.4]
  wire  RetimeWrapper_380_io_flow; // @[package.scala 93:22:@56620.4]
  wire  RetimeWrapper_380_io_in; // @[package.scala 93:22:@56620.4]
  wire  RetimeWrapper_380_io_out; // @[package.scala 93:22:@56620.4]
  wire  RetimeWrapper_381_clock; // @[package.scala 93:22:@56628.4]
  wire  RetimeWrapper_381_reset; // @[package.scala 93:22:@56628.4]
  wire  RetimeWrapper_381_io_flow; // @[package.scala 93:22:@56628.4]
  wire  RetimeWrapper_381_io_in; // @[package.scala 93:22:@56628.4]
  wire  RetimeWrapper_381_io_out; // @[package.scala 93:22:@56628.4]
  wire  RetimeWrapper_382_clock; // @[package.scala 93:22:@56636.4]
  wire  RetimeWrapper_382_reset; // @[package.scala 93:22:@56636.4]
  wire  RetimeWrapper_382_io_flow; // @[package.scala 93:22:@56636.4]
  wire  RetimeWrapper_382_io_in; // @[package.scala 93:22:@56636.4]
  wire  RetimeWrapper_382_io_out; // @[package.scala 93:22:@56636.4]
  wire  RetimeWrapper_383_clock; // @[package.scala 93:22:@56644.4]
  wire  RetimeWrapper_383_reset; // @[package.scala 93:22:@56644.4]
  wire  RetimeWrapper_383_io_flow; // @[package.scala 93:22:@56644.4]
  wire  RetimeWrapper_383_io_in; // @[package.scala 93:22:@56644.4]
  wire  RetimeWrapper_383_io_out; // @[package.scala 93:22:@56644.4]
  wire  RetimeWrapper_384_clock; // @[package.scala 93:22:@56652.4]
  wire  RetimeWrapper_384_reset; // @[package.scala 93:22:@56652.4]
  wire  RetimeWrapper_384_io_flow; // @[package.scala 93:22:@56652.4]
  wire  RetimeWrapper_384_io_in; // @[package.scala 93:22:@56652.4]
  wire  RetimeWrapper_384_io_out; // @[package.scala 93:22:@56652.4]
  wire  RetimeWrapper_385_clock; // @[package.scala 93:22:@56660.4]
  wire  RetimeWrapper_385_reset; // @[package.scala 93:22:@56660.4]
  wire  RetimeWrapper_385_io_flow; // @[package.scala 93:22:@56660.4]
  wire  RetimeWrapper_385_io_in; // @[package.scala 93:22:@56660.4]
  wire  RetimeWrapper_385_io_out; // @[package.scala 93:22:@56660.4]
  wire  RetimeWrapper_386_clock; // @[package.scala 93:22:@56668.4]
  wire  RetimeWrapper_386_reset; // @[package.scala 93:22:@56668.4]
  wire  RetimeWrapper_386_io_flow; // @[package.scala 93:22:@56668.4]
  wire  RetimeWrapper_386_io_in; // @[package.scala 93:22:@56668.4]
  wire  RetimeWrapper_386_io_out; // @[package.scala 93:22:@56668.4]
  wire  RetimeWrapper_387_clock; // @[package.scala 93:22:@56676.4]
  wire  RetimeWrapper_387_reset; // @[package.scala 93:22:@56676.4]
  wire  RetimeWrapper_387_io_flow; // @[package.scala 93:22:@56676.4]
  wire  RetimeWrapper_387_io_in; // @[package.scala 93:22:@56676.4]
  wire  RetimeWrapper_387_io_out; // @[package.scala 93:22:@56676.4]
  wire  RetimeWrapper_388_clock; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_388_reset; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_388_io_flow; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_388_io_in; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_388_io_out; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_389_clock; // @[package.scala 93:22:@56692.4]
  wire  RetimeWrapper_389_reset; // @[package.scala 93:22:@56692.4]
  wire  RetimeWrapper_389_io_flow; // @[package.scala 93:22:@56692.4]
  wire  RetimeWrapper_389_io_in; // @[package.scala 93:22:@56692.4]
  wire  RetimeWrapper_389_io_out; // @[package.scala 93:22:@56692.4]
  wire  RetimeWrapper_390_clock; // @[package.scala 93:22:@56700.4]
  wire  RetimeWrapper_390_reset; // @[package.scala 93:22:@56700.4]
  wire  RetimeWrapper_390_io_flow; // @[package.scala 93:22:@56700.4]
  wire  RetimeWrapper_390_io_in; // @[package.scala 93:22:@56700.4]
  wire  RetimeWrapper_390_io_out; // @[package.scala 93:22:@56700.4]
  wire  RetimeWrapper_391_clock; // @[package.scala 93:22:@56708.4]
  wire  RetimeWrapper_391_reset; // @[package.scala 93:22:@56708.4]
  wire  RetimeWrapper_391_io_flow; // @[package.scala 93:22:@56708.4]
  wire  RetimeWrapper_391_io_in; // @[package.scala 93:22:@56708.4]
  wire  RetimeWrapper_391_io_out; // @[package.scala 93:22:@56708.4]
  wire  RetimeWrapper_392_clock; // @[package.scala 93:22:@56716.4]
  wire  RetimeWrapper_392_reset; // @[package.scala 93:22:@56716.4]
  wire  RetimeWrapper_392_io_flow; // @[package.scala 93:22:@56716.4]
  wire  RetimeWrapper_392_io_in; // @[package.scala 93:22:@56716.4]
  wire  RetimeWrapper_392_io_out; // @[package.scala 93:22:@56716.4]
  wire  RetimeWrapper_393_clock; // @[package.scala 93:22:@56724.4]
  wire  RetimeWrapper_393_reset; // @[package.scala 93:22:@56724.4]
  wire  RetimeWrapper_393_io_flow; // @[package.scala 93:22:@56724.4]
  wire  RetimeWrapper_393_io_in; // @[package.scala 93:22:@56724.4]
  wire  RetimeWrapper_393_io_out; // @[package.scala 93:22:@56724.4]
  wire  RetimeWrapper_394_clock; // @[package.scala 93:22:@56732.4]
  wire  RetimeWrapper_394_reset; // @[package.scala 93:22:@56732.4]
  wire  RetimeWrapper_394_io_flow; // @[package.scala 93:22:@56732.4]
  wire  RetimeWrapper_394_io_in; // @[package.scala 93:22:@56732.4]
  wire  RetimeWrapper_394_io_out; // @[package.scala 93:22:@56732.4]
  wire  RetimeWrapper_395_clock; // @[package.scala 93:22:@56740.4]
  wire  RetimeWrapper_395_reset; // @[package.scala 93:22:@56740.4]
  wire  RetimeWrapper_395_io_flow; // @[package.scala 93:22:@56740.4]
  wire  RetimeWrapper_395_io_in; // @[package.scala 93:22:@56740.4]
  wire  RetimeWrapper_395_io_out; // @[package.scala 93:22:@56740.4]
  wire  RetimeWrapper_396_clock; // @[package.scala 93:22:@56748.4]
  wire  RetimeWrapper_396_reset; // @[package.scala 93:22:@56748.4]
  wire  RetimeWrapper_396_io_flow; // @[package.scala 93:22:@56748.4]
  wire  RetimeWrapper_396_io_in; // @[package.scala 93:22:@56748.4]
  wire  RetimeWrapper_396_io_out; // @[package.scala 93:22:@56748.4]
  wire  RetimeWrapper_397_clock; // @[package.scala 93:22:@56756.4]
  wire  RetimeWrapper_397_reset; // @[package.scala 93:22:@56756.4]
  wire  RetimeWrapper_397_io_flow; // @[package.scala 93:22:@56756.4]
  wire  RetimeWrapper_397_io_in; // @[package.scala 93:22:@56756.4]
  wire  RetimeWrapper_397_io_out; // @[package.scala 93:22:@56756.4]
  wire  RetimeWrapper_398_clock; // @[package.scala 93:22:@56764.4]
  wire  RetimeWrapper_398_reset; // @[package.scala 93:22:@56764.4]
  wire  RetimeWrapper_398_io_flow; // @[package.scala 93:22:@56764.4]
  wire  RetimeWrapper_398_io_in; // @[package.scala 93:22:@56764.4]
  wire  RetimeWrapper_398_io_out; // @[package.scala 93:22:@56764.4]
  wire  RetimeWrapper_399_clock; // @[package.scala 93:22:@56772.4]
  wire  RetimeWrapper_399_reset; // @[package.scala 93:22:@56772.4]
  wire  RetimeWrapper_399_io_flow; // @[package.scala 93:22:@56772.4]
  wire  RetimeWrapper_399_io_in; // @[package.scala 93:22:@56772.4]
  wire  RetimeWrapper_399_io_out; // @[package.scala 93:22:@56772.4]
  wire  RetimeWrapper_400_clock; // @[package.scala 93:22:@56860.4]
  wire  RetimeWrapper_400_reset; // @[package.scala 93:22:@56860.4]
  wire  RetimeWrapper_400_io_flow; // @[package.scala 93:22:@56860.4]
  wire  RetimeWrapper_400_io_in; // @[package.scala 93:22:@56860.4]
  wire  RetimeWrapper_400_io_out; // @[package.scala 93:22:@56860.4]
  wire  RetimeWrapper_401_clock; // @[package.scala 93:22:@56868.4]
  wire  RetimeWrapper_401_reset; // @[package.scala 93:22:@56868.4]
  wire  RetimeWrapper_401_io_flow; // @[package.scala 93:22:@56868.4]
  wire  RetimeWrapper_401_io_in; // @[package.scala 93:22:@56868.4]
  wire  RetimeWrapper_401_io_out; // @[package.scala 93:22:@56868.4]
  wire  RetimeWrapper_402_clock; // @[package.scala 93:22:@56876.4]
  wire  RetimeWrapper_402_reset; // @[package.scala 93:22:@56876.4]
  wire  RetimeWrapper_402_io_flow; // @[package.scala 93:22:@56876.4]
  wire  RetimeWrapper_402_io_in; // @[package.scala 93:22:@56876.4]
  wire  RetimeWrapper_402_io_out; // @[package.scala 93:22:@56876.4]
  wire  RetimeWrapper_403_clock; // @[package.scala 93:22:@56884.4]
  wire  RetimeWrapper_403_reset; // @[package.scala 93:22:@56884.4]
  wire  RetimeWrapper_403_io_flow; // @[package.scala 93:22:@56884.4]
  wire  RetimeWrapper_403_io_in; // @[package.scala 93:22:@56884.4]
  wire  RetimeWrapper_403_io_out; // @[package.scala 93:22:@56884.4]
  wire  RetimeWrapper_404_clock; // @[package.scala 93:22:@56892.4]
  wire  RetimeWrapper_404_reset; // @[package.scala 93:22:@56892.4]
  wire  RetimeWrapper_404_io_flow; // @[package.scala 93:22:@56892.4]
  wire  RetimeWrapper_404_io_in; // @[package.scala 93:22:@56892.4]
  wire  RetimeWrapper_404_io_out; // @[package.scala 93:22:@56892.4]
  wire  RetimeWrapper_405_clock; // @[package.scala 93:22:@56900.4]
  wire  RetimeWrapper_405_reset; // @[package.scala 93:22:@56900.4]
  wire  RetimeWrapper_405_io_flow; // @[package.scala 93:22:@56900.4]
  wire  RetimeWrapper_405_io_in; // @[package.scala 93:22:@56900.4]
  wire  RetimeWrapper_405_io_out; // @[package.scala 93:22:@56900.4]
  wire  RetimeWrapper_406_clock; // @[package.scala 93:22:@56908.4]
  wire  RetimeWrapper_406_reset; // @[package.scala 93:22:@56908.4]
  wire  RetimeWrapper_406_io_flow; // @[package.scala 93:22:@56908.4]
  wire  RetimeWrapper_406_io_in; // @[package.scala 93:22:@56908.4]
  wire  RetimeWrapper_406_io_out; // @[package.scala 93:22:@56908.4]
  wire  RetimeWrapper_407_clock; // @[package.scala 93:22:@56916.4]
  wire  RetimeWrapper_407_reset; // @[package.scala 93:22:@56916.4]
  wire  RetimeWrapper_407_io_flow; // @[package.scala 93:22:@56916.4]
  wire  RetimeWrapper_407_io_in; // @[package.scala 93:22:@56916.4]
  wire  RetimeWrapper_407_io_out; // @[package.scala 93:22:@56916.4]
  wire  RetimeWrapper_408_clock; // @[package.scala 93:22:@56924.4]
  wire  RetimeWrapper_408_reset; // @[package.scala 93:22:@56924.4]
  wire  RetimeWrapper_408_io_flow; // @[package.scala 93:22:@56924.4]
  wire  RetimeWrapper_408_io_in; // @[package.scala 93:22:@56924.4]
  wire  RetimeWrapper_408_io_out; // @[package.scala 93:22:@56924.4]
  wire  RetimeWrapper_409_clock; // @[package.scala 93:22:@56932.4]
  wire  RetimeWrapper_409_reset; // @[package.scala 93:22:@56932.4]
  wire  RetimeWrapper_409_io_flow; // @[package.scala 93:22:@56932.4]
  wire  RetimeWrapper_409_io_in; // @[package.scala 93:22:@56932.4]
  wire  RetimeWrapper_409_io_out; // @[package.scala 93:22:@56932.4]
  wire  RetimeWrapper_410_clock; // @[package.scala 93:22:@56940.4]
  wire  RetimeWrapper_410_reset; // @[package.scala 93:22:@56940.4]
  wire  RetimeWrapper_410_io_flow; // @[package.scala 93:22:@56940.4]
  wire  RetimeWrapper_410_io_in; // @[package.scala 93:22:@56940.4]
  wire  RetimeWrapper_410_io_out; // @[package.scala 93:22:@56940.4]
  wire  RetimeWrapper_411_clock; // @[package.scala 93:22:@56948.4]
  wire  RetimeWrapper_411_reset; // @[package.scala 93:22:@56948.4]
  wire  RetimeWrapper_411_io_flow; // @[package.scala 93:22:@56948.4]
  wire  RetimeWrapper_411_io_in; // @[package.scala 93:22:@56948.4]
  wire  RetimeWrapper_411_io_out; // @[package.scala 93:22:@56948.4]
  wire  RetimeWrapper_412_clock; // @[package.scala 93:22:@56956.4]
  wire  RetimeWrapper_412_reset; // @[package.scala 93:22:@56956.4]
  wire  RetimeWrapper_412_io_flow; // @[package.scala 93:22:@56956.4]
  wire  RetimeWrapper_412_io_in; // @[package.scala 93:22:@56956.4]
  wire  RetimeWrapper_412_io_out; // @[package.scala 93:22:@56956.4]
  wire  RetimeWrapper_413_clock; // @[package.scala 93:22:@56964.4]
  wire  RetimeWrapper_413_reset; // @[package.scala 93:22:@56964.4]
  wire  RetimeWrapper_413_io_flow; // @[package.scala 93:22:@56964.4]
  wire  RetimeWrapper_413_io_in; // @[package.scala 93:22:@56964.4]
  wire  RetimeWrapper_413_io_out; // @[package.scala 93:22:@56964.4]
  wire  RetimeWrapper_414_clock; // @[package.scala 93:22:@56972.4]
  wire  RetimeWrapper_414_reset; // @[package.scala 93:22:@56972.4]
  wire  RetimeWrapper_414_io_flow; // @[package.scala 93:22:@56972.4]
  wire  RetimeWrapper_414_io_in; // @[package.scala 93:22:@56972.4]
  wire  RetimeWrapper_414_io_out; // @[package.scala 93:22:@56972.4]
  wire  RetimeWrapper_415_clock; // @[package.scala 93:22:@56980.4]
  wire  RetimeWrapper_415_reset; // @[package.scala 93:22:@56980.4]
  wire  RetimeWrapper_415_io_flow; // @[package.scala 93:22:@56980.4]
  wire  RetimeWrapper_415_io_in; // @[package.scala 93:22:@56980.4]
  wire  RetimeWrapper_415_io_out; // @[package.scala 93:22:@56980.4]
  wire  RetimeWrapper_416_clock; // @[package.scala 93:22:@56988.4]
  wire  RetimeWrapper_416_reset; // @[package.scala 93:22:@56988.4]
  wire  RetimeWrapper_416_io_flow; // @[package.scala 93:22:@56988.4]
  wire  RetimeWrapper_416_io_in; // @[package.scala 93:22:@56988.4]
  wire  RetimeWrapper_416_io_out; // @[package.scala 93:22:@56988.4]
  wire  RetimeWrapper_417_clock; // @[package.scala 93:22:@56996.4]
  wire  RetimeWrapper_417_reset; // @[package.scala 93:22:@56996.4]
  wire  RetimeWrapper_417_io_flow; // @[package.scala 93:22:@56996.4]
  wire  RetimeWrapper_417_io_in; // @[package.scala 93:22:@56996.4]
  wire  RetimeWrapper_417_io_out; // @[package.scala 93:22:@56996.4]
  wire  RetimeWrapper_418_clock; // @[package.scala 93:22:@57004.4]
  wire  RetimeWrapper_418_reset; // @[package.scala 93:22:@57004.4]
  wire  RetimeWrapper_418_io_flow; // @[package.scala 93:22:@57004.4]
  wire  RetimeWrapper_418_io_in; // @[package.scala 93:22:@57004.4]
  wire  RetimeWrapper_418_io_out; // @[package.scala 93:22:@57004.4]
  wire  RetimeWrapper_419_clock; // @[package.scala 93:22:@57012.4]
  wire  RetimeWrapper_419_reset; // @[package.scala 93:22:@57012.4]
  wire  RetimeWrapper_419_io_flow; // @[package.scala 93:22:@57012.4]
  wire  RetimeWrapper_419_io_in; // @[package.scala 93:22:@57012.4]
  wire  RetimeWrapper_419_io_out; // @[package.scala 93:22:@57012.4]
  wire  RetimeWrapper_420_clock; // @[package.scala 93:22:@57100.4]
  wire  RetimeWrapper_420_reset; // @[package.scala 93:22:@57100.4]
  wire  RetimeWrapper_420_io_flow; // @[package.scala 93:22:@57100.4]
  wire  RetimeWrapper_420_io_in; // @[package.scala 93:22:@57100.4]
  wire  RetimeWrapper_420_io_out; // @[package.scala 93:22:@57100.4]
  wire  RetimeWrapper_421_clock; // @[package.scala 93:22:@57108.4]
  wire  RetimeWrapper_421_reset; // @[package.scala 93:22:@57108.4]
  wire  RetimeWrapper_421_io_flow; // @[package.scala 93:22:@57108.4]
  wire  RetimeWrapper_421_io_in; // @[package.scala 93:22:@57108.4]
  wire  RetimeWrapper_421_io_out; // @[package.scala 93:22:@57108.4]
  wire  RetimeWrapper_422_clock; // @[package.scala 93:22:@57116.4]
  wire  RetimeWrapper_422_reset; // @[package.scala 93:22:@57116.4]
  wire  RetimeWrapper_422_io_flow; // @[package.scala 93:22:@57116.4]
  wire  RetimeWrapper_422_io_in; // @[package.scala 93:22:@57116.4]
  wire  RetimeWrapper_422_io_out; // @[package.scala 93:22:@57116.4]
  wire  RetimeWrapper_423_clock; // @[package.scala 93:22:@57124.4]
  wire  RetimeWrapper_423_reset; // @[package.scala 93:22:@57124.4]
  wire  RetimeWrapper_423_io_flow; // @[package.scala 93:22:@57124.4]
  wire  RetimeWrapper_423_io_in; // @[package.scala 93:22:@57124.4]
  wire  RetimeWrapper_423_io_out; // @[package.scala 93:22:@57124.4]
  wire  RetimeWrapper_424_clock; // @[package.scala 93:22:@57132.4]
  wire  RetimeWrapper_424_reset; // @[package.scala 93:22:@57132.4]
  wire  RetimeWrapper_424_io_flow; // @[package.scala 93:22:@57132.4]
  wire  RetimeWrapper_424_io_in; // @[package.scala 93:22:@57132.4]
  wire  RetimeWrapper_424_io_out; // @[package.scala 93:22:@57132.4]
  wire  RetimeWrapper_425_clock; // @[package.scala 93:22:@57140.4]
  wire  RetimeWrapper_425_reset; // @[package.scala 93:22:@57140.4]
  wire  RetimeWrapper_425_io_flow; // @[package.scala 93:22:@57140.4]
  wire  RetimeWrapper_425_io_in; // @[package.scala 93:22:@57140.4]
  wire  RetimeWrapper_425_io_out; // @[package.scala 93:22:@57140.4]
  wire  RetimeWrapper_426_clock; // @[package.scala 93:22:@57148.4]
  wire  RetimeWrapper_426_reset; // @[package.scala 93:22:@57148.4]
  wire  RetimeWrapper_426_io_flow; // @[package.scala 93:22:@57148.4]
  wire  RetimeWrapper_426_io_in; // @[package.scala 93:22:@57148.4]
  wire  RetimeWrapper_426_io_out; // @[package.scala 93:22:@57148.4]
  wire  RetimeWrapper_427_clock; // @[package.scala 93:22:@57156.4]
  wire  RetimeWrapper_427_reset; // @[package.scala 93:22:@57156.4]
  wire  RetimeWrapper_427_io_flow; // @[package.scala 93:22:@57156.4]
  wire  RetimeWrapper_427_io_in; // @[package.scala 93:22:@57156.4]
  wire  RetimeWrapper_427_io_out; // @[package.scala 93:22:@57156.4]
  wire  RetimeWrapper_428_clock; // @[package.scala 93:22:@57164.4]
  wire  RetimeWrapper_428_reset; // @[package.scala 93:22:@57164.4]
  wire  RetimeWrapper_428_io_flow; // @[package.scala 93:22:@57164.4]
  wire  RetimeWrapper_428_io_in; // @[package.scala 93:22:@57164.4]
  wire  RetimeWrapper_428_io_out; // @[package.scala 93:22:@57164.4]
  wire  RetimeWrapper_429_clock; // @[package.scala 93:22:@57172.4]
  wire  RetimeWrapper_429_reset; // @[package.scala 93:22:@57172.4]
  wire  RetimeWrapper_429_io_flow; // @[package.scala 93:22:@57172.4]
  wire  RetimeWrapper_429_io_in; // @[package.scala 93:22:@57172.4]
  wire  RetimeWrapper_429_io_out; // @[package.scala 93:22:@57172.4]
  wire  RetimeWrapper_430_clock; // @[package.scala 93:22:@57180.4]
  wire  RetimeWrapper_430_reset; // @[package.scala 93:22:@57180.4]
  wire  RetimeWrapper_430_io_flow; // @[package.scala 93:22:@57180.4]
  wire  RetimeWrapper_430_io_in; // @[package.scala 93:22:@57180.4]
  wire  RetimeWrapper_430_io_out; // @[package.scala 93:22:@57180.4]
  wire  RetimeWrapper_431_clock; // @[package.scala 93:22:@57188.4]
  wire  RetimeWrapper_431_reset; // @[package.scala 93:22:@57188.4]
  wire  RetimeWrapper_431_io_flow; // @[package.scala 93:22:@57188.4]
  wire  RetimeWrapper_431_io_in; // @[package.scala 93:22:@57188.4]
  wire  RetimeWrapper_431_io_out; // @[package.scala 93:22:@57188.4]
  wire  RetimeWrapper_432_clock; // @[package.scala 93:22:@57196.4]
  wire  RetimeWrapper_432_reset; // @[package.scala 93:22:@57196.4]
  wire  RetimeWrapper_432_io_flow; // @[package.scala 93:22:@57196.4]
  wire  RetimeWrapper_432_io_in; // @[package.scala 93:22:@57196.4]
  wire  RetimeWrapper_432_io_out; // @[package.scala 93:22:@57196.4]
  wire  RetimeWrapper_433_clock; // @[package.scala 93:22:@57204.4]
  wire  RetimeWrapper_433_reset; // @[package.scala 93:22:@57204.4]
  wire  RetimeWrapper_433_io_flow; // @[package.scala 93:22:@57204.4]
  wire  RetimeWrapper_433_io_in; // @[package.scala 93:22:@57204.4]
  wire  RetimeWrapper_433_io_out; // @[package.scala 93:22:@57204.4]
  wire  RetimeWrapper_434_clock; // @[package.scala 93:22:@57212.4]
  wire  RetimeWrapper_434_reset; // @[package.scala 93:22:@57212.4]
  wire  RetimeWrapper_434_io_flow; // @[package.scala 93:22:@57212.4]
  wire  RetimeWrapper_434_io_in; // @[package.scala 93:22:@57212.4]
  wire  RetimeWrapper_434_io_out; // @[package.scala 93:22:@57212.4]
  wire  RetimeWrapper_435_clock; // @[package.scala 93:22:@57220.4]
  wire  RetimeWrapper_435_reset; // @[package.scala 93:22:@57220.4]
  wire  RetimeWrapper_435_io_flow; // @[package.scala 93:22:@57220.4]
  wire  RetimeWrapper_435_io_in; // @[package.scala 93:22:@57220.4]
  wire  RetimeWrapper_435_io_out; // @[package.scala 93:22:@57220.4]
  wire  RetimeWrapper_436_clock; // @[package.scala 93:22:@57228.4]
  wire  RetimeWrapper_436_reset; // @[package.scala 93:22:@57228.4]
  wire  RetimeWrapper_436_io_flow; // @[package.scala 93:22:@57228.4]
  wire  RetimeWrapper_436_io_in; // @[package.scala 93:22:@57228.4]
  wire  RetimeWrapper_436_io_out; // @[package.scala 93:22:@57228.4]
  wire  RetimeWrapper_437_clock; // @[package.scala 93:22:@57236.4]
  wire  RetimeWrapper_437_reset; // @[package.scala 93:22:@57236.4]
  wire  RetimeWrapper_437_io_flow; // @[package.scala 93:22:@57236.4]
  wire  RetimeWrapper_437_io_in; // @[package.scala 93:22:@57236.4]
  wire  RetimeWrapper_437_io_out; // @[package.scala 93:22:@57236.4]
  wire  RetimeWrapper_438_clock; // @[package.scala 93:22:@57244.4]
  wire  RetimeWrapper_438_reset; // @[package.scala 93:22:@57244.4]
  wire  RetimeWrapper_438_io_flow; // @[package.scala 93:22:@57244.4]
  wire  RetimeWrapper_438_io_in; // @[package.scala 93:22:@57244.4]
  wire  RetimeWrapper_438_io_out; // @[package.scala 93:22:@57244.4]
  wire  RetimeWrapper_439_clock; // @[package.scala 93:22:@57252.4]
  wire  RetimeWrapper_439_reset; // @[package.scala 93:22:@57252.4]
  wire  RetimeWrapper_439_io_flow; // @[package.scala 93:22:@57252.4]
  wire  RetimeWrapper_439_io_in; // @[package.scala 93:22:@57252.4]
  wire  RetimeWrapper_439_io_out; // @[package.scala 93:22:@57252.4]
  wire  RetimeWrapper_440_clock; // @[package.scala 93:22:@57340.4]
  wire  RetimeWrapper_440_reset; // @[package.scala 93:22:@57340.4]
  wire  RetimeWrapper_440_io_flow; // @[package.scala 93:22:@57340.4]
  wire  RetimeWrapper_440_io_in; // @[package.scala 93:22:@57340.4]
  wire  RetimeWrapper_440_io_out; // @[package.scala 93:22:@57340.4]
  wire  RetimeWrapper_441_clock; // @[package.scala 93:22:@57348.4]
  wire  RetimeWrapper_441_reset; // @[package.scala 93:22:@57348.4]
  wire  RetimeWrapper_441_io_flow; // @[package.scala 93:22:@57348.4]
  wire  RetimeWrapper_441_io_in; // @[package.scala 93:22:@57348.4]
  wire  RetimeWrapper_441_io_out; // @[package.scala 93:22:@57348.4]
  wire  RetimeWrapper_442_clock; // @[package.scala 93:22:@57356.4]
  wire  RetimeWrapper_442_reset; // @[package.scala 93:22:@57356.4]
  wire  RetimeWrapper_442_io_flow; // @[package.scala 93:22:@57356.4]
  wire  RetimeWrapper_442_io_in; // @[package.scala 93:22:@57356.4]
  wire  RetimeWrapper_442_io_out; // @[package.scala 93:22:@57356.4]
  wire  RetimeWrapper_443_clock; // @[package.scala 93:22:@57364.4]
  wire  RetimeWrapper_443_reset; // @[package.scala 93:22:@57364.4]
  wire  RetimeWrapper_443_io_flow; // @[package.scala 93:22:@57364.4]
  wire  RetimeWrapper_443_io_in; // @[package.scala 93:22:@57364.4]
  wire  RetimeWrapper_443_io_out; // @[package.scala 93:22:@57364.4]
  wire  RetimeWrapper_444_clock; // @[package.scala 93:22:@57372.4]
  wire  RetimeWrapper_444_reset; // @[package.scala 93:22:@57372.4]
  wire  RetimeWrapper_444_io_flow; // @[package.scala 93:22:@57372.4]
  wire  RetimeWrapper_444_io_in; // @[package.scala 93:22:@57372.4]
  wire  RetimeWrapper_444_io_out; // @[package.scala 93:22:@57372.4]
  wire  RetimeWrapper_445_clock; // @[package.scala 93:22:@57380.4]
  wire  RetimeWrapper_445_reset; // @[package.scala 93:22:@57380.4]
  wire  RetimeWrapper_445_io_flow; // @[package.scala 93:22:@57380.4]
  wire  RetimeWrapper_445_io_in; // @[package.scala 93:22:@57380.4]
  wire  RetimeWrapper_445_io_out; // @[package.scala 93:22:@57380.4]
  wire  RetimeWrapper_446_clock; // @[package.scala 93:22:@57388.4]
  wire  RetimeWrapper_446_reset; // @[package.scala 93:22:@57388.4]
  wire  RetimeWrapper_446_io_flow; // @[package.scala 93:22:@57388.4]
  wire  RetimeWrapper_446_io_in; // @[package.scala 93:22:@57388.4]
  wire  RetimeWrapper_446_io_out; // @[package.scala 93:22:@57388.4]
  wire  RetimeWrapper_447_clock; // @[package.scala 93:22:@57396.4]
  wire  RetimeWrapper_447_reset; // @[package.scala 93:22:@57396.4]
  wire  RetimeWrapper_447_io_flow; // @[package.scala 93:22:@57396.4]
  wire  RetimeWrapper_447_io_in; // @[package.scala 93:22:@57396.4]
  wire  RetimeWrapper_447_io_out; // @[package.scala 93:22:@57396.4]
  wire  RetimeWrapper_448_clock; // @[package.scala 93:22:@57404.4]
  wire  RetimeWrapper_448_reset; // @[package.scala 93:22:@57404.4]
  wire  RetimeWrapper_448_io_flow; // @[package.scala 93:22:@57404.4]
  wire  RetimeWrapper_448_io_in; // @[package.scala 93:22:@57404.4]
  wire  RetimeWrapper_448_io_out; // @[package.scala 93:22:@57404.4]
  wire  RetimeWrapper_449_clock; // @[package.scala 93:22:@57412.4]
  wire  RetimeWrapper_449_reset; // @[package.scala 93:22:@57412.4]
  wire  RetimeWrapper_449_io_flow; // @[package.scala 93:22:@57412.4]
  wire  RetimeWrapper_449_io_in; // @[package.scala 93:22:@57412.4]
  wire  RetimeWrapper_449_io_out; // @[package.scala 93:22:@57412.4]
  wire  RetimeWrapper_450_clock; // @[package.scala 93:22:@57420.4]
  wire  RetimeWrapper_450_reset; // @[package.scala 93:22:@57420.4]
  wire  RetimeWrapper_450_io_flow; // @[package.scala 93:22:@57420.4]
  wire  RetimeWrapper_450_io_in; // @[package.scala 93:22:@57420.4]
  wire  RetimeWrapper_450_io_out; // @[package.scala 93:22:@57420.4]
  wire  RetimeWrapper_451_clock; // @[package.scala 93:22:@57428.4]
  wire  RetimeWrapper_451_reset; // @[package.scala 93:22:@57428.4]
  wire  RetimeWrapper_451_io_flow; // @[package.scala 93:22:@57428.4]
  wire  RetimeWrapper_451_io_in; // @[package.scala 93:22:@57428.4]
  wire  RetimeWrapper_451_io_out; // @[package.scala 93:22:@57428.4]
  wire  RetimeWrapper_452_clock; // @[package.scala 93:22:@57436.4]
  wire  RetimeWrapper_452_reset; // @[package.scala 93:22:@57436.4]
  wire  RetimeWrapper_452_io_flow; // @[package.scala 93:22:@57436.4]
  wire  RetimeWrapper_452_io_in; // @[package.scala 93:22:@57436.4]
  wire  RetimeWrapper_452_io_out; // @[package.scala 93:22:@57436.4]
  wire  RetimeWrapper_453_clock; // @[package.scala 93:22:@57444.4]
  wire  RetimeWrapper_453_reset; // @[package.scala 93:22:@57444.4]
  wire  RetimeWrapper_453_io_flow; // @[package.scala 93:22:@57444.4]
  wire  RetimeWrapper_453_io_in; // @[package.scala 93:22:@57444.4]
  wire  RetimeWrapper_453_io_out; // @[package.scala 93:22:@57444.4]
  wire  RetimeWrapper_454_clock; // @[package.scala 93:22:@57452.4]
  wire  RetimeWrapper_454_reset; // @[package.scala 93:22:@57452.4]
  wire  RetimeWrapper_454_io_flow; // @[package.scala 93:22:@57452.4]
  wire  RetimeWrapper_454_io_in; // @[package.scala 93:22:@57452.4]
  wire  RetimeWrapper_454_io_out; // @[package.scala 93:22:@57452.4]
  wire  RetimeWrapper_455_clock; // @[package.scala 93:22:@57460.4]
  wire  RetimeWrapper_455_reset; // @[package.scala 93:22:@57460.4]
  wire  RetimeWrapper_455_io_flow; // @[package.scala 93:22:@57460.4]
  wire  RetimeWrapper_455_io_in; // @[package.scala 93:22:@57460.4]
  wire  RetimeWrapper_455_io_out; // @[package.scala 93:22:@57460.4]
  wire  RetimeWrapper_456_clock; // @[package.scala 93:22:@57468.4]
  wire  RetimeWrapper_456_reset; // @[package.scala 93:22:@57468.4]
  wire  RetimeWrapper_456_io_flow; // @[package.scala 93:22:@57468.4]
  wire  RetimeWrapper_456_io_in; // @[package.scala 93:22:@57468.4]
  wire  RetimeWrapper_456_io_out; // @[package.scala 93:22:@57468.4]
  wire  RetimeWrapper_457_clock; // @[package.scala 93:22:@57476.4]
  wire  RetimeWrapper_457_reset; // @[package.scala 93:22:@57476.4]
  wire  RetimeWrapper_457_io_flow; // @[package.scala 93:22:@57476.4]
  wire  RetimeWrapper_457_io_in; // @[package.scala 93:22:@57476.4]
  wire  RetimeWrapper_457_io_out; // @[package.scala 93:22:@57476.4]
  wire  RetimeWrapper_458_clock; // @[package.scala 93:22:@57484.4]
  wire  RetimeWrapper_458_reset; // @[package.scala 93:22:@57484.4]
  wire  RetimeWrapper_458_io_flow; // @[package.scala 93:22:@57484.4]
  wire  RetimeWrapper_458_io_in; // @[package.scala 93:22:@57484.4]
  wire  RetimeWrapper_458_io_out; // @[package.scala 93:22:@57484.4]
  wire  RetimeWrapper_459_clock; // @[package.scala 93:22:@57492.4]
  wire  RetimeWrapper_459_reset; // @[package.scala 93:22:@57492.4]
  wire  RetimeWrapper_459_io_flow; // @[package.scala 93:22:@57492.4]
  wire  RetimeWrapper_459_io_in; // @[package.scala 93:22:@57492.4]
  wire  RetimeWrapper_459_io_out; // @[package.scala 93:22:@57492.4]
  wire  RetimeWrapper_460_clock; // @[package.scala 93:22:@57580.4]
  wire  RetimeWrapper_460_reset; // @[package.scala 93:22:@57580.4]
  wire  RetimeWrapper_460_io_flow; // @[package.scala 93:22:@57580.4]
  wire  RetimeWrapper_460_io_in; // @[package.scala 93:22:@57580.4]
  wire  RetimeWrapper_460_io_out; // @[package.scala 93:22:@57580.4]
  wire  RetimeWrapper_461_clock; // @[package.scala 93:22:@57588.4]
  wire  RetimeWrapper_461_reset; // @[package.scala 93:22:@57588.4]
  wire  RetimeWrapper_461_io_flow; // @[package.scala 93:22:@57588.4]
  wire  RetimeWrapper_461_io_in; // @[package.scala 93:22:@57588.4]
  wire  RetimeWrapper_461_io_out; // @[package.scala 93:22:@57588.4]
  wire  RetimeWrapper_462_clock; // @[package.scala 93:22:@57596.4]
  wire  RetimeWrapper_462_reset; // @[package.scala 93:22:@57596.4]
  wire  RetimeWrapper_462_io_flow; // @[package.scala 93:22:@57596.4]
  wire  RetimeWrapper_462_io_in; // @[package.scala 93:22:@57596.4]
  wire  RetimeWrapper_462_io_out; // @[package.scala 93:22:@57596.4]
  wire  RetimeWrapper_463_clock; // @[package.scala 93:22:@57604.4]
  wire  RetimeWrapper_463_reset; // @[package.scala 93:22:@57604.4]
  wire  RetimeWrapper_463_io_flow; // @[package.scala 93:22:@57604.4]
  wire  RetimeWrapper_463_io_in; // @[package.scala 93:22:@57604.4]
  wire  RetimeWrapper_463_io_out; // @[package.scala 93:22:@57604.4]
  wire  RetimeWrapper_464_clock; // @[package.scala 93:22:@57612.4]
  wire  RetimeWrapper_464_reset; // @[package.scala 93:22:@57612.4]
  wire  RetimeWrapper_464_io_flow; // @[package.scala 93:22:@57612.4]
  wire  RetimeWrapper_464_io_in; // @[package.scala 93:22:@57612.4]
  wire  RetimeWrapper_464_io_out; // @[package.scala 93:22:@57612.4]
  wire  RetimeWrapper_465_clock; // @[package.scala 93:22:@57620.4]
  wire  RetimeWrapper_465_reset; // @[package.scala 93:22:@57620.4]
  wire  RetimeWrapper_465_io_flow; // @[package.scala 93:22:@57620.4]
  wire  RetimeWrapper_465_io_in; // @[package.scala 93:22:@57620.4]
  wire  RetimeWrapper_465_io_out; // @[package.scala 93:22:@57620.4]
  wire  RetimeWrapper_466_clock; // @[package.scala 93:22:@57628.4]
  wire  RetimeWrapper_466_reset; // @[package.scala 93:22:@57628.4]
  wire  RetimeWrapper_466_io_flow; // @[package.scala 93:22:@57628.4]
  wire  RetimeWrapper_466_io_in; // @[package.scala 93:22:@57628.4]
  wire  RetimeWrapper_466_io_out; // @[package.scala 93:22:@57628.4]
  wire  RetimeWrapper_467_clock; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_467_reset; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_467_io_flow; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_467_io_in; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_467_io_out; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_468_clock; // @[package.scala 93:22:@57644.4]
  wire  RetimeWrapper_468_reset; // @[package.scala 93:22:@57644.4]
  wire  RetimeWrapper_468_io_flow; // @[package.scala 93:22:@57644.4]
  wire  RetimeWrapper_468_io_in; // @[package.scala 93:22:@57644.4]
  wire  RetimeWrapper_468_io_out; // @[package.scala 93:22:@57644.4]
  wire  RetimeWrapper_469_clock; // @[package.scala 93:22:@57652.4]
  wire  RetimeWrapper_469_reset; // @[package.scala 93:22:@57652.4]
  wire  RetimeWrapper_469_io_flow; // @[package.scala 93:22:@57652.4]
  wire  RetimeWrapper_469_io_in; // @[package.scala 93:22:@57652.4]
  wire  RetimeWrapper_469_io_out; // @[package.scala 93:22:@57652.4]
  wire  RetimeWrapper_470_clock; // @[package.scala 93:22:@57660.4]
  wire  RetimeWrapper_470_reset; // @[package.scala 93:22:@57660.4]
  wire  RetimeWrapper_470_io_flow; // @[package.scala 93:22:@57660.4]
  wire  RetimeWrapper_470_io_in; // @[package.scala 93:22:@57660.4]
  wire  RetimeWrapper_470_io_out; // @[package.scala 93:22:@57660.4]
  wire  RetimeWrapper_471_clock; // @[package.scala 93:22:@57668.4]
  wire  RetimeWrapper_471_reset; // @[package.scala 93:22:@57668.4]
  wire  RetimeWrapper_471_io_flow; // @[package.scala 93:22:@57668.4]
  wire  RetimeWrapper_471_io_in; // @[package.scala 93:22:@57668.4]
  wire  RetimeWrapper_471_io_out; // @[package.scala 93:22:@57668.4]
  wire  RetimeWrapper_472_clock; // @[package.scala 93:22:@57676.4]
  wire  RetimeWrapper_472_reset; // @[package.scala 93:22:@57676.4]
  wire  RetimeWrapper_472_io_flow; // @[package.scala 93:22:@57676.4]
  wire  RetimeWrapper_472_io_in; // @[package.scala 93:22:@57676.4]
  wire  RetimeWrapper_472_io_out; // @[package.scala 93:22:@57676.4]
  wire  RetimeWrapper_473_clock; // @[package.scala 93:22:@57684.4]
  wire  RetimeWrapper_473_reset; // @[package.scala 93:22:@57684.4]
  wire  RetimeWrapper_473_io_flow; // @[package.scala 93:22:@57684.4]
  wire  RetimeWrapper_473_io_in; // @[package.scala 93:22:@57684.4]
  wire  RetimeWrapper_473_io_out; // @[package.scala 93:22:@57684.4]
  wire  RetimeWrapper_474_clock; // @[package.scala 93:22:@57692.4]
  wire  RetimeWrapper_474_reset; // @[package.scala 93:22:@57692.4]
  wire  RetimeWrapper_474_io_flow; // @[package.scala 93:22:@57692.4]
  wire  RetimeWrapper_474_io_in; // @[package.scala 93:22:@57692.4]
  wire  RetimeWrapper_474_io_out; // @[package.scala 93:22:@57692.4]
  wire  RetimeWrapper_475_clock; // @[package.scala 93:22:@57700.4]
  wire  RetimeWrapper_475_reset; // @[package.scala 93:22:@57700.4]
  wire  RetimeWrapper_475_io_flow; // @[package.scala 93:22:@57700.4]
  wire  RetimeWrapper_475_io_in; // @[package.scala 93:22:@57700.4]
  wire  RetimeWrapper_475_io_out; // @[package.scala 93:22:@57700.4]
  wire  RetimeWrapper_476_clock; // @[package.scala 93:22:@57708.4]
  wire  RetimeWrapper_476_reset; // @[package.scala 93:22:@57708.4]
  wire  RetimeWrapper_476_io_flow; // @[package.scala 93:22:@57708.4]
  wire  RetimeWrapper_476_io_in; // @[package.scala 93:22:@57708.4]
  wire  RetimeWrapper_476_io_out; // @[package.scala 93:22:@57708.4]
  wire  RetimeWrapper_477_clock; // @[package.scala 93:22:@57716.4]
  wire  RetimeWrapper_477_reset; // @[package.scala 93:22:@57716.4]
  wire  RetimeWrapper_477_io_flow; // @[package.scala 93:22:@57716.4]
  wire  RetimeWrapper_477_io_in; // @[package.scala 93:22:@57716.4]
  wire  RetimeWrapper_477_io_out; // @[package.scala 93:22:@57716.4]
  wire  RetimeWrapper_478_clock; // @[package.scala 93:22:@57724.4]
  wire  RetimeWrapper_478_reset; // @[package.scala 93:22:@57724.4]
  wire  RetimeWrapper_478_io_flow; // @[package.scala 93:22:@57724.4]
  wire  RetimeWrapper_478_io_in; // @[package.scala 93:22:@57724.4]
  wire  RetimeWrapper_478_io_out; // @[package.scala 93:22:@57724.4]
  wire  RetimeWrapper_479_clock; // @[package.scala 93:22:@57732.4]
  wire  RetimeWrapper_479_reset; // @[package.scala 93:22:@57732.4]
  wire  RetimeWrapper_479_io_flow; // @[package.scala 93:22:@57732.4]
  wire  RetimeWrapper_479_io_in; // @[package.scala 93:22:@57732.4]
  wire  RetimeWrapper_479_io_out; // @[package.scala 93:22:@57732.4]
  wire  RetimeWrapper_480_clock; // @[package.scala 93:22:@57820.4]
  wire  RetimeWrapper_480_reset; // @[package.scala 93:22:@57820.4]
  wire  RetimeWrapper_480_io_flow; // @[package.scala 93:22:@57820.4]
  wire  RetimeWrapper_480_io_in; // @[package.scala 93:22:@57820.4]
  wire  RetimeWrapper_480_io_out; // @[package.scala 93:22:@57820.4]
  wire  RetimeWrapper_481_clock; // @[package.scala 93:22:@57828.4]
  wire  RetimeWrapper_481_reset; // @[package.scala 93:22:@57828.4]
  wire  RetimeWrapper_481_io_flow; // @[package.scala 93:22:@57828.4]
  wire  RetimeWrapper_481_io_in; // @[package.scala 93:22:@57828.4]
  wire  RetimeWrapper_481_io_out; // @[package.scala 93:22:@57828.4]
  wire  RetimeWrapper_482_clock; // @[package.scala 93:22:@57836.4]
  wire  RetimeWrapper_482_reset; // @[package.scala 93:22:@57836.4]
  wire  RetimeWrapper_482_io_flow; // @[package.scala 93:22:@57836.4]
  wire  RetimeWrapper_482_io_in; // @[package.scala 93:22:@57836.4]
  wire  RetimeWrapper_482_io_out; // @[package.scala 93:22:@57836.4]
  wire  RetimeWrapper_483_clock; // @[package.scala 93:22:@57844.4]
  wire  RetimeWrapper_483_reset; // @[package.scala 93:22:@57844.4]
  wire  RetimeWrapper_483_io_flow; // @[package.scala 93:22:@57844.4]
  wire  RetimeWrapper_483_io_in; // @[package.scala 93:22:@57844.4]
  wire  RetimeWrapper_483_io_out; // @[package.scala 93:22:@57844.4]
  wire  RetimeWrapper_484_clock; // @[package.scala 93:22:@57852.4]
  wire  RetimeWrapper_484_reset; // @[package.scala 93:22:@57852.4]
  wire  RetimeWrapper_484_io_flow; // @[package.scala 93:22:@57852.4]
  wire  RetimeWrapper_484_io_in; // @[package.scala 93:22:@57852.4]
  wire  RetimeWrapper_484_io_out; // @[package.scala 93:22:@57852.4]
  wire  RetimeWrapper_485_clock; // @[package.scala 93:22:@57860.4]
  wire  RetimeWrapper_485_reset; // @[package.scala 93:22:@57860.4]
  wire  RetimeWrapper_485_io_flow; // @[package.scala 93:22:@57860.4]
  wire  RetimeWrapper_485_io_in; // @[package.scala 93:22:@57860.4]
  wire  RetimeWrapper_485_io_out; // @[package.scala 93:22:@57860.4]
  wire  RetimeWrapper_486_clock; // @[package.scala 93:22:@57868.4]
  wire  RetimeWrapper_486_reset; // @[package.scala 93:22:@57868.4]
  wire  RetimeWrapper_486_io_flow; // @[package.scala 93:22:@57868.4]
  wire  RetimeWrapper_486_io_in; // @[package.scala 93:22:@57868.4]
  wire  RetimeWrapper_486_io_out; // @[package.scala 93:22:@57868.4]
  wire  RetimeWrapper_487_clock; // @[package.scala 93:22:@57876.4]
  wire  RetimeWrapper_487_reset; // @[package.scala 93:22:@57876.4]
  wire  RetimeWrapper_487_io_flow; // @[package.scala 93:22:@57876.4]
  wire  RetimeWrapper_487_io_in; // @[package.scala 93:22:@57876.4]
  wire  RetimeWrapper_487_io_out; // @[package.scala 93:22:@57876.4]
  wire  RetimeWrapper_488_clock; // @[package.scala 93:22:@57884.4]
  wire  RetimeWrapper_488_reset; // @[package.scala 93:22:@57884.4]
  wire  RetimeWrapper_488_io_flow; // @[package.scala 93:22:@57884.4]
  wire  RetimeWrapper_488_io_in; // @[package.scala 93:22:@57884.4]
  wire  RetimeWrapper_488_io_out; // @[package.scala 93:22:@57884.4]
  wire  RetimeWrapper_489_clock; // @[package.scala 93:22:@57892.4]
  wire  RetimeWrapper_489_reset; // @[package.scala 93:22:@57892.4]
  wire  RetimeWrapper_489_io_flow; // @[package.scala 93:22:@57892.4]
  wire  RetimeWrapper_489_io_in; // @[package.scala 93:22:@57892.4]
  wire  RetimeWrapper_489_io_out; // @[package.scala 93:22:@57892.4]
  wire  RetimeWrapper_490_clock; // @[package.scala 93:22:@57900.4]
  wire  RetimeWrapper_490_reset; // @[package.scala 93:22:@57900.4]
  wire  RetimeWrapper_490_io_flow; // @[package.scala 93:22:@57900.4]
  wire  RetimeWrapper_490_io_in; // @[package.scala 93:22:@57900.4]
  wire  RetimeWrapper_490_io_out; // @[package.scala 93:22:@57900.4]
  wire  RetimeWrapper_491_clock; // @[package.scala 93:22:@57908.4]
  wire  RetimeWrapper_491_reset; // @[package.scala 93:22:@57908.4]
  wire  RetimeWrapper_491_io_flow; // @[package.scala 93:22:@57908.4]
  wire  RetimeWrapper_491_io_in; // @[package.scala 93:22:@57908.4]
  wire  RetimeWrapper_491_io_out; // @[package.scala 93:22:@57908.4]
  wire  RetimeWrapper_492_clock; // @[package.scala 93:22:@57916.4]
  wire  RetimeWrapper_492_reset; // @[package.scala 93:22:@57916.4]
  wire  RetimeWrapper_492_io_flow; // @[package.scala 93:22:@57916.4]
  wire  RetimeWrapper_492_io_in; // @[package.scala 93:22:@57916.4]
  wire  RetimeWrapper_492_io_out; // @[package.scala 93:22:@57916.4]
  wire  RetimeWrapper_493_clock; // @[package.scala 93:22:@57924.4]
  wire  RetimeWrapper_493_reset; // @[package.scala 93:22:@57924.4]
  wire  RetimeWrapper_493_io_flow; // @[package.scala 93:22:@57924.4]
  wire  RetimeWrapper_493_io_in; // @[package.scala 93:22:@57924.4]
  wire  RetimeWrapper_493_io_out; // @[package.scala 93:22:@57924.4]
  wire  RetimeWrapper_494_clock; // @[package.scala 93:22:@57932.4]
  wire  RetimeWrapper_494_reset; // @[package.scala 93:22:@57932.4]
  wire  RetimeWrapper_494_io_flow; // @[package.scala 93:22:@57932.4]
  wire  RetimeWrapper_494_io_in; // @[package.scala 93:22:@57932.4]
  wire  RetimeWrapper_494_io_out; // @[package.scala 93:22:@57932.4]
  wire  RetimeWrapper_495_clock; // @[package.scala 93:22:@57940.4]
  wire  RetimeWrapper_495_reset; // @[package.scala 93:22:@57940.4]
  wire  RetimeWrapper_495_io_flow; // @[package.scala 93:22:@57940.4]
  wire  RetimeWrapper_495_io_in; // @[package.scala 93:22:@57940.4]
  wire  RetimeWrapper_495_io_out; // @[package.scala 93:22:@57940.4]
  wire  RetimeWrapper_496_clock; // @[package.scala 93:22:@57948.4]
  wire  RetimeWrapper_496_reset; // @[package.scala 93:22:@57948.4]
  wire  RetimeWrapper_496_io_flow; // @[package.scala 93:22:@57948.4]
  wire  RetimeWrapper_496_io_in; // @[package.scala 93:22:@57948.4]
  wire  RetimeWrapper_496_io_out; // @[package.scala 93:22:@57948.4]
  wire  RetimeWrapper_497_clock; // @[package.scala 93:22:@57956.4]
  wire  RetimeWrapper_497_reset; // @[package.scala 93:22:@57956.4]
  wire  RetimeWrapper_497_io_flow; // @[package.scala 93:22:@57956.4]
  wire  RetimeWrapper_497_io_in; // @[package.scala 93:22:@57956.4]
  wire  RetimeWrapper_497_io_out; // @[package.scala 93:22:@57956.4]
  wire  RetimeWrapper_498_clock; // @[package.scala 93:22:@57964.4]
  wire  RetimeWrapper_498_reset; // @[package.scala 93:22:@57964.4]
  wire  RetimeWrapper_498_io_flow; // @[package.scala 93:22:@57964.4]
  wire  RetimeWrapper_498_io_in; // @[package.scala 93:22:@57964.4]
  wire  RetimeWrapper_498_io_out; // @[package.scala 93:22:@57964.4]
  wire  RetimeWrapper_499_clock; // @[package.scala 93:22:@57972.4]
  wire  RetimeWrapper_499_reset; // @[package.scala 93:22:@57972.4]
  wire  RetimeWrapper_499_io_flow; // @[package.scala 93:22:@57972.4]
  wire  RetimeWrapper_499_io_in; // @[package.scala 93:22:@57972.4]
  wire  RetimeWrapper_499_io_out; // @[package.scala 93:22:@57972.4]
  wire  RetimeWrapper_500_clock; // @[package.scala 93:22:@58060.4]
  wire  RetimeWrapper_500_reset; // @[package.scala 93:22:@58060.4]
  wire  RetimeWrapper_500_io_flow; // @[package.scala 93:22:@58060.4]
  wire  RetimeWrapper_500_io_in; // @[package.scala 93:22:@58060.4]
  wire  RetimeWrapper_500_io_out; // @[package.scala 93:22:@58060.4]
  wire  RetimeWrapper_501_clock; // @[package.scala 93:22:@58068.4]
  wire  RetimeWrapper_501_reset; // @[package.scala 93:22:@58068.4]
  wire  RetimeWrapper_501_io_flow; // @[package.scala 93:22:@58068.4]
  wire  RetimeWrapper_501_io_in; // @[package.scala 93:22:@58068.4]
  wire  RetimeWrapper_501_io_out; // @[package.scala 93:22:@58068.4]
  wire  RetimeWrapper_502_clock; // @[package.scala 93:22:@58076.4]
  wire  RetimeWrapper_502_reset; // @[package.scala 93:22:@58076.4]
  wire  RetimeWrapper_502_io_flow; // @[package.scala 93:22:@58076.4]
  wire  RetimeWrapper_502_io_in; // @[package.scala 93:22:@58076.4]
  wire  RetimeWrapper_502_io_out; // @[package.scala 93:22:@58076.4]
  wire  RetimeWrapper_503_clock; // @[package.scala 93:22:@58084.4]
  wire  RetimeWrapper_503_reset; // @[package.scala 93:22:@58084.4]
  wire  RetimeWrapper_503_io_flow; // @[package.scala 93:22:@58084.4]
  wire  RetimeWrapper_503_io_in; // @[package.scala 93:22:@58084.4]
  wire  RetimeWrapper_503_io_out; // @[package.scala 93:22:@58084.4]
  wire  RetimeWrapper_504_clock; // @[package.scala 93:22:@58092.4]
  wire  RetimeWrapper_504_reset; // @[package.scala 93:22:@58092.4]
  wire  RetimeWrapper_504_io_flow; // @[package.scala 93:22:@58092.4]
  wire  RetimeWrapper_504_io_in; // @[package.scala 93:22:@58092.4]
  wire  RetimeWrapper_504_io_out; // @[package.scala 93:22:@58092.4]
  wire  RetimeWrapper_505_clock; // @[package.scala 93:22:@58100.4]
  wire  RetimeWrapper_505_reset; // @[package.scala 93:22:@58100.4]
  wire  RetimeWrapper_505_io_flow; // @[package.scala 93:22:@58100.4]
  wire  RetimeWrapper_505_io_in; // @[package.scala 93:22:@58100.4]
  wire  RetimeWrapper_505_io_out; // @[package.scala 93:22:@58100.4]
  wire  RetimeWrapper_506_clock; // @[package.scala 93:22:@58108.4]
  wire  RetimeWrapper_506_reset; // @[package.scala 93:22:@58108.4]
  wire  RetimeWrapper_506_io_flow; // @[package.scala 93:22:@58108.4]
  wire  RetimeWrapper_506_io_in; // @[package.scala 93:22:@58108.4]
  wire  RetimeWrapper_506_io_out; // @[package.scala 93:22:@58108.4]
  wire  RetimeWrapper_507_clock; // @[package.scala 93:22:@58116.4]
  wire  RetimeWrapper_507_reset; // @[package.scala 93:22:@58116.4]
  wire  RetimeWrapper_507_io_flow; // @[package.scala 93:22:@58116.4]
  wire  RetimeWrapper_507_io_in; // @[package.scala 93:22:@58116.4]
  wire  RetimeWrapper_507_io_out; // @[package.scala 93:22:@58116.4]
  wire  RetimeWrapper_508_clock; // @[package.scala 93:22:@58124.4]
  wire  RetimeWrapper_508_reset; // @[package.scala 93:22:@58124.4]
  wire  RetimeWrapper_508_io_flow; // @[package.scala 93:22:@58124.4]
  wire  RetimeWrapper_508_io_in; // @[package.scala 93:22:@58124.4]
  wire  RetimeWrapper_508_io_out; // @[package.scala 93:22:@58124.4]
  wire  RetimeWrapper_509_clock; // @[package.scala 93:22:@58132.4]
  wire  RetimeWrapper_509_reset; // @[package.scala 93:22:@58132.4]
  wire  RetimeWrapper_509_io_flow; // @[package.scala 93:22:@58132.4]
  wire  RetimeWrapper_509_io_in; // @[package.scala 93:22:@58132.4]
  wire  RetimeWrapper_509_io_out; // @[package.scala 93:22:@58132.4]
  wire  RetimeWrapper_510_clock; // @[package.scala 93:22:@58140.4]
  wire  RetimeWrapper_510_reset; // @[package.scala 93:22:@58140.4]
  wire  RetimeWrapper_510_io_flow; // @[package.scala 93:22:@58140.4]
  wire  RetimeWrapper_510_io_in; // @[package.scala 93:22:@58140.4]
  wire  RetimeWrapper_510_io_out; // @[package.scala 93:22:@58140.4]
  wire  RetimeWrapper_511_clock; // @[package.scala 93:22:@58148.4]
  wire  RetimeWrapper_511_reset; // @[package.scala 93:22:@58148.4]
  wire  RetimeWrapper_511_io_flow; // @[package.scala 93:22:@58148.4]
  wire  RetimeWrapper_511_io_in; // @[package.scala 93:22:@58148.4]
  wire  RetimeWrapper_511_io_out; // @[package.scala 93:22:@58148.4]
  wire  RetimeWrapper_512_clock; // @[package.scala 93:22:@58156.4]
  wire  RetimeWrapper_512_reset; // @[package.scala 93:22:@58156.4]
  wire  RetimeWrapper_512_io_flow; // @[package.scala 93:22:@58156.4]
  wire  RetimeWrapper_512_io_in; // @[package.scala 93:22:@58156.4]
  wire  RetimeWrapper_512_io_out; // @[package.scala 93:22:@58156.4]
  wire  RetimeWrapper_513_clock; // @[package.scala 93:22:@58164.4]
  wire  RetimeWrapper_513_reset; // @[package.scala 93:22:@58164.4]
  wire  RetimeWrapper_513_io_flow; // @[package.scala 93:22:@58164.4]
  wire  RetimeWrapper_513_io_in; // @[package.scala 93:22:@58164.4]
  wire  RetimeWrapper_513_io_out; // @[package.scala 93:22:@58164.4]
  wire  RetimeWrapper_514_clock; // @[package.scala 93:22:@58172.4]
  wire  RetimeWrapper_514_reset; // @[package.scala 93:22:@58172.4]
  wire  RetimeWrapper_514_io_flow; // @[package.scala 93:22:@58172.4]
  wire  RetimeWrapper_514_io_in; // @[package.scala 93:22:@58172.4]
  wire  RetimeWrapper_514_io_out; // @[package.scala 93:22:@58172.4]
  wire  RetimeWrapper_515_clock; // @[package.scala 93:22:@58180.4]
  wire  RetimeWrapper_515_reset; // @[package.scala 93:22:@58180.4]
  wire  RetimeWrapper_515_io_flow; // @[package.scala 93:22:@58180.4]
  wire  RetimeWrapper_515_io_in; // @[package.scala 93:22:@58180.4]
  wire  RetimeWrapper_515_io_out; // @[package.scala 93:22:@58180.4]
  wire  RetimeWrapper_516_clock; // @[package.scala 93:22:@58188.4]
  wire  RetimeWrapper_516_reset; // @[package.scala 93:22:@58188.4]
  wire  RetimeWrapper_516_io_flow; // @[package.scala 93:22:@58188.4]
  wire  RetimeWrapper_516_io_in; // @[package.scala 93:22:@58188.4]
  wire  RetimeWrapper_516_io_out; // @[package.scala 93:22:@58188.4]
  wire  RetimeWrapper_517_clock; // @[package.scala 93:22:@58196.4]
  wire  RetimeWrapper_517_reset; // @[package.scala 93:22:@58196.4]
  wire  RetimeWrapper_517_io_flow; // @[package.scala 93:22:@58196.4]
  wire  RetimeWrapper_517_io_in; // @[package.scala 93:22:@58196.4]
  wire  RetimeWrapper_517_io_out; // @[package.scala 93:22:@58196.4]
  wire  RetimeWrapper_518_clock; // @[package.scala 93:22:@58204.4]
  wire  RetimeWrapper_518_reset; // @[package.scala 93:22:@58204.4]
  wire  RetimeWrapper_518_io_flow; // @[package.scala 93:22:@58204.4]
  wire  RetimeWrapper_518_io_in; // @[package.scala 93:22:@58204.4]
  wire  RetimeWrapper_518_io_out; // @[package.scala 93:22:@58204.4]
  wire  RetimeWrapper_519_clock; // @[package.scala 93:22:@58212.4]
  wire  RetimeWrapper_519_reset; // @[package.scala 93:22:@58212.4]
  wire  RetimeWrapper_519_io_flow; // @[package.scala 93:22:@58212.4]
  wire  RetimeWrapper_519_io_in; // @[package.scala 93:22:@58212.4]
  wire  RetimeWrapper_519_io_out; // @[package.scala 93:22:@58212.4]
  wire  RetimeWrapper_520_clock; // @[package.scala 93:22:@58300.4]
  wire  RetimeWrapper_520_reset; // @[package.scala 93:22:@58300.4]
  wire  RetimeWrapper_520_io_flow; // @[package.scala 93:22:@58300.4]
  wire  RetimeWrapper_520_io_in; // @[package.scala 93:22:@58300.4]
  wire  RetimeWrapper_520_io_out; // @[package.scala 93:22:@58300.4]
  wire  RetimeWrapper_521_clock; // @[package.scala 93:22:@58308.4]
  wire  RetimeWrapper_521_reset; // @[package.scala 93:22:@58308.4]
  wire  RetimeWrapper_521_io_flow; // @[package.scala 93:22:@58308.4]
  wire  RetimeWrapper_521_io_in; // @[package.scala 93:22:@58308.4]
  wire  RetimeWrapper_521_io_out; // @[package.scala 93:22:@58308.4]
  wire  RetimeWrapper_522_clock; // @[package.scala 93:22:@58316.4]
  wire  RetimeWrapper_522_reset; // @[package.scala 93:22:@58316.4]
  wire  RetimeWrapper_522_io_flow; // @[package.scala 93:22:@58316.4]
  wire  RetimeWrapper_522_io_in; // @[package.scala 93:22:@58316.4]
  wire  RetimeWrapper_522_io_out; // @[package.scala 93:22:@58316.4]
  wire  RetimeWrapper_523_clock; // @[package.scala 93:22:@58324.4]
  wire  RetimeWrapper_523_reset; // @[package.scala 93:22:@58324.4]
  wire  RetimeWrapper_523_io_flow; // @[package.scala 93:22:@58324.4]
  wire  RetimeWrapper_523_io_in; // @[package.scala 93:22:@58324.4]
  wire  RetimeWrapper_523_io_out; // @[package.scala 93:22:@58324.4]
  wire  RetimeWrapper_524_clock; // @[package.scala 93:22:@58332.4]
  wire  RetimeWrapper_524_reset; // @[package.scala 93:22:@58332.4]
  wire  RetimeWrapper_524_io_flow; // @[package.scala 93:22:@58332.4]
  wire  RetimeWrapper_524_io_in; // @[package.scala 93:22:@58332.4]
  wire  RetimeWrapper_524_io_out; // @[package.scala 93:22:@58332.4]
  wire  RetimeWrapper_525_clock; // @[package.scala 93:22:@58340.4]
  wire  RetimeWrapper_525_reset; // @[package.scala 93:22:@58340.4]
  wire  RetimeWrapper_525_io_flow; // @[package.scala 93:22:@58340.4]
  wire  RetimeWrapper_525_io_in; // @[package.scala 93:22:@58340.4]
  wire  RetimeWrapper_525_io_out; // @[package.scala 93:22:@58340.4]
  wire  RetimeWrapper_526_clock; // @[package.scala 93:22:@58348.4]
  wire  RetimeWrapper_526_reset; // @[package.scala 93:22:@58348.4]
  wire  RetimeWrapper_526_io_flow; // @[package.scala 93:22:@58348.4]
  wire  RetimeWrapper_526_io_in; // @[package.scala 93:22:@58348.4]
  wire  RetimeWrapper_526_io_out; // @[package.scala 93:22:@58348.4]
  wire  RetimeWrapper_527_clock; // @[package.scala 93:22:@58356.4]
  wire  RetimeWrapper_527_reset; // @[package.scala 93:22:@58356.4]
  wire  RetimeWrapper_527_io_flow; // @[package.scala 93:22:@58356.4]
  wire  RetimeWrapper_527_io_in; // @[package.scala 93:22:@58356.4]
  wire  RetimeWrapper_527_io_out; // @[package.scala 93:22:@58356.4]
  wire  RetimeWrapper_528_clock; // @[package.scala 93:22:@58364.4]
  wire  RetimeWrapper_528_reset; // @[package.scala 93:22:@58364.4]
  wire  RetimeWrapper_528_io_flow; // @[package.scala 93:22:@58364.4]
  wire  RetimeWrapper_528_io_in; // @[package.scala 93:22:@58364.4]
  wire  RetimeWrapper_528_io_out; // @[package.scala 93:22:@58364.4]
  wire  RetimeWrapper_529_clock; // @[package.scala 93:22:@58372.4]
  wire  RetimeWrapper_529_reset; // @[package.scala 93:22:@58372.4]
  wire  RetimeWrapper_529_io_flow; // @[package.scala 93:22:@58372.4]
  wire  RetimeWrapper_529_io_in; // @[package.scala 93:22:@58372.4]
  wire  RetimeWrapper_529_io_out; // @[package.scala 93:22:@58372.4]
  wire  RetimeWrapper_530_clock; // @[package.scala 93:22:@58380.4]
  wire  RetimeWrapper_530_reset; // @[package.scala 93:22:@58380.4]
  wire  RetimeWrapper_530_io_flow; // @[package.scala 93:22:@58380.4]
  wire  RetimeWrapper_530_io_in; // @[package.scala 93:22:@58380.4]
  wire  RetimeWrapper_530_io_out; // @[package.scala 93:22:@58380.4]
  wire  RetimeWrapper_531_clock; // @[package.scala 93:22:@58388.4]
  wire  RetimeWrapper_531_reset; // @[package.scala 93:22:@58388.4]
  wire  RetimeWrapper_531_io_flow; // @[package.scala 93:22:@58388.4]
  wire  RetimeWrapper_531_io_in; // @[package.scala 93:22:@58388.4]
  wire  RetimeWrapper_531_io_out; // @[package.scala 93:22:@58388.4]
  wire  RetimeWrapper_532_clock; // @[package.scala 93:22:@58396.4]
  wire  RetimeWrapper_532_reset; // @[package.scala 93:22:@58396.4]
  wire  RetimeWrapper_532_io_flow; // @[package.scala 93:22:@58396.4]
  wire  RetimeWrapper_532_io_in; // @[package.scala 93:22:@58396.4]
  wire  RetimeWrapper_532_io_out; // @[package.scala 93:22:@58396.4]
  wire  RetimeWrapper_533_clock; // @[package.scala 93:22:@58404.4]
  wire  RetimeWrapper_533_reset; // @[package.scala 93:22:@58404.4]
  wire  RetimeWrapper_533_io_flow; // @[package.scala 93:22:@58404.4]
  wire  RetimeWrapper_533_io_in; // @[package.scala 93:22:@58404.4]
  wire  RetimeWrapper_533_io_out; // @[package.scala 93:22:@58404.4]
  wire  RetimeWrapper_534_clock; // @[package.scala 93:22:@58412.4]
  wire  RetimeWrapper_534_reset; // @[package.scala 93:22:@58412.4]
  wire  RetimeWrapper_534_io_flow; // @[package.scala 93:22:@58412.4]
  wire  RetimeWrapper_534_io_in; // @[package.scala 93:22:@58412.4]
  wire  RetimeWrapper_534_io_out; // @[package.scala 93:22:@58412.4]
  wire  RetimeWrapper_535_clock; // @[package.scala 93:22:@58420.4]
  wire  RetimeWrapper_535_reset; // @[package.scala 93:22:@58420.4]
  wire  RetimeWrapper_535_io_flow; // @[package.scala 93:22:@58420.4]
  wire  RetimeWrapper_535_io_in; // @[package.scala 93:22:@58420.4]
  wire  RetimeWrapper_535_io_out; // @[package.scala 93:22:@58420.4]
  wire  RetimeWrapper_536_clock; // @[package.scala 93:22:@58428.4]
  wire  RetimeWrapper_536_reset; // @[package.scala 93:22:@58428.4]
  wire  RetimeWrapper_536_io_flow; // @[package.scala 93:22:@58428.4]
  wire  RetimeWrapper_536_io_in; // @[package.scala 93:22:@58428.4]
  wire  RetimeWrapper_536_io_out; // @[package.scala 93:22:@58428.4]
  wire  RetimeWrapper_537_clock; // @[package.scala 93:22:@58436.4]
  wire  RetimeWrapper_537_reset; // @[package.scala 93:22:@58436.4]
  wire  RetimeWrapper_537_io_flow; // @[package.scala 93:22:@58436.4]
  wire  RetimeWrapper_537_io_in; // @[package.scala 93:22:@58436.4]
  wire  RetimeWrapper_537_io_out; // @[package.scala 93:22:@58436.4]
  wire  RetimeWrapper_538_clock; // @[package.scala 93:22:@58444.4]
  wire  RetimeWrapper_538_reset; // @[package.scala 93:22:@58444.4]
  wire  RetimeWrapper_538_io_flow; // @[package.scala 93:22:@58444.4]
  wire  RetimeWrapper_538_io_in; // @[package.scala 93:22:@58444.4]
  wire  RetimeWrapper_538_io_out; // @[package.scala 93:22:@58444.4]
  wire  RetimeWrapper_539_clock; // @[package.scala 93:22:@58452.4]
  wire  RetimeWrapper_539_reset; // @[package.scala 93:22:@58452.4]
  wire  RetimeWrapper_539_io_flow; // @[package.scala 93:22:@58452.4]
  wire  RetimeWrapper_539_io_in; // @[package.scala 93:22:@58452.4]
  wire  RetimeWrapper_539_io_out; // @[package.scala 93:22:@58452.4]
  wire  RetimeWrapper_540_clock; // @[package.scala 93:22:@58540.4]
  wire  RetimeWrapper_540_reset; // @[package.scala 93:22:@58540.4]
  wire  RetimeWrapper_540_io_flow; // @[package.scala 93:22:@58540.4]
  wire  RetimeWrapper_540_io_in; // @[package.scala 93:22:@58540.4]
  wire  RetimeWrapper_540_io_out; // @[package.scala 93:22:@58540.4]
  wire  RetimeWrapper_541_clock; // @[package.scala 93:22:@58548.4]
  wire  RetimeWrapper_541_reset; // @[package.scala 93:22:@58548.4]
  wire  RetimeWrapper_541_io_flow; // @[package.scala 93:22:@58548.4]
  wire  RetimeWrapper_541_io_in; // @[package.scala 93:22:@58548.4]
  wire  RetimeWrapper_541_io_out; // @[package.scala 93:22:@58548.4]
  wire  RetimeWrapper_542_clock; // @[package.scala 93:22:@58556.4]
  wire  RetimeWrapper_542_reset; // @[package.scala 93:22:@58556.4]
  wire  RetimeWrapper_542_io_flow; // @[package.scala 93:22:@58556.4]
  wire  RetimeWrapper_542_io_in; // @[package.scala 93:22:@58556.4]
  wire  RetimeWrapper_542_io_out; // @[package.scala 93:22:@58556.4]
  wire  RetimeWrapper_543_clock; // @[package.scala 93:22:@58564.4]
  wire  RetimeWrapper_543_reset; // @[package.scala 93:22:@58564.4]
  wire  RetimeWrapper_543_io_flow; // @[package.scala 93:22:@58564.4]
  wire  RetimeWrapper_543_io_in; // @[package.scala 93:22:@58564.4]
  wire  RetimeWrapper_543_io_out; // @[package.scala 93:22:@58564.4]
  wire  RetimeWrapper_544_clock; // @[package.scala 93:22:@58572.4]
  wire  RetimeWrapper_544_reset; // @[package.scala 93:22:@58572.4]
  wire  RetimeWrapper_544_io_flow; // @[package.scala 93:22:@58572.4]
  wire  RetimeWrapper_544_io_in; // @[package.scala 93:22:@58572.4]
  wire  RetimeWrapper_544_io_out; // @[package.scala 93:22:@58572.4]
  wire  RetimeWrapper_545_clock; // @[package.scala 93:22:@58580.4]
  wire  RetimeWrapper_545_reset; // @[package.scala 93:22:@58580.4]
  wire  RetimeWrapper_545_io_flow; // @[package.scala 93:22:@58580.4]
  wire  RetimeWrapper_545_io_in; // @[package.scala 93:22:@58580.4]
  wire  RetimeWrapper_545_io_out; // @[package.scala 93:22:@58580.4]
  wire  RetimeWrapper_546_clock; // @[package.scala 93:22:@58588.4]
  wire  RetimeWrapper_546_reset; // @[package.scala 93:22:@58588.4]
  wire  RetimeWrapper_546_io_flow; // @[package.scala 93:22:@58588.4]
  wire  RetimeWrapper_546_io_in; // @[package.scala 93:22:@58588.4]
  wire  RetimeWrapper_546_io_out; // @[package.scala 93:22:@58588.4]
  wire  RetimeWrapper_547_clock; // @[package.scala 93:22:@58596.4]
  wire  RetimeWrapper_547_reset; // @[package.scala 93:22:@58596.4]
  wire  RetimeWrapper_547_io_flow; // @[package.scala 93:22:@58596.4]
  wire  RetimeWrapper_547_io_in; // @[package.scala 93:22:@58596.4]
  wire  RetimeWrapper_547_io_out; // @[package.scala 93:22:@58596.4]
  wire  RetimeWrapper_548_clock; // @[package.scala 93:22:@58604.4]
  wire  RetimeWrapper_548_reset; // @[package.scala 93:22:@58604.4]
  wire  RetimeWrapper_548_io_flow; // @[package.scala 93:22:@58604.4]
  wire  RetimeWrapper_548_io_in; // @[package.scala 93:22:@58604.4]
  wire  RetimeWrapper_548_io_out; // @[package.scala 93:22:@58604.4]
  wire  RetimeWrapper_549_clock; // @[package.scala 93:22:@58612.4]
  wire  RetimeWrapper_549_reset; // @[package.scala 93:22:@58612.4]
  wire  RetimeWrapper_549_io_flow; // @[package.scala 93:22:@58612.4]
  wire  RetimeWrapper_549_io_in; // @[package.scala 93:22:@58612.4]
  wire  RetimeWrapper_549_io_out; // @[package.scala 93:22:@58612.4]
  wire  RetimeWrapper_550_clock; // @[package.scala 93:22:@58620.4]
  wire  RetimeWrapper_550_reset; // @[package.scala 93:22:@58620.4]
  wire  RetimeWrapper_550_io_flow; // @[package.scala 93:22:@58620.4]
  wire  RetimeWrapper_550_io_in; // @[package.scala 93:22:@58620.4]
  wire  RetimeWrapper_550_io_out; // @[package.scala 93:22:@58620.4]
  wire  RetimeWrapper_551_clock; // @[package.scala 93:22:@58628.4]
  wire  RetimeWrapper_551_reset; // @[package.scala 93:22:@58628.4]
  wire  RetimeWrapper_551_io_flow; // @[package.scala 93:22:@58628.4]
  wire  RetimeWrapper_551_io_in; // @[package.scala 93:22:@58628.4]
  wire  RetimeWrapper_551_io_out; // @[package.scala 93:22:@58628.4]
  wire  RetimeWrapper_552_clock; // @[package.scala 93:22:@58636.4]
  wire  RetimeWrapper_552_reset; // @[package.scala 93:22:@58636.4]
  wire  RetimeWrapper_552_io_flow; // @[package.scala 93:22:@58636.4]
  wire  RetimeWrapper_552_io_in; // @[package.scala 93:22:@58636.4]
  wire  RetimeWrapper_552_io_out; // @[package.scala 93:22:@58636.4]
  wire  RetimeWrapper_553_clock; // @[package.scala 93:22:@58644.4]
  wire  RetimeWrapper_553_reset; // @[package.scala 93:22:@58644.4]
  wire  RetimeWrapper_553_io_flow; // @[package.scala 93:22:@58644.4]
  wire  RetimeWrapper_553_io_in; // @[package.scala 93:22:@58644.4]
  wire  RetimeWrapper_553_io_out; // @[package.scala 93:22:@58644.4]
  wire  RetimeWrapper_554_clock; // @[package.scala 93:22:@58652.4]
  wire  RetimeWrapper_554_reset; // @[package.scala 93:22:@58652.4]
  wire  RetimeWrapper_554_io_flow; // @[package.scala 93:22:@58652.4]
  wire  RetimeWrapper_554_io_in; // @[package.scala 93:22:@58652.4]
  wire  RetimeWrapper_554_io_out; // @[package.scala 93:22:@58652.4]
  wire  RetimeWrapper_555_clock; // @[package.scala 93:22:@58660.4]
  wire  RetimeWrapper_555_reset; // @[package.scala 93:22:@58660.4]
  wire  RetimeWrapper_555_io_flow; // @[package.scala 93:22:@58660.4]
  wire  RetimeWrapper_555_io_in; // @[package.scala 93:22:@58660.4]
  wire  RetimeWrapper_555_io_out; // @[package.scala 93:22:@58660.4]
  wire  RetimeWrapper_556_clock; // @[package.scala 93:22:@58668.4]
  wire  RetimeWrapper_556_reset; // @[package.scala 93:22:@58668.4]
  wire  RetimeWrapper_556_io_flow; // @[package.scala 93:22:@58668.4]
  wire  RetimeWrapper_556_io_in; // @[package.scala 93:22:@58668.4]
  wire  RetimeWrapper_556_io_out; // @[package.scala 93:22:@58668.4]
  wire  RetimeWrapper_557_clock; // @[package.scala 93:22:@58676.4]
  wire  RetimeWrapper_557_reset; // @[package.scala 93:22:@58676.4]
  wire  RetimeWrapper_557_io_flow; // @[package.scala 93:22:@58676.4]
  wire  RetimeWrapper_557_io_in; // @[package.scala 93:22:@58676.4]
  wire  RetimeWrapper_557_io_out; // @[package.scala 93:22:@58676.4]
  wire  RetimeWrapper_558_clock; // @[package.scala 93:22:@58684.4]
  wire  RetimeWrapper_558_reset; // @[package.scala 93:22:@58684.4]
  wire  RetimeWrapper_558_io_flow; // @[package.scala 93:22:@58684.4]
  wire  RetimeWrapper_558_io_in; // @[package.scala 93:22:@58684.4]
  wire  RetimeWrapper_558_io_out; // @[package.scala 93:22:@58684.4]
  wire  RetimeWrapper_559_clock; // @[package.scala 93:22:@58692.4]
  wire  RetimeWrapper_559_reset; // @[package.scala 93:22:@58692.4]
  wire  RetimeWrapper_559_io_flow; // @[package.scala 93:22:@58692.4]
  wire  RetimeWrapper_559_io_in; // @[package.scala 93:22:@58692.4]
  wire  RetimeWrapper_559_io_out; // @[package.scala 93:22:@58692.4]
  wire  RetimeWrapper_560_clock; // @[package.scala 93:22:@58780.4]
  wire  RetimeWrapper_560_reset; // @[package.scala 93:22:@58780.4]
  wire  RetimeWrapper_560_io_flow; // @[package.scala 93:22:@58780.4]
  wire  RetimeWrapper_560_io_in; // @[package.scala 93:22:@58780.4]
  wire  RetimeWrapper_560_io_out; // @[package.scala 93:22:@58780.4]
  wire  RetimeWrapper_561_clock; // @[package.scala 93:22:@58788.4]
  wire  RetimeWrapper_561_reset; // @[package.scala 93:22:@58788.4]
  wire  RetimeWrapper_561_io_flow; // @[package.scala 93:22:@58788.4]
  wire  RetimeWrapper_561_io_in; // @[package.scala 93:22:@58788.4]
  wire  RetimeWrapper_561_io_out; // @[package.scala 93:22:@58788.4]
  wire  RetimeWrapper_562_clock; // @[package.scala 93:22:@58796.4]
  wire  RetimeWrapper_562_reset; // @[package.scala 93:22:@58796.4]
  wire  RetimeWrapper_562_io_flow; // @[package.scala 93:22:@58796.4]
  wire  RetimeWrapper_562_io_in; // @[package.scala 93:22:@58796.4]
  wire  RetimeWrapper_562_io_out; // @[package.scala 93:22:@58796.4]
  wire  RetimeWrapper_563_clock; // @[package.scala 93:22:@58804.4]
  wire  RetimeWrapper_563_reset; // @[package.scala 93:22:@58804.4]
  wire  RetimeWrapper_563_io_flow; // @[package.scala 93:22:@58804.4]
  wire  RetimeWrapper_563_io_in; // @[package.scala 93:22:@58804.4]
  wire  RetimeWrapper_563_io_out; // @[package.scala 93:22:@58804.4]
  wire  RetimeWrapper_564_clock; // @[package.scala 93:22:@58812.4]
  wire  RetimeWrapper_564_reset; // @[package.scala 93:22:@58812.4]
  wire  RetimeWrapper_564_io_flow; // @[package.scala 93:22:@58812.4]
  wire  RetimeWrapper_564_io_in; // @[package.scala 93:22:@58812.4]
  wire  RetimeWrapper_564_io_out; // @[package.scala 93:22:@58812.4]
  wire  RetimeWrapper_565_clock; // @[package.scala 93:22:@58820.4]
  wire  RetimeWrapper_565_reset; // @[package.scala 93:22:@58820.4]
  wire  RetimeWrapper_565_io_flow; // @[package.scala 93:22:@58820.4]
  wire  RetimeWrapper_565_io_in; // @[package.scala 93:22:@58820.4]
  wire  RetimeWrapper_565_io_out; // @[package.scala 93:22:@58820.4]
  wire  RetimeWrapper_566_clock; // @[package.scala 93:22:@58828.4]
  wire  RetimeWrapper_566_reset; // @[package.scala 93:22:@58828.4]
  wire  RetimeWrapper_566_io_flow; // @[package.scala 93:22:@58828.4]
  wire  RetimeWrapper_566_io_in; // @[package.scala 93:22:@58828.4]
  wire  RetimeWrapper_566_io_out; // @[package.scala 93:22:@58828.4]
  wire  RetimeWrapper_567_clock; // @[package.scala 93:22:@58836.4]
  wire  RetimeWrapper_567_reset; // @[package.scala 93:22:@58836.4]
  wire  RetimeWrapper_567_io_flow; // @[package.scala 93:22:@58836.4]
  wire  RetimeWrapper_567_io_in; // @[package.scala 93:22:@58836.4]
  wire  RetimeWrapper_567_io_out; // @[package.scala 93:22:@58836.4]
  wire  RetimeWrapper_568_clock; // @[package.scala 93:22:@58844.4]
  wire  RetimeWrapper_568_reset; // @[package.scala 93:22:@58844.4]
  wire  RetimeWrapper_568_io_flow; // @[package.scala 93:22:@58844.4]
  wire  RetimeWrapper_568_io_in; // @[package.scala 93:22:@58844.4]
  wire  RetimeWrapper_568_io_out; // @[package.scala 93:22:@58844.4]
  wire  RetimeWrapper_569_clock; // @[package.scala 93:22:@58852.4]
  wire  RetimeWrapper_569_reset; // @[package.scala 93:22:@58852.4]
  wire  RetimeWrapper_569_io_flow; // @[package.scala 93:22:@58852.4]
  wire  RetimeWrapper_569_io_in; // @[package.scala 93:22:@58852.4]
  wire  RetimeWrapper_569_io_out; // @[package.scala 93:22:@58852.4]
  wire  RetimeWrapper_570_clock; // @[package.scala 93:22:@58860.4]
  wire  RetimeWrapper_570_reset; // @[package.scala 93:22:@58860.4]
  wire  RetimeWrapper_570_io_flow; // @[package.scala 93:22:@58860.4]
  wire  RetimeWrapper_570_io_in; // @[package.scala 93:22:@58860.4]
  wire  RetimeWrapper_570_io_out; // @[package.scala 93:22:@58860.4]
  wire  RetimeWrapper_571_clock; // @[package.scala 93:22:@58868.4]
  wire  RetimeWrapper_571_reset; // @[package.scala 93:22:@58868.4]
  wire  RetimeWrapper_571_io_flow; // @[package.scala 93:22:@58868.4]
  wire  RetimeWrapper_571_io_in; // @[package.scala 93:22:@58868.4]
  wire  RetimeWrapper_571_io_out; // @[package.scala 93:22:@58868.4]
  wire  RetimeWrapper_572_clock; // @[package.scala 93:22:@58876.4]
  wire  RetimeWrapper_572_reset; // @[package.scala 93:22:@58876.4]
  wire  RetimeWrapper_572_io_flow; // @[package.scala 93:22:@58876.4]
  wire  RetimeWrapper_572_io_in; // @[package.scala 93:22:@58876.4]
  wire  RetimeWrapper_572_io_out; // @[package.scala 93:22:@58876.4]
  wire  RetimeWrapper_573_clock; // @[package.scala 93:22:@58884.4]
  wire  RetimeWrapper_573_reset; // @[package.scala 93:22:@58884.4]
  wire  RetimeWrapper_573_io_flow; // @[package.scala 93:22:@58884.4]
  wire  RetimeWrapper_573_io_in; // @[package.scala 93:22:@58884.4]
  wire  RetimeWrapper_573_io_out; // @[package.scala 93:22:@58884.4]
  wire  RetimeWrapper_574_clock; // @[package.scala 93:22:@58892.4]
  wire  RetimeWrapper_574_reset; // @[package.scala 93:22:@58892.4]
  wire  RetimeWrapper_574_io_flow; // @[package.scala 93:22:@58892.4]
  wire  RetimeWrapper_574_io_in; // @[package.scala 93:22:@58892.4]
  wire  RetimeWrapper_574_io_out; // @[package.scala 93:22:@58892.4]
  wire  RetimeWrapper_575_clock; // @[package.scala 93:22:@58900.4]
  wire  RetimeWrapper_575_reset; // @[package.scala 93:22:@58900.4]
  wire  RetimeWrapper_575_io_flow; // @[package.scala 93:22:@58900.4]
  wire  RetimeWrapper_575_io_in; // @[package.scala 93:22:@58900.4]
  wire  RetimeWrapper_575_io_out; // @[package.scala 93:22:@58900.4]
  wire  RetimeWrapper_576_clock; // @[package.scala 93:22:@58908.4]
  wire  RetimeWrapper_576_reset; // @[package.scala 93:22:@58908.4]
  wire  RetimeWrapper_576_io_flow; // @[package.scala 93:22:@58908.4]
  wire  RetimeWrapper_576_io_in; // @[package.scala 93:22:@58908.4]
  wire  RetimeWrapper_576_io_out; // @[package.scala 93:22:@58908.4]
  wire  RetimeWrapper_577_clock; // @[package.scala 93:22:@58916.4]
  wire  RetimeWrapper_577_reset; // @[package.scala 93:22:@58916.4]
  wire  RetimeWrapper_577_io_flow; // @[package.scala 93:22:@58916.4]
  wire  RetimeWrapper_577_io_in; // @[package.scala 93:22:@58916.4]
  wire  RetimeWrapper_577_io_out; // @[package.scala 93:22:@58916.4]
  wire  RetimeWrapper_578_clock; // @[package.scala 93:22:@58924.4]
  wire  RetimeWrapper_578_reset; // @[package.scala 93:22:@58924.4]
  wire  RetimeWrapper_578_io_flow; // @[package.scala 93:22:@58924.4]
  wire  RetimeWrapper_578_io_in; // @[package.scala 93:22:@58924.4]
  wire  RetimeWrapper_578_io_out; // @[package.scala 93:22:@58924.4]
  wire  RetimeWrapper_579_clock; // @[package.scala 93:22:@58932.4]
  wire  RetimeWrapper_579_reset; // @[package.scala 93:22:@58932.4]
  wire  RetimeWrapper_579_io_flow; // @[package.scala 93:22:@58932.4]
  wire  RetimeWrapper_579_io_in; // @[package.scala 93:22:@58932.4]
  wire  RetimeWrapper_579_io_out; // @[package.scala 93:22:@58932.4]
  wire  RetimeWrapper_580_clock; // @[package.scala 93:22:@59020.4]
  wire  RetimeWrapper_580_reset; // @[package.scala 93:22:@59020.4]
  wire  RetimeWrapper_580_io_flow; // @[package.scala 93:22:@59020.4]
  wire  RetimeWrapper_580_io_in; // @[package.scala 93:22:@59020.4]
  wire  RetimeWrapper_580_io_out; // @[package.scala 93:22:@59020.4]
  wire  RetimeWrapper_581_clock; // @[package.scala 93:22:@59028.4]
  wire  RetimeWrapper_581_reset; // @[package.scala 93:22:@59028.4]
  wire  RetimeWrapper_581_io_flow; // @[package.scala 93:22:@59028.4]
  wire  RetimeWrapper_581_io_in; // @[package.scala 93:22:@59028.4]
  wire  RetimeWrapper_581_io_out; // @[package.scala 93:22:@59028.4]
  wire  RetimeWrapper_582_clock; // @[package.scala 93:22:@59036.4]
  wire  RetimeWrapper_582_reset; // @[package.scala 93:22:@59036.4]
  wire  RetimeWrapper_582_io_flow; // @[package.scala 93:22:@59036.4]
  wire  RetimeWrapper_582_io_in; // @[package.scala 93:22:@59036.4]
  wire  RetimeWrapper_582_io_out; // @[package.scala 93:22:@59036.4]
  wire  RetimeWrapper_583_clock; // @[package.scala 93:22:@59044.4]
  wire  RetimeWrapper_583_reset; // @[package.scala 93:22:@59044.4]
  wire  RetimeWrapper_583_io_flow; // @[package.scala 93:22:@59044.4]
  wire  RetimeWrapper_583_io_in; // @[package.scala 93:22:@59044.4]
  wire  RetimeWrapper_583_io_out; // @[package.scala 93:22:@59044.4]
  wire  RetimeWrapper_584_clock; // @[package.scala 93:22:@59052.4]
  wire  RetimeWrapper_584_reset; // @[package.scala 93:22:@59052.4]
  wire  RetimeWrapper_584_io_flow; // @[package.scala 93:22:@59052.4]
  wire  RetimeWrapper_584_io_in; // @[package.scala 93:22:@59052.4]
  wire  RetimeWrapper_584_io_out; // @[package.scala 93:22:@59052.4]
  wire  RetimeWrapper_585_clock; // @[package.scala 93:22:@59060.4]
  wire  RetimeWrapper_585_reset; // @[package.scala 93:22:@59060.4]
  wire  RetimeWrapper_585_io_flow; // @[package.scala 93:22:@59060.4]
  wire  RetimeWrapper_585_io_in; // @[package.scala 93:22:@59060.4]
  wire  RetimeWrapper_585_io_out; // @[package.scala 93:22:@59060.4]
  wire  RetimeWrapper_586_clock; // @[package.scala 93:22:@59068.4]
  wire  RetimeWrapper_586_reset; // @[package.scala 93:22:@59068.4]
  wire  RetimeWrapper_586_io_flow; // @[package.scala 93:22:@59068.4]
  wire  RetimeWrapper_586_io_in; // @[package.scala 93:22:@59068.4]
  wire  RetimeWrapper_586_io_out; // @[package.scala 93:22:@59068.4]
  wire  RetimeWrapper_587_clock; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_587_reset; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_587_io_flow; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_587_io_in; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_587_io_out; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_588_clock; // @[package.scala 93:22:@59084.4]
  wire  RetimeWrapper_588_reset; // @[package.scala 93:22:@59084.4]
  wire  RetimeWrapper_588_io_flow; // @[package.scala 93:22:@59084.4]
  wire  RetimeWrapper_588_io_in; // @[package.scala 93:22:@59084.4]
  wire  RetimeWrapper_588_io_out; // @[package.scala 93:22:@59084.4]
  wire  RetimeWrapper_589_clock; // @[package.scala 93:22:@59092.4]
  wire  RetimeWrapper_589_reset; // @[package.scala 93:22:@59092.4]
  wire  RetimeWrapper_589_io_flow; // @[package.scala 93:22:@59092.4]
  wire  RetimeWrapper_589_io_in; // @[package.scala 93:22:@59092.4]
  wire  RetimeWrapper_589_io_out; // @[package.scala 93:22:@59092.4]
  wire  RetimeWrapper_590_clock; // @[package.scala 93:22:@59100.4]
  wire  RetimeWrapper_590_reset; // @[package.scala 93:22:@59100.4]
  wire  RetimeWrapper_590_io_flow; // @[package.scala 93:22:@59100.4]
  wire  RetimeWrapper_590_io_in; // @[package.scala 93:22:@59100.4]
  wire  RetimeWrapper_590_io_out; // @[package.scala 93:22:@59100.4]
  wire  RetimeWrapper_591_clock; // @[package.scala 93:22:@59108.4]
  wire  RetimeWrapper_591_reset; // @[package.scala 93:22:@59108.4]
  wire  RetimeWrapper_591_io_flow; // @[package.scala 93:22:@59108.4]
  wire  RetimeWrapper_591_io_in; // @[package.scala 93:22:@59108.4]
  wire  RetimeWrapper_591_io_out; // @[package.scala 93:22:@59108.4]
  wire  RetimeWrapper_592_clock; // @[package.scala 93:22:@59116.4]
  wire  RetimeWrapper_592_reset; // @[package.scala 93:22:@59116.4]
  wire  RetimeWrapper_592_io_flow; // @[package.scala 93:22:@59116.4]
  wire  RetimeWrapper_592_io_in; // @[package.scala 93:22:@59116.4]
  wire  RetimeWrapper_592_io_out; // @[package.scala 93:22:@59116.4]
  wire  RetimeWrapper_593_clock; // @[package.scala 93:22:@59124.4]
  wire  RetimeWrapper_593_reset; // @[package.scala 93:22:@59124.4]
  wire  RetimeWrapper_593_io_flow; // @[package.scala 93:22:@59124.4]
  wire  RetimeWrapper_593_io_in; // @[package.scala 93:22:@59124.4]
  wire  RetimeWrapper_593_io_out; // @[package.scala 93:22:@59124.4]
  wire  RetimeWrapper_594_clock; // @[package.scala 93:22:@59132.4]
  wire  RetimeWrapper_594_reset; // @[package.scala 93:22:@59132.4]
  wire  RetimeWrapper_594_io_flow; // @[package.scala 93:22:@59132.4]
  wire  RetimeWrapper_594_io_in; // @[package.scala 93:22:@59132.4]
  wire  RetimeWrapper_594_io_out; // @[package.scala 93:22:@59132.4]
  wire  RetimeWrapper_595_clock; // @[package.scala 93:22:@59140.4]
  wire  RetimeWrapper_595_reset; // @[package.scala 93:22:@59140.4]
  wire  RetimeWrapper_595_io_flow; // @[package.scala 93:22:@59140.4]
  wire  RetimeWrapper_595_io_in; // @[package.scala 93:22:@59140.4]
  wire  RetimeWrapper_595_io_out; // @[package.scala 93:22:@59140.4]
  wire  RetimeWrapper_596_clock; // @[package.scala 93:22:@59148.4]
  wire  RetimeWrapper_596_reset; // @[package.scala 93:22:@59148.4]
  wire  RetimeWrapper_596_io_flow; // @[package.scala 93:22:@59148.4]
  wire  RetimeWrapper_596_io_in; // @[package.scala 93:22:@59148.4]
  wire  RetimeWrapper_596_io_out; // @[package.scala 93:22:@59148.4]
  wire  RetimeWrapper_597_clock; // @[package.scala 93:22:@59156.4]
  wire  RetimeWrapper_597_reset; // @[package.scala 93:22:@59156.4]
  wire  RetimeWrapper_597_io_flow; // @[package.scala 93:22:@59156.4]
  wire  RetimeWrapper_597_io_in; // @[package.scala 93:22:@59156.4]
  wire  RetimeWrapper_597_io_out; // @[package.scala 93:22:@59156.4]
  wire  RetimeWrapper_598_clock; // @[package.scala 93:22:@59164.4]
  wire  RetimeWrapper_598_reset; // @[package.scala 93:22:@59164.4]
  wire  RetimeWrapper_598_io_flow; // @[package.scala 93:22:@59164.4]
  wire  RetimeWrapper_598_io_in; // @[package.scala 93:22:@59164.4]
  wire  RetimeWrapper_598_io_out; // @[package.scala 93:22:@59164.4]
  wire  RetimeWrapper_599_clock; // @[package.scala 93:22:@59172.4]
  wire  RetimeWrapper_599_reset; // @[package.scala 93:22:@59172.4]
  wire  RetimeWrapper_599_io_flow; // @[package.scala 93:22:@59172.4]
  wire  RetimeWrapper_599_io_in; // @[package.scala 93:22:@59172.4]
  wire  RetimeWrapper_599_io_out; // @[package.scala 93:22:@59172.4]
  wire  _T_1212; // @[MemPrimitives.scala 82:210:@44959.4]
  wire  _T_1214; // @[MemPrimitives.scala 82:210:@44960.4]
  wire  _T_1215; // @[MemPrimitives.scala 82:228:@44961.4]
  wire  _T_1216; // @[MemPrimitives.scala 83:102:@44962.4]
  wire  _T_1218; // @[MemPrimitives.scala 82:210:@44963.4]
  wire  _T_1220; // @[MemPrimitives.scala 82:210:@44964.4]
  wire  _T_1221; // @[MemPrimitives.scala 82:228:@44965.4]
  wire  _T_1222; // @[MemPrimitives.scala 83:102:@44966.4]
  wire  _T_1224; // @[MemPrimitives.scala 82:210:@44967.4]
  wire  _T_1226; // @[MemPrimitives.scala 82:210:@44968.4]
  wire  _T_1227; // @[MemPrimitives.scala 82:228:@44969.4]
  wire  _T_1228; // @[MemPrimitives.scala 83:102:@44970.4]
  wire  _T_1230; // @[MemPrimitives.scala 82:210:@44971.4]
  wire  _T_1232; // @[MemPrimitives.scala 82:210:@44972.4]
  wire  _T_1233; // @[MemPrimitives.scala 82:228:@44973.4]
  wire  _T_1234; // @[MemPrimitives.scala 83:102:@44974.4]
  wire [16:0] _T_1236; // @[Cat.scala 30:58:@44976.4]
  wire [16:0] _T_1238; // @[Cat.scala 30:58:@44978.4]
  wire [16:0] _T_1240; // @[Cat.scala 30:58:@44980.4]
  wire [16:0] _T_1242; // @[Cat.scala 30:58:@44982.4]
  wire [16:0] _T_1243; // @[Mux.scala 31:69:@44983.4]
  wire [16:0] _T_1244; // @[Mux.scala 31:69:@44984.4]
  wire [16:0] _T_1245; // @[Mux.scala 31:69:@44985.4]
  wire  _T_1250; // @[MemPrimitives.scala 82:210:@44992.4]
  wire  _T_1252; // @[MemPrimitives.scala 82:210:@44993.4]
  wire  _T_1253; // @[MemPrimitives.scala 82:228:@44994.4]
  wire  _T_1254; // @[MemPrimitives.scala 83:102:@44995.4]
  wire  _T_1256; // @[MemPrimitives.scala 82:210:@44996.4]
  wire  _T_1258; // @[MemPrimitives.scala 82:210:@44997.4]
  wire  _T_1259; // @[MemPrimitives.scala 82:228:@44998.4]
  wire  _T_1260; // @[MemPrimitives.scala 83:102:@44999.4]
  wire  _T_1262; // @[MemPrimitives.scala 82:210:@45000.4]
  wire  _T_1264; // @[MemPrimitives.scala 82:210:@45001.4]
  wire  _T_1265; // @[MemPrimitives.scala 82:228:@45002.4]
  wire  _T_1266; // @[MemPrimitives.scala 83:102:@45003.4]
  wire  _T_1268; // @[MemPrimitives.scala 82:210:@45004.4]
  wire  _T_1270; // @[MemPrimitives.scala 82:210:@45005.4]
  wire  _T_1271; // @[MemPrimitives.scala 82:228:@45006.4]
  wire  _T_1272; // @[MemPrimitives.scala 83:102:@45007.4]
  wire [16:0] _T_1274; // @[Cat.scala 30:58:@45009.4]
  wire [16:0] _T_1276; // @[Cat.scala 30:58:@45011.4]
  wire [16:0] _T_1278; // @[Cat.scala 30:58:@45013.4]
  wire [16:0] _T_1280; // @[Cat.scala 30:58:@45015.4]
  wire [16:0] _T_1281; // @[Mux.scala 31:69:@45016.4]
  wire [16:0] _T_1282; // @[Mux.scala 31:69:@45017.4]
  wire [16:0] _T_1283; // @[Mux.scala 31:69:@45018.4]
  wire  _T_1290; // @[MemPrimitives.scala 82:210:@45026.4]
  wire  _T_1291; // @[MemPrimitives.scala 82:228:@45027.4]
  wire  _T_1292; // @[MemPrimitives.scala 83:102:@45028.4]
  wire  _T_1296; // @[MemPrimitives.scala 82:210:@45030.4]
  wire  _T_1297; // @[MemPrimitives.scala 82:228:@45031.4]
  wire  _T_1298; // @[MemPrimitives.scala 83:102:@45032.4]
  wire  _T_1302; // @[MemPrimitives.scala 82:210:@45034.4]
  wire  _T_1303; // @[MemPrimitives.scala 82:228:@45035.4]
  wire  _T_1304; // @[MemPrimitives.scala 83:102:@45036.4]
  wire  _T_1308; // @[MemPrimitives.scala 82:210:@45038.4]
  wire  _T_1309; // @[MemPrimitives.scala 82:228:@45039.4]
  wire  _T_1310; // @[MemPrimitives.scala 83:102:@45040.4]
  wire [16:0] _T_1312; // @[Cat.scala 30:58:@45042.4]
  wire [16:0] _T_1314; // @[Cat.scala 30:58:@45044.4]
  wire [16:0] _T_1316; // @[Cat.scala 30:58:@45046.4]
  wire [16:0] _T_1318; // @[Cat.scala 30:58:@45048.4]
  wire [16:0] _T_1319; // @[Mux.scala 31:69:@45049.4]
  wire [16:0] _T_1320; // @[Mux.scala 31:69:@45050.4]
  wire [16:0] _T_1321; // @[Mux.scala 31:69:@45051.4]
  wire  _T_1328; // @[MemPrimitives.scala 82:210:@45059.4]
  wire  _T_1329; // @[MemPrimitives.scala 82:228:@45060.4]
  wire  _T_1330; // @[MemPrimitives.scala 83:102:@45061.4]
  wire  _T_1334; // @[MemPrimitives.scala 82:210:@45063.4]
  wire  _T_1335; // @[MemPrimitives.scala 82:228:@45064.4]
  wire  _T_1336; // @[MemPrimitives.scala 83:102:@45065.4]
  wire  _T_1340; // @[MemPrimitives.scala 82:210:@45067.4]
  wire  _T_1341; // @[MemPrimitives.scala 82:228:@45068.4]
  wire  _T_1342; // @[MemPrimitives.scala 83:102:@45069.4]
  wire  _T_1346; // @[MemPrimitives.scala 82:210:@45071.4]
  wire  _T_1347; // @[MemPrimitives.scala 82:228:@45072.4]
  wire  _T_1348; // @[MemPrimitives.scala 83:102:@45073.4]
  wire [16:0] _T_1350; // @[Cat.scala 30:58:@45075.4]
  wire [16:0] _T_1352; // @[Cat.scala 30:58:@45077.4]
  wire [16:0] _T_1354; // @[Cat.scala 30:58:@45079.4]
  wire [16:0] _T_1356; // @[Cat.scala 30:58:@45081.4]
  wire [16:0] _T_1357; // @[Mux.scala 31:69:@45082.4]
  wire [16:0] _T_1358; // @[Mux.scala 31:69:@45083.4]
  wire [16:0] _T_1359; // @[Mux.scala 31:69:@45084.4]
  wire  _T_1366; // @[MemPrimitives.scala 82:210:@45092.4]
  wire  _T_1367; // @[MemPrimitives.scala 82:228:@45093.4]
  wire  _T_1368; // @[MemPrimitives.scala 83:102:@45094.4]
  wire  _T_1372; // @[MemPrimitives.scala 82:210:@45096.4]
  wire  _T_1373; // @[MemPrimitives.scala 82:228:@45097.4]
  wire  _T_1374; // @[MemPrimitives.scala 83:102:@45098.4]
  wire  _T_1378; // @[MemPrimitives.scala 82:210:@45100.4]
  wire  _T_1379; // @[MemPrimitives.scala 82:228:@45101.4]
  wire  _T_1380; // @[MemPrimitives.scala 83:102:@45102.4]
  wire  _T_1384; // @[MemPrimitives.scala 82:210:@45104.4]
  wire  _T_1385; // @[MemPrimitives.scala 82:228:@45105.4]
  wire  _T_1386; // @[MemPrimitives.scala 83:102:@45106.4]
  wire [16:0] _T_1388; // @[Cat.scala 30:58:@45108.4]
  wire [16:0] _T_1390; // @[Cat.scala 30:58:@45110.4]
  wire [16:0] _T_1392; // @[Cat.scala 30:58:@45112.4]
  wire [16:0] _T_1394; // @[Cat.scala 30:58:@45114.4]
  wire [16:0] _T_1395; // @[Mux.scala 31:69:@45115.4]
  wire [16:0] _T_1396; // @[Mux.scala 31:69:@45116.4]
  wire [16:0] _T_1397; // @[Mux.scala 31:69:@45117.4]
  wire  _T_1404; // @[MemPrimitives.scala 82:210:@45125.4]
  wire  _T_1405; // @[MemPrimitives.scala 82:228:@45126.4]
  wire  _T_1406; // @[MemPrimitives.scala 83:102:@45127.4]
  wire  _T_1410; // @[MemPrimitives.scala 82:210:@45129.4]
  wire  _T_1411; // @[MemPrimitives.scala 82:228:@45130.4]
  wire  _T_1412; // @[MemPrimitives.scala 83:102:@45131.4]
  wire  _T_1416; // @[MemPrimitives.scala 82:210:@45133.4]
  wire  _T_1417; // @[MemPrimitives.scala 82:228:@45134.4]
  wire  _T_1418; // @[MemPrimitives.scala 83:102:@45135.4]
  wire  _T_1422; // @[MemPrimitives.scala 82:210:@45137.4]
  wire  _T_1423; // @[MemPrimitives.scala 82:228:@45138.4]
  wire  _T_1424; // @[MemPrimitives.scala 83:102:@45139.4]
  wire [16:0] _T_1426; // @[Cat.scala 30:58:@45141.4]
  wire [16:0] _T_1428; // @[Cat.scala 30:58:@45143.4]
  wire [16:0] _T_1430; // @[Cat.scala 30:58:@45145.4]
  wire [16:0] _T_1432; // @[Cat.scala 30:58:@45147.4]
  wire [16:0] _T_1433; // @[Mux.scala 31:69:@45148.4]
  wire [16:0] _T_1434; // @[Mux.scala 31:69:@45149.4]
  wire [16:0] _T_1435; // @[Mux.scala 31:69:@45150.4]
  wire  _T_1442; // @[MemPrimitives.scala 82:210:@45158.4]
  wire  _T_1443; // @[MemPrimitives.scala 82:228:@45159.4]
  wire  _T_1444; // @[MemPrimitives.scala 83:102:@45160.4]
  wire  _T_1448; // @[MemPrimitives.scala 82:210:@45162.4]
  wire  _T_1449; // @[MemPrimitives.scala 82:228:@45163.4]
  wire  _T_1450; // @[MemPrimitives.scala 83:102:@45164.4]
  wire  _T_1454; // @[MemPrimitives.scala 82:210:@45166.4]
  wire  _T_1455; // @[MemPrimitives.scala 82:228:@45167.4]
  wire  _T_1456; // @[MemPrimitives.scala 83:102:@45168.4]
  wire  _T_1460; // @[MemPrimitives.scala 82:210:@45170.4]
  wire  _T_1461; // @[MemPrimitives.scala 82:228:@45171.4]
  wire  _T_1462; // @[MemPrimitives.scala 83:102:@45172.4]
  wire [16:0] _T_1464; // @[Cat.scala 30:58:@45174.4]
  wire [16:0] _T_1466; // @[Cat.scala 30:58:@45176.4]
  wire [16:0] _T_1468; // @[Cat.scala 30:58:@45178.4]
  wire [16:0] _T_1470; // @[Cat.scala 30:58:@45180.4]
  wire [16:0] _T_1471; // @[Mux.scala 31:69:@45181.4]
  wire [16:0] _T_1472; // @[Mux.scala 31:69:@45182.4]
  wire [16:0] _T_1473; // @[Mux.scala 31:69:@45183.4]
  wire  _T_1480; // @[MemPrimitives.scala 82:210:@45191.4]
  wire  _T_1481; // @[MemPrimitives.scala 82:228:@45192.4]
  wire  _T_1482; // @[MemPrimitives.scala 83:102:@45193.4]
  wire  _T_1486; // @[MemPrimitives.scala 82:210:@45195.4]
  wire  _T_1487; // @[MemPrimitives.scala 82:228:@45196.4]
  wire  _T_1488; // @[MemPrimitives.scala 83:102:@45197.4]
  wire  _T_1492; // @[MemPrimitives.scala 82:210:@45199.4]
  wire  _T_1493; // @[MemPrimitives.scala 82:228:@45200.4]
  wire  _T_1494; // @[MemPrimitives.scala 83:102:@45201.4]
  wire  _T_1498; // @[MemPrimitives.scala 82:210:@45203.4]
  wire  _T_1499; // @[MemPrimitives.scala 82:228:@45204.4]
  wire  _T_1500; // @[MemPrimitives.scala 83:102:@45205.4]
  wire [16:0] _T_1502; // @[Cat.scala 30:58:@45207.4]
  wire [16:0] _T_1504; // @[Cat.scala 30:58:@45209.4]
  wire [16:0] _T_1506; // @[Cat.scala 30:58:@45211.4]
  wire [16:0] _T_1508; // @[Cat.scala 30:58:@45213.4]
  wire [16:0] _T_1509; // @[Mux.scala 31:69:@45214.4]
  wire [16:0] _T_1510; // @[Mux.scala 31:69:@45215.4]
  wire [16:0] _T_1511; // @[Mux.scala 31:69:@45216.4]
  wire  _T_1518; // @[MemPrimitives.scala 82:210:@45224.4]
  wire  _T_1519; // @[MemPrimitives.scala 82:228:@45225.4]
  wire  _T_1520; // @[MemPrimitives.scala 83:102:@45226.4]
  wire  _T_1524; // @[MemPrimitives.scala 82:210:@45228.4]
  wire  _T_1525; // @[MemPrimitives.scala 82:228:@45229.4]
  wire  _T_1526; // @[MemPrimitives.scala 83:102:@45230.4]
  wire  _T_1530; // @[MemPrimitives.scala 82:210:@45232.4]
  wire  _T_1531; // @[MemPrimitives.scala 82:228:@45233.4]
  wire  _T_1532; // @[MemPrimitives.scala 83:102:@45234.4]
  wire  _T_1536; // @[MemPrimitives.scala 82:210:@45236.4]
  wire  _T_1537; // @[MemPrimitives.scala 82:228:@45237.4]
  wire  _T_1538; // @[MemPrimitives.scala 83:102:@45238.4]
  wire [16:0] _T_1540; // @[Cat.scala 30:58:@45240.4]
  wire [16:0] _T_1542; // @[Cat.scala 30:58:@45242.4]
  wire [16:0] _T_1544; // @[Cat.scala 30:58:@45244.4]
  wire [16:0] _T_1546; // @[Cat.scala 30:58:@45246.4]
  wire [16:0] _T_1547; // @[Mux.scala 31:69:@45247.4]
  wire [16:0] _T_1548; // @[Mux.scala 31:69:@45248.4]
  wire [16:0] _T_1549; // @[Mux.scala 31:69:@45249.4]
  wire  _T_1556; // @[MemPrimitives.scala 82:210:@45257.4]
  wire  _T_1557; // @[MemPrimitives.scala 82:228:@45258.4]
  wire  _T_1558; // @[MemPrimitives.scala 83:102:@45259.4]
  wire  _T_1562; // @[MemPrimitives.scala 82:210:@45261.4]
  wire  _T_1563; // @[MemPrimitives.scala 82:228:@45262.4]
  wire  _T_1564; // @[MemPrimitives.scala 83:102:@45263.4]
  wire  _T_1568; // @[MemPrimitives.scala 82:210:@45265.4]
  wire  _T_1569; // @[MemPrimitives.scala 82:228:@45266.4]
  wire  _T_1570; // @[MemPrimitives.scala 83:102:@45267.4]
  wire  _T_1574; // @[MemPrimitives.scala 82:210:@45269.4]
  wire  _T_1575; // @[MemPrimitives.scala 82:228:@45270.4]
  wire  _T_1576; // @[MemPrimitives.scala 83:102:@45271.4]
  wire [16:0] _T_1578; // @[Cat.scala 30:58:@45273.4]
  wire [16:0] _T_1580; // @[Cat.scala 30:58:@45275.4]
  wire [16:0] _T_1582; // @[Cat.scala 30:58:@45277.4]
  wire [16:0] _T_1584; // @[Cat.scala 30:58:@45279.4]
  wire [16:0] _T_1585; // @[Mux.scala 31:69:@45280.4]
  wire [16:0] _T_1586; // @[Mux.scala 31:69:@45281.4]
  wire [16:0] _T_1587; // @[Mux.scala 31:69:@45282.4]
  wire  _T_1592; // @[MemPrimitives.scala 82:210:@45289.4]
  wire  _T_1595; // @[MemPrimitives.scala 82:228:@45291.4]
  wire  _T_1596; // @[MemPrimitives.scala 83:102:@45292.4]
  wire  _T_1598; // @[MemPrimitives.scala 82:210:@45293.4]
  wire  _T_1601; // @[MemPrimitives.scala 82:228:@45295.4]
  wire  _T_1602; // @[MemPrimitives.scala 83:102:@45296.4]
  wire  _T_1604; // @[MemPrimitives.scala 82:210:@45297.4]
  wire  _T_1607; // @[MemPrimitives.scala 82:228:@45299.4]
  wire  _T_1608; // @[MemPrimitives.scala 83:102:@45300.4]
  wire  _T_1610; // @[MemPrimitives.scala 82:210:@45301.4]
  wire  _T_1613; // @[MemPrimitives.scala 82:228:@45303.4]
  wire  _T_1614; // @[MemPrimitives.scala 83:102:@45304.4]
  wire [16:0] _T_1616; // @[Cat.scala 30:58:@45306.4]
  wire [16:0] _T_1618; // @[Cat.scala 30:58:@45308.4]
  wire [16:0] _T_1620; // @[Cat.scala 30:58:@45310.4]
  wire [16:0] _T_1622; // @[Cat.scala 30:58:@45312.4]
  wire [16:0] _T_1623; // @[Mux.scala 31:69:@45313.4]
  wire [16:0] _T_1624; // @[Mux.scala 31:69:@45314.4]
  wire [16:0] _T_1625; // @[Mux.scala 31:69:@45315.4]
  wire  _T_1630; // @[MemPrimitives.scala 82:210:@45322.4]
  wire  _T_1633; // @[MemPrimitives.scala 82:228:@45324.4]
  wire  _T_1634; // @[MemPrimitives.scala 83:102:@45325.4]
  wire  _T_1636; // @[MemPrimitives.scala 82:210:@45326.4]
  wire  _T_1639; // @[MemPrimitives.scala 82:228:@45328.4]
  wire  _T_1640; // @[MemPrimitives.scala 83:102:@45329.4]
  wire  _T_1642; // @[MemPrimitives.scala 82:210:@45330.4]
  wire  _T_1645; // @[MemPrimitives.scala 82:228:@45332.4]
  wire  _T_1646; // @[MemPrimitives.scala 83:102:@45333.4]
  wire  _T_1648; // @[MemPrimitives.scala 82:210:@45334.4]
  wire  _T_1651; // @[MemPrimitives.scala 82:228:@45336.4]
  wire  _T_1652; // @[MemPrimitives.scala 83:102:@45337.4]
  wire [16:0] _T_1654; // @[Cat.scala 30:58:@45339.4]
  wire [16:0] _T_1656; // @[Cat.scala 30:58:@45341.4]
  wire [16:0] _T_1658; // @[Cat.scala 30:58:@45343.4]
  wire [16:0] _T_1660; // @[Cat.scala 30:58:@45345.4]
  wire [16:0] _T_1661; // @[Mux.scala 31:69:@45346.4]
  wire [16:0] _T_1662; // @[Mux.scala 31:69:@45347.4]
  wire [16:0] _T_1663; // @[Mux.scala 31:69:@45348.4]
  wire  _T_1671; // @[MemPrimitives.scala 82:228:@45357.4]
  wire  _T_1672; // @[MemPrimitives.scala 83:102:@45358.4]
  wire  _T_1677; // @[MemPrimitives.scala 82:228:@45361.4]
  wire  _T_1678; // @[MemPrimitives.scala 83:102:@45362.4]
  wire  _T_1683; // @[MemPrimitives.scala 82:228:@45365.4]
  wire  _T_1684; // @[MemPrimitives.scala 83:102:@45366.4]
  wire  _T_1689; // @[MemPrimitives.scala 82:228:@45369.4]
  wire  _T_1690; // @[MemPrimitives.scala 83:102:@45370.4]
  wire [16:0] _T_1692; // @[Cat.scala 30:58:@45372.4]
  wire [16:0] _T_1694; // @[Cat.scala 30:58:@45374.4]
  wire [16:0] _T_1696; // @[Cat.scala 30:58:@45376.4]
  wire [16:0] _T_1698; // @[Cat.scala 30:58:@45378.4]
  wire [16:0] _T_1699; // @[Mux.scala 31:69:@45379.4]
  wire [16:0] _T_1700; // @[Mux.scala 31:69:@45380.4]
  wire [16:0] _T_1701; // @[Mux.scala 31:69:@45381.4]
  wire  _T_1709; // @[MemPrimitives.scala 82:228:@45390.4]
  wire  _T_1710; // @[MemPrimitives.scala 83:102:@45391.4]
  wire  _T_1715; // @[MemPrimitives.scala 82:228:@45394.4]
  wire  _T_1716; // @[MemPrimitives.scala 83:102:@45395.4]
  wire  _T_1721; // @[MemPrimitives.scala 82:228:@45398.4]
  wire  _T_1722; // @[MemPrimitives.scala 83:102:@45399.4]
  wire  _T_1727; // @[MemPrimitives.scala 82:228:@45402.4]
  wire  _T_1728; // @[MemPrimitives.scala 83:102:@45403.4]
  wire [16:0] _T_1730; // @[Cat.scala 30:58:@45405.4]
  wire [16:0] _T_1732; // @[Cat.scala 30:58:@45407.4]
  wire [16:0] _T_1734; // @[Cat.scala 30:58:@45409.4]
  wire [16:0] _T_1736; // @[Cat.scala 30:58:@45411.4]
  wire [16:0] _T_1737; // @[Mux.scala 31:69:@45412.4]
  wire [16:0] _T_1738; // @[Mux.scala 31:69:@45413.4]
  wire [16:0] _T_1739; // @[Mux.scala 31:69:@45414.4]
  wire  _T_1747; // @[MemPrimitives.scala 82:228:@45423.4]
  wire  _T_1748; // @[MemPrimitives.scala 83:102:@45424.4]
  wire  _T_1753; // @[MemPrimitives.scala 82:228:@45427.4]
  wire  _T_1754; // @[MemPrimitives.scala 83:102:@45428.4]
  wire  _T_1759; // @[MemPrimitives.scala 82:228:@45431.4]
  wire  _T_1760; // @[MemPrimitives.scala 83:102:@45432.4]
  wire  _T_1765; // @[MemPrimitives.scala 82:228:@45435.4]
  wire  _T_1766; // @[MemPrimitives.scala 83:102:@45436.4]
  wire [16:0] _T_1768; // @[Cat.scala 30:58:@45438.4]
  wire [16:0] _T_1770; // @[Cat.scala 30:58:@45440.4]
  wire [16:0] _T_1772; // @[Cat.scala 30:58:@45442.4]
  wire [16:0] _T_1774; // @[Cat.scala 30:58:@45444.4]
  wire [16:0] _T_1775; // @[Mux.scala 31:69:@45445.4]
  wire [16:0] _T_1776; // @[Mux.scala 31:69:@45446.4]
  wire [16:0] _T_1777; // @[Mux.scala 31:69:@45447.4]
  wire  _T_1785; // @[MemPrimitives.scala 82:228:@45456.4]
  wire  _T_1786; // @[MemPrimitives.scala 83:102:@45457.4]
  wire  _T_1791; // @[MemPrimitives.scala 82:228:@45460.4]
  wire  _T_1792; // @[MemPrimitives.scala 83:102:@45461.4]
  wire  _T_1797; // @[MemPrimitives.scala 82:228:@45464.4]
  wire  _T_1798; // @[MemPrimitives.scala 83:102:@45465.4]
  wire  _T_1803; // @[MemPrimitives.scala 82:228:@45468.4]
  wire  _T_1804; // @[MemPrimitives.scala 83:102:@45469.4]
  wire [16:0] _T_1806; // @[Cat.scala 30:58:@45471.4]
  wire [16:0] _T_1808; // @[Cat.scala 30:58:@45473.4]
  wire [16:0] _T_1810; // @[Cat.scala 30:58:@45475.4]
  wire [16:0] _T_1812; // @[Cat.scala 30:58:@45477.4]
  wire [16:0] _T_1813; // @[Mux.scala 31:69:@45478.4]
  wire [16:0] _T_1814; // @[Mux.scala 31:69:@45479.4]
  wire [16:0] _T_1815; // @[Mux.scala 31:69:@45480.4]
  wire  _T_1823; // @[MemPrimitives.scala 82:228:@45489.4]
  wire  _T_1824; // @[MemPrimitives.scala 83:102:@45490.4]
  wire  _T_1829; // @[MemPrimitives.scala 82:228:@45493.4]
  wire  _T_1830; // @[MemPrimitives.scala 83:102:@45494.4]
  wire  _T_1835; // @[MemPrimitives.scala 82:228:@45497.4]
  wire  _T_1836; // @[MemPrimitives.scala 83:102:@45498.4]
  wire  _T_1841; // @[MemPrimitives.scala 82:228:@45501.4]
  wire  _T_1842; // @[MemPrimitives.scala 83:102:@45502.4]
  wire [16:0] _T_1844; // @[Cat.scala 30:58:@45504.4]
  wire [16:0] _T_1846; // @[Cat.scala 30:58:@45506.4]
  wire [16:0] _T_1848; // @[Cat.scala 30:58:@45508.4]
  wire [16:0] _T_1850; // @[Cat.scala 30:58:@45510.4]
  wire [16:0] _T_1851; // @[Mux.scala 31:69:@45511.4]
  wire [16:0] _T_1852; // @[Mux.scala 31:69:@45512.4]
  wire [16:0] _T_1853; // @[Mux.scala 31:69:@45513.4]
  wire  _T_1861; // @[MemPrimitives.scala 82:228:@45522.4]
  wire  _T_1862; // @[MemPrimitives.scala 83:102:@45523.4]
  wire  _T_1867; // @[MemPrimitives.scala 82:228:@45526.4]
  wire  _T_1868; // @[MemPrimitives.scala 83:102:@45527.4]
  wire  _T_1873; // @[MemPrimitives.scala 82:228:@45530.4]
  wire  _T_1874; // @[MemPrimitives.scala 83:102:@45531.4]
  wire  _T_1879; // @[MemPrimitives.scala 82:228:@45534.4]
  wire  _T_1880; // @[MemPrimitives.scala 83:102:@45535.4]
  wire [16:0] _T_1882; // @[Cat.scala 30:58:@45537.4]
  wire [16:0] _T_1884; // @[Cat.scala 30:58:@45539.4]
  wire [16:0] _T_1886; // @[Cat.scala 30:58:@45541.4]
  wire [16:0] _T_1888; // @[Cat.scala 30:58:@45543.4]
  wire [16:0] _T_1889; // @[Mux.scala 31:69:@45544.4]
  wire [16:0] _T_1890; // @[Mux.scala 31:69:@45545.4]
  wire [16:0] _T_1891; // @[Mux.scala 31:69:@45546.4]
  wire  _T_1899; // @[MemPrimitives.scala 82:228:@45555.4]
  wire  _T_1900; // @[MemPrimitives.scala 83:102:@45556.4]
  wire  _T_1905; // @[MemPrimitives.scala 82:228:@45559.4]
  wire  _T_1906; // @[MemPrimitives.scala 83:102:@45560.4]
  wire  _T_1911; // @[MemPrimitives.scala 82:228:@45563.4]
  wire  _T_1912; // @[MemPrimitives.scala 83:102:@45564.4]
  wire  _T_1917; // @[MemPrimitives.scala 82:228:@45567.4]
  wire  _T_1918; // @[MemPrimitives.scala 83:102:@45568.4]
  wire [16:0] _T_1920; // @[Cat.scala 30:58:@45570.4]
  wire [16:0] _T_1922; // @[Cat.scala 30:58:@45572.4]
  wire [16:0] _T_1924; // @[Cat.scala 30:58:@45574.4]
  wire [16:0] _T_1926; // @[Cat.scala 30:58:@45576.4]
  wire [16:0] _T_1927; // @[Mux.scala 31:69:@45577.4]
  wire [16:0] _T_1928; // @[Mux.scala 31:69:@45578.4]
  wire [16:0] _T_1929; // @[Mux.scala 31:69:@45579.4]
  wire  _T_1937; // @[MemPrimitives.scala 82:228:@45588.4]
  wire  _T_1938; // @[MemPrimitives.scala 83:102:@45589.4]
  wire  _T_1943; // @[MemPrimitives.scala 82:228:@45592.4]
  wire  _T_1944; // @[MemPrimitives.scala 83:102:@45593.4]
  wire  _T_1949; // @[MemPrimitives.scala 82:228:@45596.4]
  wire  _T_1950; // @[MemPrimitives.scala 83:102:@45597.4]
  wire  _T_1955; // @[MemPrimitives.scala 82:228:@45600.4]
  wire  _T_1956; // @[MemPrimitives.scala 83:102:@45601.4]
  wire [16:0] _T_1958; // @[Cat.scala 30:58:@45603.4]
  wire [16:0] _T_1960; // @[Cat.scala 30:58:@45605.4]
  wire [16:0] _T_1962; // @[Cat.scala 30:58:@45607.4]
  wire [16:0] _T_1964; // @[Cat.scala 30:58:@45609.4]
  wire [16:0] _T_1965; // @[Mux.scala 31:69:@45610.4]
  wire [16:0] _T_1966; // @[Mux.scala 31:69:@45611.4]
  wire [16:0] _T_1967; // @[Mux.scala 31:69:@45612.4]
  wire  _T_1972; // @[MemPrimitives.scala 82:210:@45619.4]
  wire  _T_1975; // @[MemPrimitives.scala 82:228:@45621.4]
  wire  _T_1976; // @[MemPrimitives.scala 83:102:@45622.4]
  wire  _T_1978; // @[MemPrimitives.scala 82:210:@45623.4]
  wire  _T_1981; // @[MemPrimitives.scala 82:228:@45625.4]
  wire  _T_1982; // @[MemPrimitives.scala 83:102:@45626.4]
  wire  _T_1984; // @[MemPrimitives.scala 82:210:@45627.4]
  wire  _T_1987; // @[MemPrimitives.scala 82:228:@45629.4]
  wire  _T_1988; // @[MemPrimitives.scala 83:102:@45630.4]
  wire  _T_1990; // @[MemPrimitives.scala 82:210:@45631.4]
  wire  _T_1993; // @[MemPrimitives.scala 82:228:@45633.4]
  wire  _T_1994; // @[MemPrimitives.scala 83:102:@45634.4]
  wire [16:0] _T_1996; // @[Cat.scala 30:58:@45636.4]
  wire [16:0] _T_1998; // @[Cat.scala 30:58:@45638.4]
  wire [16:0] _T_2000; // @[Cat.scala 30:58:@45640.4]
  wire [16:0] _T_2002; // @[Cat.scala 30:58:@45642.4]
  wire [16:0] _T_2003; // @[Mux.scala 31:69:@45643.4]
  wire [16:0] _T_2004; // @[Mux.scala 31:69:@45644.4]
  wire [16:0] _T_2005; // @[Mux.scala 31:69:@45645.4]
  wire  _T_2010; // @[MemPrimitives.scala 82:210:@45652.4]
  wire  _T_2013; // @[MemPrimitives.scala 82:228:@45654.4]
  wire  _T_2014; // @[MemPrimitives.scala 83:102:@45655.4]
  wire  _T_2016; // @[MemPrimitives.scala 82:210:@45656.4]
  wire  _T_2019; // @[MemPrimitives.scala 82:228:@45658.4]
  wire  _T_2020; // @[MemPrimitives.scala 83:102:@45659.4]
  wire  _T_2022; // @[MemPrimitives.scala 82:210:@45660.4]
  wire  _T_2025; // @[MemPrimitives.scala 82:228:@45662.4]
  wire  _T_2026; // @[MemPrimitives.scala 83:102:@45663.4]
  wire  _T_2028; // @[MemPrimitives.scala 82:210:@45664.4]
  wire  _T_2031; // @[MemPrimitives.scala 82:228:@45666.4]
  wire  _T_2032; // @[MemPrimitives.scala 83:102:@45667.4]
  wire [16:0] _T_2034; // @[Cat.scala 30:58:@45669.4]
  wire [16:0] _T_2036; // @[Cat.scala 30:58:@45671.4]
  wire [16:0] _T_2038; // @[Cat.scala 30:58:@45673.4]
  wire [16:0] _T_2040; // @[Cat.scala 30:58:@45675.4]
  wire [16:0] _T_2041; // @[Mux.scala 31:69:@45676.4]
  wire [16:0] _T_2042; // @[Mux.scala 31:69:@45677.4]
  wire [16:0] _T_2043; // @[Mux.scala 31:69:@45678.4]
  wire  _T_2051; // @[MemPrimitives.scala 82:228:@45687.4]
  wire  _T_2052; // @[MemPrimitives.scala 83:102:@45688.4]
  wire  _T_2057; // @[MemPrimitives.scala 82:228:@45691.4]
  wire  _T_2058; // @[MemPrimitives.scala 83:102:@45692.4]
  wire  _T_2063; // @[MemPrimitives.scala 82:228:@45695.4]
  wire  _T_2064; // @[MemPrimitives.scala 83:102:@45696.4]
  wire  _T_2069; // @[MemPrimitives.scala 82:228:@45699.4]
  wire  _T_2070; // @[MemPrimitives.scala 83:102:@45700.4]
  wire [16:0] _T_2072; // @[Cat.scala 30:58:@45702.4]
  wire [16:0] _T_2074; // @[Cat.scala 30:58:@45704.4]
  wire [16:0] _T_2076; // @[Cat.scala 30:58:@45706.4]
  wire [16:0] _T_2078; // @[Cat.scala 30:58:@45708.4]
  wire [16:0] _T_2079; // @[Mux.scala 31:69:@45709.4]
  wire [16:0] _T_2080; // @[Mux.scala 31:69:@45710.4]
  wire [16:0] _T_2081; // @[Mux.scala 31:69:@45711.4]
  wire  _T_2089; // @[MemPrimitives.scala 82:228:@45720.4]
  wire  _T_2090; // @[MemPrimitives.scala 83:102:@45721.4]
  wire  _T_2095; // @[MemPrimitives.scala 82:228:@45724.4]
  wire  _T_2096; // @[MemPrimitives.scala 83:102:@45725.4]
  wire  _T_2101; // @[MemPrimitives.scala 82:228:@45728.4]
  wire  _T_2102; // @[MemPrimitives.scala 83:102:@45729.4]
  wire  _T_2107; // @[MemPrimitives.scala 82:228:@45732.4]
  wire  _T_2108; // @[MemPrimitives.scala 83:102:@45733.4]
  wire [16:0] _T_2110; // @[Cat.scala 30:58:@45735.4]
  wire [16:0] _T_2112; // @[Cat.scala 30:58:@45737.4]
  wire [16:0] _T_2114; // @[Cat.scala 30:58:@45739.4]
  wire [16:0] _T_2116; // @[Cat.scala 30:58:@45741.4]
  wire [16:0] _T_2117; // @[Mux.scala 31:69:@45742.4]
  wire [16:0] _T_2118; // @[Mux.scala 31:69:@45743.4]
  wire [16:0] _T_2119; // @[Mux.scala 31:69:@45744.4]
  wire  _T_2127; // @[MemPrimitives.scala 82:228:@45753.4]
  wire  _T_2128; // @[MemPrimitives.scala 83:102:@45754.4]
  wire  _T_2133; // @[MemPrimitives.scala 82:228:@45757.4]
  wire  _T_2134; // @[MemPrimitives.scala 83:102:@45758.4]
  wire  _T_2139; // @[MemPrimitives.scala 82:228:@45761.4]
  wire  _T_2140; // @[MemPrimitives.scala 83:102:@45762.4]
  wire  _T_2145; // @[MemPrimitives.scala 82:228:@45765.4]
  wire  _T_2146; // @[MemPrimitives.scala 83:102:@45766.4]
  wire [16:0] _T_2148; // @[Cat.scala 30:58:@45768.4]
  wire [16:0] _T_2150; // @[Cat.scala 30:58:@45770.4]
  wire [16:0] _T_2152; // @[Cat.scala 30:58:@45772.4]
  wire [16:0] _T_2154; // @[Cat.scala 30:58:@45774.4]
  wire [16:0] _T_2155; // @[Mux.scala 31:69:@45775.4]
  wire [16:0] _T_2156; // @[Mux.scala 31:69:@45776.4]
  wire [16:0] _T_2157; // @[Mux.scala 31:69:@45777.4]
  wire  _T_2165; // @[MemPrimitives.scala 82:228:@45786.4]
  wire  _T_2166; // @[MemPrimitives.scala 83:102:@45787.4]
  wire  _T_2171; // @[MemPrimitives.scala 82:228:@45790.4]
  wire  _T_2172; // @[MemPrimitives.scala 83:102:@45791.4]
  wire  _T_2177; // @[MemPrimitives.scala 82:228:@45794.4]
  wire  _T_2178; // @[MemPrimitives.scala 83:102:@45795.4]
  wire  _T_2183; // @[MemPrimitives.scala 82:228:@45798.4]
  wire  _T_2184; // @[MemPrimitives.scala 83:102:@45799.4]
  wire [16:0] _T_2186; // @[Cat.scala 30:58:@45801.4]
  wire [16:0] _T_2188; // @[Cat.scala 30:58:@45803.4]
  wire [16:0] _T_2190; // @[Cat.scala 30:58:@45805.4]
  wire [16:0] _T_2192; // @[Cat.scala 30:58:@45807.4]
  wire [16:0] _T_2193; // @[Mux.scala 31:69:@45808.4]
  wire [16:0] _T_2194; // @[Mux.scala 31:69:@45809.4]
  wire [16:0] _T_2195; // @[Mux.scala 31:69:@45810.4]
  wire  _T_2203; // @[MemPrimitives.scala 82:228:@45819.4]
  wire  _T_2204; // @[MemPrimitives.scala 83:102:@45820.4]
  wire  _T_2209; // @[MemPrimitives.scala 82:228:@45823.4]
  wire  _T_2210; // @[MemPrimitives.scala 83:102:@45824.4]
  wire  _T_2215; // @[MemPrimitives.scala 82:228:@45827.4]
  wire  _T_2216; // @[MemPrimitives.scala 83:102:@45828.4]
  wire  _T_2221; // @[MemPrimitives.scala 82:228:@45831.4]
  wire  _T_2222; // @[MemPrimitives.scala 83:102:@45832.4]
  wire [16:0] _T_2224; // @[Cat.scala 30:58:@45834.4]
  wire [16:0] _T_2226; // @[Cat.scala 30:58:@45836.4]
  wire [16:0] _T_2228; // @[Cat.scala 30:58:@45838.4]
  wire [16:0] _T_2230; // @[Cat.scala 30:58:@45840.4]
  wire [16:0] _T_2231; // @[Mux.scala 31:69:@45841.4]
  wire [16:0] _T_2232; // @[Mux.scala 31:69:@45842.4]
  wire [16:0] _T_2233; // @[Mux.scala 31:69:@45843.4]
  wire  _T_2241; // @[MemPrimitives.scala 82:228:@45852.4]
  wire  _T_2242; // @[MemPrimitives.scala 83:102:@45853.4]
  wire  _T_2247; // @[MemPrimitives.scala 82:228:@45856.4]
  wire  _T_2248; // @[MemPrimitives.scala 83:102:@45857.4]
  wire  _T_2253; // @[MemPrimitives.scala 82:228:@45860.4]
  wire  _T_2254; // @[MemPrimitives.scala 83:102:@45861.4]
  wire  _T_2259; // @[MemPrimitives.scala 82:228:@45864.4]
  wire  _T_2260; // @[MemPrimitives.scala 83:102:@45865.4]
  wire [16:0] _T_2262; // @[Cat.scala 30:58:@45867.4]
  wire [16:0] _T_2264; // @[Cat.scala 30:58:@45869.4]
  wire [16:0] _T_2266; // @[Cat.scala 30:58:@45871.4]
  wire [16:0] _T_2268; // @[Cat.scala 30:58:@45873.4]
  wire [16:0] _T_2269; // @[Mux.scala 31:69:@45874.4]
  wire [16:0] _T_2270; // @[Mux.scala 31:69:@45875.4]
  wire [16:0] _T_2271; // @[Mux.scala 31:69:@45876.4]
  wire  _T_2279; // @[MemPrimitives.scala 82:228:@45885.4]
  wire  _T_2280; // @[MemPrimitives.scala 83:102:@45886.4]
  wire  _T_2285; // @[MemPrimitives.scala 82:228:@45889.4]
  wire  _T_2286; // @[MemPrimitives.scala 83:102:@45890.4]
  wire  _T_2291; // @[MemPrimitives.scala 82:228:@45893.4]
  wire  _T_2292; // @[MemPrimitives.scala 83:102:@45894.4]
  wire  _T_2297; // @[MemPrimitives.scala 82:228:@45897.4]
  wire  _T_2298; // @[MemPrimitives.scala 83:102:@45898.4]
  wire [16:0] _T_2300; // @[Cat.scala 30:58:@45900.4]
  wire [16:0] _T_2302; // @[Cat.scala 30:58:@45902.4]
  wire [16:0] _T_2304; // @[Cat.scala 30:58:@45904.4]
  wire [16:0] _T_2306; // @[Cat.scala 30:58:@45906.4]
  wire [16:0] _T_2307; // @[Mux.scala 31:69:@45907.4]
  wire [16:0] _T_2308; // @[Mux.scala 31:69:@45908.4]
  wire [16:0] _T_2309; // @[Mux.scala 31:69:@45909.4]
  wire  _T_2317; // @[MemPrimitives.scala 82:228:@45918.4]
  wire  _T_2318; // @[MemPrimitives.scala 83:102:@45919.4]
  wire  _T_2323; // @[MemPrimitives.scala 82:228:@45922.4]
  wire  _T_2324; // @[MemPrimitives.scala 83:102:@45923.4]
  wire  _T_2329; // @[MemPrimitives.scala 82:228:@45926.4]
  wire  _T_2330; // @[MemPrimitives.scala 83:102:@45927.4]
  wire  _T_2335; // @[MemPrimitives.scala 82:228:@45930.4]
  wire  _T_2336; // @[MemPrimitives.scala 83:102:@45931.4]
  wire [16:0] _T_2338; // @[Cat.scala 30:58:@45933.4]
  wire [16:0] _T_2340; // @[Cat.scala 30:58:@45935.4]
  wire [16:0] _T_2342; // @[Cat.scala 30:58:@45937.4]
  wire [16:0] _T_2344; // @[Cat.scala 30:58:@45939.4]
  wire [16:0] _T_2345; // @[Mux.scala 31:69:@45940.4]
  wire [16:0] _T_2346; // @[Mux.scala 31:69:@45941.4]
  wire [16:0] _T_2347; // @[Mux.scala 31:69:@45942.4]
  wire  _T_2352; // @[MemPrimitives.scala 82:210:@45949.4]
  wire  _T_2355; // @[MemPrimitives.scala 82:228:@45951.4]
  wire  _T_2356; // @[MemPrimitives.scala 83:102:@45952.4]
  wire  _T_2358; // @[MemPrimitives.scala 82:210:@45953.4]
  wire  _T_2361; // @[MemPrimitives.scala 82:228:@45955.4]
  wire  _T_2362; // @[MemPrimitives.scala 83:102:@45956.4]
  wire  _T_2364; // @[MemPrimitives.scala 82:210:@45957.4]
  wire  _T_2367; // @[MemPrimitives.scala 82:228:@45959.4]
  wire  _T_2368; // @[MemPrimitives.scala 83:102:@45960.4]
  wire  _T_2370; // @[MemPrimitives.scala 82:210:@45961.4]
  wire  _T_2373; // @[MemPrimitives.scala 82:228:@45963.4]
  wire  _T_2374; // @[MemPrimitives.scala 83:102:@45964.4]
  wire [16:0] _T_2376; // @[Cat.scala 30:58:@45966.4]
  wire [16:0] _T_2378; // @[Cat.scala 30:58:@45968.4]
  wire [16:0] _T_2380; // @[Cat.scala 30:58:@45970.4]
  wire [16:0] _T_2382; // @[Cat.scala 30:58:@45972.4]
  wire [16:0] _T_2383; // @[Mux.scala 31:69:@45973.4]
  wire [16:0] _T_2384; // @[Mux.scala 31:69:@45974.4]
  wire [16:0] _T_2385; // @[Mux.scala 31:69:@45975.4]
  wire  _T_2390; // @[MemPrimitives.scala 82:210:@45982.4]
  wire  _T_2393; // @[MemPrimitives.scala 82:228:@45984.4]
  wire  _T_2394; // @[MemPrimitives.scala 83:102:@45985.4]
  wire  _T_2396; // @[MemPrimitives.scala 82:210:@45986.4]
  wire  _T_2399; // @[MemPrimitives.scala 82:228:@45988.4]
  wire  _T_2400; // @[MemPrimitives.scala 83:102:@45989.4]
  wire  _T_2402; // @[MemPrimitives.scala 82:210:@45990.4]
  wire  _T_2405; // @[MemPrimitives.scala 82:228:@45992.4]
  wire  _T_2406; // @[MemPrimitives.scala 83:102:@45993.4]
  wire  _T_2408; // @[MemPrimitives.scala 82:210:@45994.4]
  wire  _T_2411; // @[MemPrimitives.scala 82:228:@45996.4]
  wire  _T_2412; // @[MemPrimitives.scala 83:102:@45997.4]
  wire [16:0] _T_2414; // @[Cat.scala 30:58:@45999.4]
  wire [16:0] _T_2416; // @[Cat.scala 30:58:@46001.4]
  wire [16:0] _T_2418; // @[Cat.scala 30:58:@46003.4]
  wire [16:0] _T_2420; // @[Cat.scala 30:58:@46005.4]
  wire [16:0] _T_2421; // @[Mux.scala 31:69:@46006.4]
  wire [16:0] _T_2422; // @[Mux.scala 31:69:@46007.4]
  wire [16:0] _T_2423; // @[Mux.scala 31:69:@46008.4]
  wire  _T_2431; // @[MemPrimitives.scala 82:228:@46017.4]
  wire  _T_2432; // @[MemPrimitives.scala 83:102:@46018.4]
  wire  _T_2437; // @[MemPrimitives.scala 82:228:@46021.4]
  wire  _T_2438; // @[MemPrimitives.scala 83:102:@46022.4]
  wire  _T_2443; // @[MemPrimitives.scala 82:228:@46025.4]
  wire  _T_2444; // @[MemPrimitives.scala 83:102:@46026.4]
  wire  _T_2449; // @[MemPrimitives.scala 82:228:@46029.4]
  wire  _T_2450; // @[MemPrimitives.scala 83:102:@46030.4]
  wire [16:0] _T_2452; // @[Cat.scala 30:58:@46032.4]
  wire [16:0] _T_2454; // @[Cat.scala 30:58:@46034.4]
  wire [16:0] _T_2456; // @[Cat.scala 30:58:@46036.4]
  wire [16:0] _T_2458; // @[Cat.scala 30:58:@46038.4]
  wire [16:0] _T_2459; // @[Mux.scala 31:69:@46039.4]
  wire [16:0] _T_2460; // @[Mux.scala 31:69:@46040.4]
  wire [16:0] _T_2461; // @[Mux.scala 31:69:@46041.4]
  wire  _T_2469; // @[MemPrimitives.scala 82:228:@46050.4]
  wire  _T_2470; // @[MemPrimitives.scala 83:102:@46051.4]
  wire  _T_2475; // @[MemPrimitives.scala 82:228:@46054.4]
  wire  _T_2476; // @[MemPrimitives.scala 83:102:@46055.4]
  wire  _T_2481; // @[MemPrimitives.scala 82:228:@46058.4]
  wire  _T_2482; // @[MemPrimitives.scala 83:102:@46059.4]
  wire  _T_2487; // @[MemPrimitives.scala 82:228:@46062.4]
  wire  _T_2488; // @[MemPrimitives.scala 83:102:@46063.4]
  wire [16:0] _T_2490; // @[Cat.scala 30:58:@46065.4]
  wire [16:0] _T_2492; // @[Cat.scala 30:58:@46067.4]
  wire [16:0] _T_2494; // @[Cat.scala 30:58:@46069.4]
  wire [16:0] _T_2496; // @[Cat.scala 30:58:@46071.4]
  wire [16:0] _T_2497; // @[Mux.scala 31:69:@46072.4]
  wire [16:0] _T_2498; // @[Mux.scala 31:69:@46073.4]
  wire [16:0] _T_2499; // @[Mux.scala 31:69:@46074.4]
  wire  _T_2507; // @[MemPrimitives.scala 82:228:@46083.4]
  wire  _T_2508; // @[MemPrimitives.scala 83:102:@46084.4]
  wire  _T_2513; // @[MemPrimitives.scala 82:228:@46087.4]
  wire  _T_2514; // @[MemPrimitives.scala 83:102:@46088.4]
  wire  _T_2519; // @[MemPrimitives.scala 82:228:@46091.4]
  wire  _T_2520; // @[MemPrimitives.scala 83:102:@46092.4]
  wire  _T_2525; // @[MemPrimitives.scala 82:228:@46095.4]
  wire  _T_2526; // @[MemPrimitives.scala 83:102:@46096.4]
  wire [16:0] _T_2528; // @[Cat.scala 30:58:@46098.4]
  wire [16:0] _T_2530; // @[Cat.scala 30:58:@46100.4]
  wire [16:0] _T_2532; // @[Cat.scala 30:58:@46102.4]
  wire [16:0] _T_2534; // @[Cat.scala 30:58:@46104.4]
  wire [16:0] _T_2535; // @[Mux.scala 31:69:@46105.4]
  wire [16:0] _T_2536; // @[Mux.scala 31:69:@46106.4]
  wire [16:0] _T_2537; // @[Mux.scala 31:69:@46107.4]
  wire  _T_2545; // @[MemPrimitives.scala 82:228:@46116.4]
  wire  _T_2546; // @[MemPrimitives.scala 83:102:@46117.4]
  wire  _T_2551; // @[MemPrimitives.scala 82:228:@46120.4]
  wire  _T_2552; // @[MemPrimitives.scala 83:102:@46121.4]
  wire  _T_2557; // @[MemPrimitives.scala 82:228:@46124.4]
  wire  _T_2558; // @[MemPrimitives.scala 83:102:@46125.4]
  wire  _T_2563; // @[MemPrimitives.scala 82:228:@46128.4]
  wire  _T_2564; // @[MemPrimitives.scala 83:102:@46129.4]
  wire [16:0] _T_2566; // @[Cat.scala 30:58:@46131.4]
  wire [16:0] _T_2568; // @[Cat.scala 30:58:@46133.4]
  wire [16:0] _T_2570; // @[Cat.scala 30:58:@46135.4]
  wire [16:0] _T_2572; // @[Cat.scala 30:58:@46137.4]
  wire [16:0] _T_2573; // @[Mux.scala 31:69:@46138.4]
  wire [16:0] _T_2574; // @[Mux.scala 31:69:@46139.4]
  wire [16:0] _T_2575; // @[Mux.scala 31:69:@46140.4]
  wire  _T_2583; // @[MemPrimitives.scala 82:228:@46149.4]
  wire  _T_2584; // @[MemPrimitives.scala 83:102:@46150.4]
  wire  _T_2589; // @[MemPrimitives.scala 82:228:@46153.4]
  wire  _T_2590; // @[MemPrimitives.scala 83:102:@46154.4]
  wire  _T_2595; // @[MemPrimitives.scala 82:228:@46157.4]
  wire  _T_2596; // @[MemPrimitives.scala 83:102:@46158.4]
  wire  _T_2601; // @[MemPrimitives.scala 82:228:@46161.4]
  wire  _T_2602; // @[MemPrimitives.scala 83:102:@46162.4]
  wire [16:0] _T_2604; // @[Cat.scala 30:58:@46164.4]
  wire [16:0] _T_2606; // @[Cat.scala 30:58:@46166.4]
  wire [16:0] _T_2608; // @[Cat.scala 30:58:@46168.4]
  wire [16:0] _T_2610; // @[Cat.scala 30:58:@46170.4]
  wire [16:0] _T_2611; // @[Mux.scala 31:69:@46171.4]
  wire [16:0] _T_2612; // @[Mux.scala 31:69:@46172.4]
  wire [16:0] _T_2613; // @[Mux.scala 31:69:@46173.4]
  wire  _T_2621; // @[MemPrimitives.scala 82:228:@46182.4]
  wire  _T_2622; // @[MemPrimitives.scala 83:102:@46183.4]
  wire  _T_2627; // @[MemPrimitives.scala 82:228:@46186.4]
  wire  _T_2628; // @[MemPrimitives.scala 83:102:@46187.4]
  wire  _T_2633; // @[MemPrimitives.scala 82:228:@46190.4]
  wire  _T_2634; // @[MemPrimitives.scala 83:102:@46191.4]
  wire  _T_2639; // @[MemPrimitives.scala 82:228:@46194.4]
  wire  _T_2640; // @[MemPrimitives.scala 83:102:@46195.4]
  wire [16:0] _T_2642; // @[Cat.scala 30:58:@46197.4]
  wire [16:0] _T_2644; // @[Cat.scala 30:58:@46199.4]
  wire [16:0] _T_2646; // @[Cat.scala 30:58:@46201.4]
  wire [16:0] _T_2648; // @[Cat.scala 30:58:@46203.4]
  wire [16:0] _T_2649; // @[Mux.scala 31:69:@46204.4]
  wire [16:0] _T_2650; // @[Mux.scala 31:69:@46205.4]
  wire [16:0] _T_2651; // @[Mux.scala 31:69:@46206.4]
  wire  _T_2659; // @[MemPrimitives.scala 82:228:@46215.4]
  wire  _T_2660; // @[MemPrimitives.scala 83:102:@46216.4]
  wire  _T_2665; // @[MemPrimitives.scala 82:228:@46219.4]
  wire  _T_2666; // @[MemPrimitives.scala 83:102:@46220.4]
  wire  _T_2671; // @[MemPrimitives.scala 82:228:@46223.4]
  wire  _T_2672; // @[MemPrimitives.scala 83:102:@46224.4]
  wire  _T_2677; // @[MemPrimitives.scala 82:228:@46227.4]
  wire  _T_2678; // @[MemPrimitives.scala 83:102:@46228.4]
  wire [16:0] _T_2680; // @[Cat.scala 30:58:@46230.4]
  wire [16:0] _T_2682; // @[Cat.scala 30:58:@46232.4]
  wire [16:0] _T_2684; // @[Cat.scala 30:58:@46234.4]
  wire [16:0] _T_2686; // @[Cat.scala 30:58:@46236.4]
  wire [16:0] _T_2687; // @[Mux.scala 31:69:@46237.4]
  wire [16:0] _T_2688; // @[Mux.scala 31:69:@46238.4]
  wire [16:0] _T_2689; // @[Mux.scala 31:69:@46239.4]
  wire  _T_2697; // @[MemPrimitives.scala 82:228:@46248.4]
  wire  _T_2698; // @[MemPrimitives.scala 83:102:@46249.4]
  wire  _T_2703; // @[MemPrimitives.scala 82:228:@46252.4]
  wire  _T_2704; // @[MemPrimitives.scala 83:102:@46253.4]
  wire  _T_2709; // @[MemPrimitives.scala 82:228:@46256.4]
  wire  _T_2710; // @[MemPrimitives.scala 83:102:@46257.4]
  wire  _T_2715; // @[MemPrimitives.scala 82:228:@46260.4]
  wire  _T_2716; // @[MemPrimitives.scala 83:102:@46261.4]
  wire [16:0] _T_2718; // @[Cat.scala 30:58:@46263.4]
  wire [16:0] _T_2720; // @[Cat.scala 30:58:@46265.4]
  wire [16:0] _T_2722; // @[Cat.scala 30:58:@46267.4]
  wire [16:0] _T_2724; // @[Cat.scala 30:58:@46269.4]
  wire [16:0] _T_2725; // @[Mux.scala 31:69:@46270.4]
  wire [16:0] _T_2726; // @[Mux.scala 31:69:@46271.4]
  wire [16:0] _T_2727; // @[Mux.scala 31:69:@46272.4]
  wire  _T_2732; // @[MemPrimitives.scala 110:210:@46279.4]
  wire  _T_2734; // @[MemPrimitives.scala 110:210:@46280.4]
  wire  _T_2735; // @[MemPrimitives.scala 110:228:@46281.4]
  wire  _T_2738; // @[MemPrimitives.scala 110:210:@46283.4]
  wire  _T_2740; // @[MemPrimitives.scala 110:210:@46284.4]
  wire  _T_2741; // @[MemPrimitives.scala 110:228:@46285.4]
  wire  _T_2744; // @[MemPrimitives.scala 110:210:@46287.4]
  wire  _T_2746; // @[MemPrimitives.scala 110:210:@46288.4]
  wire  _T_2747; // @[MemPrimitives.scala 110:228:@46289.4]
  wire  _T_2750; // @[MemPrimitives.scala 110:210:@46291.4]
  wire  _T_2752; // @[MemPrimitives.scala 110:210:@46292.4]
  wire  _T_2753; // @[MemPrimitives.scala 110:228:@46293.4]
  wire  _T_2756; // @[MemPrimitives.scala 110:210:@46295.4]
  wire  _T_2758; // @[MemPrimitives.scala 110:210:@46296.4]
  wire  _T_2759; // @[MemPrimitives.scala 110:228:@46297.4]
  wire  _T_2762; // @[MemPrimitives.scala 110:210:@46299.4]
  wire  _T_2764; // @[MemPrimitives.scala 110:210:@46300.4]
  wire  _T_2765; // @[MemPrimitives.scala 110:228:@46301.4]
  wire  _T_2768; // @[MemPrimitives.scala 110:210:@46303.4]
  wire  _T_2770; // @[MemPrimitives.scala 110:210:@46304.4]
  wire  _T_2771; // @[MemPrimitives.scala 110:228:@46305.4]
  wire  _T_2774; // @[MemPrimitives.scala 110:210:@46307.4]
  wire  _T_2776; // @[MemPrimitives.scala 110:210:@46308.4]
  wire  _T_2777; // @[MemPrimitives.scala 110:228:@46309.4]
  wire  _T_2780; // @[MemPrimitives.scala 110:210:@46311.4]
  wire  _T_2782; // @[MemPrimitives.scala 110:210:@46312.4]
  wire  _T_2783; // @[MemPrimitives.scala 110:228:@46313.4]
  wire  _T_2786; // @[MemPrimitives.scala 110:210:@46315.4]
  wire  _T_2788; // @[MemPrimitives.scala 110:210:@46316.4]
  wire  _T_2789; // @[MemPrimitives.scala 110:228:@46317.4]
  wire  _T_2792; // @[MemPrimitives.scala 110:210:@46319.4]
  wire  _T_2794; // @[MemPrimitives.scala 110:210:@46320.4]
  wire  _T_2795; // @[MemPrimitives.scala 110:228:@46321.4]
  wire  _T_2798; // @[MemPrimitives.scala 110:210:@46323.4]
  wire  _T_2800; // @[MemPrimitives.scala 110:210:@46324.4]
  wire  _T_2801; // @[MemPrimitives.scala 110:228:@46325.4]
  wire  _T_2804; // @[MemPrimitives.scala 110:210:@46327.4]
  wire  _T_2806; // @[MemPrimitives.scala 110:210:@46328.4]
  wire  _T_2807; // @[MemPrimitives.scala 110:228:@46329.4]
  wire  _T_2810; // @[MemPrimitives.scala 110:210:@46331.4]
  wire  _T_2812; // @[MemPrimitives.scala 110:210:@46332.4]
  wire  _T_2813; // @[MemPrimitives.scala 110:228:@46333.4]
  wire  _T_2816; // @[MemPrimitives.scala 110:210:@46335.4]
  wire  _T_2818; // @[MemPrimitives.scala 110:210:@46336.4]
  wire  _T_2819; // @[MemPrimitives.scala 110:228:@46337.4]
  wire  _T_2821; // @[MemPrimitives.scala 123:41:@46357.4]
  wire  _T_2822; // @[MemPrimitives.scala 123:41:@46358.4]
  wire  _T_2823; // @[MemPrimitives.scala 123:41:@46359.4]
  wire  _T_2824; // @[MemPrimitives.scala 123:41:@46360.4]
  wire  _T_2825; // @[MemPrimitives.scala 123:41:@46361.4]
  wire  _T_2826; // @[MemPrimitives.scala 123:41:@46362.4]
  wire  _T_2827; // @[MemPrimitives.scala 123:41:@46363.4]
  wire  _T_2828; // @[MemPrimitives.scala 123:41:@46364.4]
  wire  _T_2829; // @[MemPrimitives.scala 123:41:@46365.4]
  wire  _T_2830; // @[MemPrimitives.scala 123:41:@46366.4]
  wire  _T_2831; // @[MemPrimitives.scala 123:41:@46367.4]
  wire  _T_2832; // @[MemPrimitives.scala 123:41:@46368.4]
  wire  _T_2833; // @[MemPrimitives.scala 123:41:@46369.4]
  wire  _T_2834; // @[MemPrimitives.scala 123:41:@46370.4]
  wire  _T_2835; // @[MemPrimitives.scala 123:41:@46371.4]
  wire [9:0] _T_2837; // @[Cat.scala 30:58:@46373.4]
  wire [9:0] _T_2839; // @[Cat.scala 30:58:@46375.4]
  wire [9:0] _T_2841; // @[Cat.scala 30:58:@46377.4]
  wire [9:0] _T_2843; // @[Cat.scala 30:58:@46379.4]
  wire [9:0] _T_2845; // @[Cat.scala 30:58:@46381.4]
  wire [9:0] _T_2847; // @[Cat.scala 30:58:@46383.4]
  wire [9:0] _T_2849; // @[Cat.scala 30:58:@46385.4]
  wire [9:0] _T_2851; // @[Cat.scala 30:58:@46387.4]
  wire [9:0] _T_2853; // @[Cat.scala 30:58:@46389.4]
  wire [9:0] _T_2855; // @[Cat.scala 30:58:@46391.4]
  wire [9:0] _T_2857; // @[Cat.scala 30:58:@46393.4]
  wire [9:0] _T_2859; // @[Cat.scala 30:58:@46395.4]
  wire [9:0] _T_2861; // @[Cat.scala 30:58:@46397.4]
  wire [9:0] _T_2863; // @[Cat.scala 30:58:@46399.4]
  wire [9:0] _T_2865; // @[Cat.scala 30:58:@46401.4]
  wire [9:0] _T_2866; // @[Mux.scala 31:69:@46402.4]
  wire [9:0] _T_2867; // @[Mux.scala 31:69:@46403.4]
  wire [9:0] _T_2868; // @[Mux.scala 31:69:@46404.4]
  wire [9:0] _T_2869; // @[Mux.scala 31:69:@46405.4]
  wire [9:0] _T_2870; // @[Mux.scala 31:69:@46406.4]
  wire [9:0] _T_2871; // @[Mux.scala 31:69:@46407.4]
  wire [9:0] _T_2872; // @[Mux.scala 31:69:@46408.4]
  wire [9:0] _T_2873; // @[Mux.scala 31:69:@46409.4]
  wire [9:0] _T_2874; // @[Mux.scala 31:69:@46410.4]
  wire [9:0] _T_2875; // @[Mux.scala 31:69:@46411.4]
  wire [9:0] _T_2876; // @[Mux.scala 31:69:@46412.4]
  wire [9:0] _T_2877; // @[Mux.scala 31:69:@46413.4]
  wire [9:0] _T_2878; // @[Mux.scala 31:69:@46414.4]
  wire [9:0] _T_2879; // @[Mux.scala 31:69:@46415.4]
  wire  _T_2884; // @[MemPrimitives.scala 110:210:@46422.4]
  wire  _T_2886; // @[MemPrimitives.scala 110:210:@46423.4]
  wire  _T_2887; // @[MemPrimitives.scala 110:228:@46424.4]
  wire  _T_2890; // @[MemPrimitives.scala 110:210:@46426.4]
  wire  _T_2892; // @[MemPrimitives.scala 110:210:@46427.4]
  wire  _T_2893; // @[MemPrimitives.scala 110:228:@46428.4]
  wire  _T_2896; // @[MemPrimitives.scala 110:210:@46430.4]
  wire  _T_2898; // @[MemPrimitives.scala 110:210:@46431.4]
  wire  _T_2899; // @[MemPrimitives.scala 110:228:@46432.4]
  wire  _T_2902; // @[MemPrimitives.scala 110:210:@46434.4]
  wire  _T_2904; // @[MemPrimitives.scala 110:210:@46435.4]
  wire  _T_2905; // @[MemPrimitives.scala 110:228:@46436.4]
  wire  _T_2908; // @[MemPrimitives.scala 110:210:@46438.4]
  wire  _T_2910; // @[MemPrimitives.scala 110:210:@46439.4]
  wire  _T_2911; // @[MemPrimitives.scala 110:228:@46440.4]
  wire  _T_2914; // @[MemPrimitives.scala 110:210:@46442.4]
  wire  _T_2916; // @[MemPrimitives.scala 110:210:@46443.4]
  wire  _T_2917; // @[MemPrimitives.scala 110:228:@46444.4]
  wire  _T_2920; // @[MemPrimitives.scala 110:210:@46446.4]
  wire  _T_2922; // @[MemPrimitives.scala 110:210:@46447.4]
  wire  _T_2923; // @[MemPrimitives.scala 110:228:@46448.4]
  wire  _T_2926; // @[MemPrimitives.scala 110:210:@46450.4]
  wire  _T_2928; // @[MemPrimitives.scala 110:210:@46451.4]
  wire  _T_2929; // @[MemPrimitives.scala 110:228:@46452.4]
  wire  _T_2932; // @[MemPrimitives.scala 110:210:@46454.4]
  wire  _T_2934; // @[MemPrimitives.scala 110:210:@46455.4]
  wire  _T_2935; // @[MemPrimitives.scala 110:228:@46456.4]
  wire  _T_2938; // @[MemPrimitives.scala 110:210:@46458.4]
  wire  _T_2940; // @[MemPrimitives.scala 110:210:@46459.4]
  wire  _T_2941; // @[MemPrimitives.scala 110:228:@46460.4]
  wire  _T_2944; // @[MemPrimitives.scala 110:210:@46462.4]
  wire  _T_2946; // @[MemPrimitives.scala 110:210:@46463.4]
  wire  _T_2947; // @[MemPrimitives.scala 110:228:@46464.4]
  wire  _T_2950; // @[MemPrimitives.scala 110:210:@46466.4]
  wire  _T_2952; // @[MemPrimitives.scala 110:210:@46467.4]
  wire  _T_2953; // @[MemPrimitives.scala 110:228:@46468.4]
  wire  _T_2956; // @[MemPrimitives.scala 110:210:@46470.4]
  wire  _T_2958; // @[MemPrimitives.scala 110:210:@46471.4]
  wire  _T_2959; // @[MemPrimitives.scala 110:228:@46472.4]
  wire  _T_2962; // @[MemPrimitives.scala 110:210:@46474.4]
  wire  _T_2964; // @[MemPrimitives.scala 110:210:@46475.4]
  wire  _T_2965; // @[MemPrimitives.scala 110:228:@46476.4]
  wire  _T_2968; // @[MemPrimitives.scala 110:210:@46478.4]
  wire  _T_2970; // @[MemPrimitives.scala 110:210:@46479.4]
  wire  _T_2971; // @[MemPrimitives.scala 110:228:@46480.4]
  wire  _T_2973; // @[MemPrimitives.scala 123:41:@46500.4]
  wire  _T_2974; // @[MemPrimitives.scala 123:41:@46501.4]
  wire  _T_2975; // @[MemPrimitives.scala 123:41:@46502.4]
  wire  _T_2976; // @[MemPrimitives.scala 123:41:@46503.4]
  wire  _T_2977; // @[MemPrimitives.scala 123:41:@46504.4]
  wire  _T_2978; // @[MemPrimitives.scala 123:41:@46505.4]
  wire  _T_2979; // @[MemPrimitives.scala 123:41:@46506.4]
  wire  _T_2980; // @[MemPrimitives.scala 123:41:@46507.4]
  wire  _T_2981; // @[MemPrimitives.scala 123:41:@46508.4]
  wire  _T_2982; // @[MemPrimitives.scala 123:41:@46509.4]
  wire  _T_2983; // @[MemPrimitives.scala 123:41:@46510.4]
  wire  _T_2984; // @[MemPrimitives.scala 123:41:@46511.4]
  wire  _T_2985; // @[MemPrimitives.scala 123:41:@46512.4]
  wire  _T_2986; // @[MemPrimitives.scala 123:41:@46513.4]
  wire  _T_2987; // @[MemPrimitives.scala 123:41:@46514.4]
  wire [9:0] _T_2989; // @[Cat.scala 30:58:@46516.4]
  wire [9:0] _T_2991; // @[Cat.scala 30:58:@46518.4]
  wire [9:0] _T_2993; // @[Cat.scala 30:58:@46520.4]
  wire [9:0] _T_2995; // @[Cat.scala 30:58:@46522.4]
  wire [9:0] _T_2997; // @[Cat.scala 30:58:@46524.4]
  wire [9:0] _T_2999; // @[Cat.scala 30:58:@46526.4]
  wire [9:0] _T_3001; // @[Cat.scala 30:58:@46528.4]
  wire [9:0] _T_3003; // @[Cat.scala 30:58:@46530.4]
  wire [9:0] _T_3005; // @[Cat.scala 30:58:@46532.4]
  wire [9:0] _T_3007; // @[Cat.scala 30:58:@46534.4]
  wire [9:0] _T_3009; // @[Cat.scala 30:58:@46536.4]
  wire [9:0] _T_3011; // @[Cat.scala 30:58:@46538.4]
  wire [9:0] _T_3013; // @[Cat.scala 30:58:@46540.4]
  wire [9:0] _T_3015; // @[Cat.scala 30:58:@46542.4]
  wire [9:0] _T_3017; // @[Cat.scala 30:58:@46544.4]
  wire [9:0] _T_3018; // @[Mux.scala 31:69:@46545.4]
  wire [9:0] _T_3019; // @[Mux.scala 31:69:@46546.4]
  wire [9:0] _T_3020; // @[Mux.scala 31:69:@46547.4]
  wire [9:0] _T_3021; // @[Mux.scala 31:69:@46548.4]
  wire [9:0] _T_3022; // @[Mux.scala 31:69:@46549.4]
  wire [9:0] _T_3023; // @[Mux.scala 31:69:@46550.4]
  wire [9:0] _T_3024; // @[Mux.scala 31:69:@46551.4]
  wire [9:0] _T_3025; // @[Mux.scala 31:69:@46552.4]
  wire [9:0] _T_3026; // @[Mux.scala 31:69:@46553.4]
  wire [9:0] _T_3027; // @[Mux.scala 31:69:@46554.4]
  wire [9:0] _T_3028; // @[Mux.scala 31:69:@46555.4]
  wire [9:0] _T_3029; // @[Mux.scala 31:69:@46556.4]
  wire [9:0] _T_3030; // @[Mux.scala 31:69:@46557.4]
  wire [9:0] _T_3031; // @[Mux.scala 31:69:@46558.4]
  wire  _T_3038; // @[MemPrimitives.scala 110:210:@46566.4]
  wire  _T_3039; // @[MemPrimitives.scala 110:228:@46567.4]
  wire  _T_3044; // @[MemPrimitives.scala 110:210:@46570.4]
  wire  _T_3045; // @[MemPrimitives.scala 110:228:@46571.4]
  wire  _T_3050; // @[MemPrimitives.scala 110:210:@46574.4]
  wire  _T_3051; // @[MemPrimitives.scala 110:228:@46575.4]
  wire  _T_3056; // @[MemPrimitives.scala 110:210:@46578.4]
  wire  _T_3057; // @[MemPrimitives.scala 110:228:@46579.4]
  wire  _T_3062; // @[MemPrimitives.scala 110:210:@46582.4]
  wire  _T_3063; // @[MemPrimitives.scala 110:228:@46583.4]
  wire  _T_3068; // @[MemPrimitives.scala 110:210:@46586.4]
  wire  _T_3069; // @[MemPrimitives.scala 110:228:@46587.4]
  wire  _T_3074; // @[MemPrimitives.scala 110:210:@46590.4]
  wire  _T_3075; // @[MemPrimitives.scala 110:228:@46591.4]
  wire  _T_3080; // @[MemPrimitives.scala 110:210:@46594.4]
  wire  _T_3081; // @[MemPrimitives.scala 110:228:@46595.4]
  wire  _T_3086; // @[MemPrimitives.scala 110:210:@46598.4]
  wire  _T_3087; // @[MemPrimitives.scala 110:228:@46599.4]
  wire  _T_3092; // @[MemPrimitives.scala 110:210:@46602.4]
  wire  _T_3093; // @[MemPrimitives.scala 110:228:@46603.4]
  wire  _T_3098; // @[MemPrimitives.scala 110:210:@46606.4]
  wire  _T_3099; // @[MemPrimitives.scala 110:228:@46607.4]
  wire  _T_3104; // @[MemPrimitives.scala 110:210:@46610.4]
  wire  _T_3105; // @[MemPrimitives.scala 110:228:@46611.4]
  wire  _T_3110; // @[MemPrimitives.scala 110:210:@46614.4]
  wire  _T_3111; // @[MemPrimitives.scala 110:228:@46615.4]
  wire  _T_3116; // @[MemPrimitives.scala 110:210:@46618.4]
  wire  _T_3117; // @[MemPrimitives.scala 110:228:@46619.4]
  wire  _T_3122; // @[MemPrimitives.scala 110:210:@46622.4]
  wire  _T_3123; // @[MemPrimitives.scala 110:228:@46623.4]
  wire  _T_3125; // @[MemPrimitives.scala 123:41:@46643.4]
  wire  _T_3126; // @[MemPrimitives.scala 123:41:@46644.4]
  wire  _T_3127; // @[MemPrimitives.scala 123:41:@46645.4]
  wire  _T_3128; // @[MemPrimitives.scala 123:41:@46646.4]
  wire  _T_3129; // @[MemPrimitives.scala 123:41:@46647.4]
  wire  _T_3130; // @[MemPrimitives.scala 123:41:@46648.4]
  wire  _T_3131; // @[MemPrimitives.scala 123:41:@46649.4]
  wire  _T_3132; // @[MemPrimitives.scala 123:41:@46650.4]
  wire  _T_3133; // @[MemPrimitives.scala 123:41:@46651.4]
  wire  _T_3134; // @[MemPrimitives.scala 123:41:@46652.4]
  wire  _T_3135; // @[MemPrimitives.scala 123:41:@46653.4]
  wire  _T_3136; // @[MemPrimitives.scala 123:41:@46654.4]
  wire  _T_3137; // @[MemPrimitives.scala 123:41:@46655.4]
  wire  _T_3138; // @[MemPrimitives.scala 123:41:@46656.4]
  wire  _T_3139; // @[MemPrimitives.scala 123:41:@46657.4]
  wire [9:0] _T_3141; // @[Cat.scala 30:58:@46659.4]
  wire [9:0] _T_3143; // @[Cat.scala 30:58:@46661.4]
  wire [9:0] _T_3145; // @[Cat.scala 30:58:@46663.4]
  wire [9:0] _T_3147; // @[Cat.scala 30:58:@46665.4]
  wire [9:0] _T_3149; // @[Cat.scala 30:58:@46667.4]
  wire [9:0] _T_3151; // @[Cat.scala 30:58:@46669.4]
  wire [9:0] _T_3153; // @[Cat.scala 30:58:@46671.4]
  wire [9:0] _T_3155; // @[Cat.scala 30:58:@46673.4]
  wire [9:0] _T_3157; // @[Cat.scala 30:58:@46675.4]
  wire [9:0] _T_3159; // @[Cat.scala 30:58:@46677.4]
  wire [9:0] _T_3161; // @[Cat.scala 30:58:@46679.4]
  wire [9:0] _T_3163; // @[Cat.scala 30:58:@46681.4]
  wire [9:0] _T_3165; // @[Cat.scala 30:58:@46683.4]
  wire [9:0] _T_3167; // @[Cat.scala 30:58:@46685.4]
  wire [9:0] _T_3169; // @[Cat.scala 30:58:@46687.4]
  wire [9:0] _T_3170; // @[Mux.scala 31:69:@46688.4]
  wire [9:0] _T_3171; // @[Mux.scala 31:69:@46689.4]
  wire [9:0] _T_3172; // @[Mux.scala 31:69:@46690.4]
  wire [9:0] _T_3173; // @[Mux.scala 31:69:@46691.4]
  wire [9:0] _T_3174; // @[Mux.scala 31:69:@46692.4]
  wire [9:0] _T_3175; // @[Mux.scala 31:69:@46693.4]
  wire [9:0] _T_3176; // @[Mux.scala 31:69:@46694.4]
  wire [9:0] _T_3177; // @[Mux.scala 31:69:@46695.4]
  wire [9:0] _T_3178; // @[Mux.scala 31:69:@46696.4]
  wire [9:0] _T_3179; // @[Mux.scala 31:69:@46697.4]
  wire [9:0] _T_3180; // @[Mux.scala 31:69:@46698.4]
  wire [9:0] _T_3181; // @[Mux.scala 31:69:@46699.4]
  wire [9:0] _T_3182; // @[Mux.scala 31:69:@46700.4]
  wire [9:0] _T_3183; // @[Mux.scala 31:69:@46701.4]
  wire  _T_3190; // @[MemPrimitives.scala 110:210:@46709.4]
  wire  _T_3191; // @[MemPrimitives.scala 110:228:@46710.4]
  wire  _T_3196; // @[MemPrimitives.scala 110:210:@46713.4]
  wire  _T_3197; // @[MemPrimitives.scala 110:228:@46714.4]
  wire  _T_3202; // @[MemPrimitives.scala 110:210:@46717.4]
  wire  _T_3203; // @[MemPrimitives.scala 110:228:@46718.4]
  wire  _T_3208; // @[MemPrimitives.scala 110:210:@46721.4]
  wire  _T_3209; // @[MemPrimitives.scala 110:228:@46722.4]
  wire  _T_3214; // @[MemPrimitives.scala 110:210:@46725.4]
  wire  _T_3215; // @[MemPrimitives.scala 110:228:@46726.4]
  wire  _T_3220; // @[MemPrimitives.scala 110:210:@46729.4]
  wire  _T_3221; // @[MemPrimitives.scala 110:228:@46730.4]
  wire  _T_3226; // @[MemPrimitives.scala 110:210:@46733.4]
  wire  _T_3227; // @[MemPrimitives.scala 110:228:@46734.4]
  wire  _T_3232; // @[MemPrimitives.scala 110:210:@46737.4]
  wire  _T_3233; // @[MemPrimitives.scala 110:228:@46738.4]
  wire  _T_3238; // @[MemPrimitives.scala 110:210:@46741.4]
  wire  _T_3239; // @[MemPrimitives.scala 110:228:@46742.4]
  wire  _T_3244; // @[MemPrimitives.scala 110:210:@46745.4]
  wire  _T_3245; // @[MemPrimitives.scala 110:228:@46746.4]
  wire  _T_3250; // @[MemPrimitives.scala 110:210:@46749.4]
  wire  _T_3251; // @[MemPrimitives.scala 110:228:@46750.4]
  wire  _T_3256; // @[MemPrimitives.scala 110:210:@46753.4]
  wire  _T_3257; // @[MemPrimitives.scala 110:228:@46754.4]
  wire  _T_3262; // @[MemPrimitives.scala 110:210:@46757.4]
  wire  _T_3263; // @[MemPrimitives.scala 110:228:@46758.4]
  wire  _T_3268; // @[MemPrimitives.scala 110:210:@46761.4]
  wire  _T_3269; // @[MemPrimitives.scala 110:228:@46762.4]
  wire  _T_3274; // @[MemPrimitives.scala 110:210:@46765.4]
  wire  _T_3275; // @[MemPrimitives.scala 110:228:@46766.4]
  wire  _T_3277; // @[MemPrimitives.scala 123:41:@46786.4]
  wire  _T_3278; // @[MemPrimitives.scala 123:41:@46787.4]
  wire  _T_3279; // @[MemPrimitives.scala 123:41:@46788.4]
  wire  _T_3280; // @[MemPrimitives.scala 123:41:@46789.4]
  wire  _T_3281; // @[MemPrimitives.scala 123:41:@46790.4]
  wire  _T_3282; // @[MemPrimitives.scala 123:41:@46791.4]
  wire  _T_3283; // @[MemPrimitives.scala 123:41:@46792.4]
  wire  _T_3284; // @[MemPrimitives.scala 123:41:@46793.4]
  wire  _T_3285; // @[MemPrimitives.scala 123:41:@46794.4]
  wire  _T_3286; // @[MemPrimitives.scala 123:41:@46795.4]
  wire  _T_3287; // @[MemPrimitives.scala 123:41:@46796.4]
  wire  _T_3288; // @[MemPrimitives.scala 123:41:@46797.4]
  wire  _T_3289; // @[MemPrimitives.scala 123:41:@46798.4]
  wire  _T_3290; // @[MemPrimitives.scala 123:41:@46799.4]
  wire  _T_3291; // @[MemPrimitives.scala 123:41:@46800.4]
  wire [9:0] _T_3293; // @[Cat.scala 30:58:@46802.4]
  wire [9:0] _T_3295; // @[Cat.scala 30:58:@46804.4]
  wire [9:0] _T_3297; // @[Cat.scala 30:58:@46806.4]
  wire [9:0] _T_3299; // @[Cat.scala 30:58:@46808.4]
  wire [9:0] _T_3301; // @[Cat.scala 30:58:@46810.4]
  wire [9:0] _T_3303; // @[Cat.scala 30:58:@46812.4]
  wire [9:0] _T_3305; // @[Cat.scala 30:58:@46814.4]
  wire [9:0] _T_3307; // @[Cat.scala 30:58:@46816.4]
  wire [9:0] _T_3309; // @[Cat.scala 30:58:@46818.4]
  wire [9:0] _T_3311; // @[Cat.scala 30:58:@46820.4]
  wire [9:0] _T_3313; // @[Cat.scala 30:58:@46822.4]
  wire [9:0] _T_3315; // @[Cat.scala 30:58:@46824.4]
  wire [9:0] _T_3317; // @[Cat.scala 30:58:@46826.4]
  wire [9:0] _T_3319; // @[Cat.scala 30:58:@46828.4]
  wire [9:0] _T_3321; // @[Cat.scala 30:58:@46830.4]
  wire [9:0] _T_3322; // @[Mux.scala 31:69:@46831.4]
  wire [9:0] _T_3323; // @[Mux.scala 31:69:@46832.4]
  wire [9:0] _T_3324; // @[Mux.scala 31:69:@46833.4]
  wire [9:0] _T_3325; // @[Mux.scala 31:69:@46834.4]
  wire [9:0] _T_3326; // @[Mux.scala 31:69:@46835.4]
  wire [9:0] _T_3327; // @[Mux.scala 31:69:@46836.4]
  wire [9:0] _T_3328; // @[Mux.scala 31:69:@46837.4]
  wire [9:0] _T_3329; // @[Mux.scala 31:69:@46838.4]
  wire [9:0] _T_3330; // @[Mux.scala 31:69:@46839.4]
  wire [9:0] _T_3331; // @[Mux.scala 31:69:@46840.4]
  wire [9:0] _T_3332; // @[Mux.scala 31:69:@46841.4]
  wire [9:0] _T_3333; // @[Mux.scala 31:69:@46842.4]
  wire [9:0] _T_3334; // @[Mux.scala 31:69:@46843.4]
  wire [9:0] _T_3335; // @[Mux.scala 31:69:@46844.4]
  wire  _T_3342; // @[MemPrimitives.scala 110:210:@46852.4]
  wire  _T_3343; // @[MemPrimitives.scala 110:228:@46853.4]
  wire  _T_3348; // @[MemPrimitives.scala 110:210:@46856.4]
  wire  _T_3349; // @[MemPrimitives.scala 110:228:@46857.4]
  wire  _T_3354; // @[MemPrimitives.scala 110:210:@46860.4]
  wire  _T_3355; // @[MemPrimitives.scala 110:228:@46861.4]
  wire  _T_3360; // @[MemPrimitives.scala 110:210:@46864.4]
  wire  _T_3361; // @[MemPrimitives.scala 110:228:@46865.4]
  wire  _T_3366; // @[MemPrimitives.scala 110:210:@46868.4]
  wire  _T_3367; // @[MemPrimitives.scala 110:228:@46869.4]
  wire  _T_3372; // @[MemPrimitives.scala 110:210:@46872.4]
  wire  _T_3373; // @[MemPrimitives.scala 110:228:@46873.4]
  wire  _T_3378; // @[MemPrimitives.scala 110:210:@46876.4]
  wire  _T_3379; // @[MemPrimitives.scala 110:228:@46877.4]
  wire  _T_3384; // @[MemPrimitives.scala 110:210:@46880.4]
  wire  _T_3385; // @[MemPrimitives.scala 110:228:@46881.4]
  wire  _T_3390; // @[MemPrimitives.scala 110:210:@46884.4]
  wire  _T_3391; // @[MemPrimitives.scala 110:228:@46885.4]
  wire  _T_3396; // @[MemPrimitives.scala 110:210:@46888.4]
  wire  _T_3397; // @[MemPrimitives.scala 110:228:@46889.4]
  wire  _T_3402; // @[MemPrimitives.scala 110:210:@46892.4]
  wire  _T_3403; // @[MemPrimitives.scala 110:228:@46893.4]
  wire  _T_3408; // @[MemPrimitives.scala 110:210:@46896.4]
  wire  _T_3409; // @[MemPrimitives.scala 110:228:@46897.4]
  wire  _T_3414; // @[MemPrimitives.scala 110:210:@46900.4]
  wire  _T_3415; // @[MemPrimitives.scala 110:228:@46901.4]
  wire  _T_3420; // @[MemPrimitives.scala 110:210:@46904.4]
  wire  _T_3421; // @[MemPrimitives.scala 110:228:@46905.4]
  wire  _T_3426; // @[MemPrimitives.scala 110:210:@46908.4]
  wire  _T_3427; // @[MemPrimitives.scala 110:228:@46909.4]
  wire  _T_3429; // @[MemPrimitives.scala 123:41:@46929.4]
  wire  _T_3430; // @[MemPrimitives.scala 123:41:@46930.4]
  wire  _T_3431; // @[MemPrimitives.scala 123:41:@46931.4]
  wire  _T_3432; // @[MemPrimitives.scala 123:41:@46932.4]
  wire  _T_3433; // @[MemPrimitives.scala 123:41:@46933.4]
  wire  _T_3434; // @[MemPrimitives.scala 123:41:@46934.4]
  wire  _T_3435; // @[MemPrimitives.scala 123:41:@46935.4]
  wire  _T_3436; // @[MemPrimitives.scala 123:41:@46936.4]
  wire  _T_3437; // @[MemPrimitives.scala 123:41:@46937.4]
  wire  _T_3438; // @[MemPrimitives.scala 123:41:@46938.4]
  wire  _T_3439; // @[MemPrimitives.scala 123:41:@46939.4]
  wire  _T_3440; // @[MemPrimitives.scala 123:41:@46940.4]
  wire  _T_3441; // @[MemPrimitives.scala 123:41:@46941.4]
  wire  _T_3442; // @[MemPrimitives.scala 123:41:@46942.4]
  wire  _T_3443; // @[MemPrimitives.scala 123:41:@46943.4]
  wire [9:0] _T_3445; // @[Cat.scala 30:58:@46945.4]
  wire [9:0] _T_3447; // @[Cat.scala 30:58:@46947.4]
  wire [9:0] _T_3449; // @[Cat.scala 30:58:@46949.4]
  wire [9:0] _T_3451; // @[Cat.scala 30:58:@46951.4]
  wire [9:0] _T_3453; // @[Cat.scala 30:58:@46953.4]
  wire [9:0] _T_3455; // @[Cat.scala 30:58:@46955.4]
  wire [9:0] _T_3457; // @[Cat.scala 30:58:@46957.4]
  wire [9:0] _T_3459; // @[Cat.scala 30:58:@46959.4]
  wire [9:0] _T_3461; // @[Cat.scala 30:58:@46961.4]
  wire [9:0] _T_3463; // @[Cat.scala 30:58:@46963.4]
  wire [9:0] _T_3465; // @[Cat.scala 30:58:@46965.4]
  wire [9:0] _T_3467; // @[Cat.scala 30:58:@46967.4]
  wire [9:0] _T_3469; // @[Cat.scala 30:58:@46969.4]
  wire [9:0] _T_3471; // @[Cat.scala 30:58:@46971.4]
  wire [9:0] _T_3473; // @[Cat.scala 30:58:@46973.4]
  wire [9:0] _T_3474; // @[Mux.scala 31:69:@46974.4]
  wire [9:0] _T_3475; // @[Mux.scala 31:69:@46975.4]
  wire [9:0] _T_3476; // @[Mux.scala 31:69:@46976.4]
  wire [9:0] _T_3477; // @[Mux.scala 31:69:@46977.4]
  wire [9:0] _T_3478; // @[Mux.scala 31:69:@46978.4]
  wire [9:0] _T_3479; // @[Mux.scala 31:69:@46979.4]
  wire [9:0] _T_3480; // @[Mux.scala 31:69:@46980.4]
  wire [9:0] _T_3481; // @[Mux.scala 31:69:@46981.4]
  wire [9:0] _T_3482; // @[Mux.scala 31:69:@46982.4]
  wire [9:0] _T_3483; // @[Mux.scala 31:69:@46983.4]
  wire [9:0] _T_3484; // @[Mux.scala 31:69:@46984.4]
  wire [9:0] _T_3485; // @[Mux.scala 31:69:@46985.4]
  wire [9:0] _T_3486; // @[Mux.scala 31:69:@46986.4]
  wire [9:0] _T_3487; // @[Mux.scala 31:69:@46987.4]
  wire  _T_3494; // @[MemPrimitives.scala 110:210:@46995.4]
  wire  _T_3495; // @[MemPrimitives.scala 110:228:@46996.4]
  wire  _T_3500; // @[MemPrimitives.scala 110:210:@46999.4]
  wire  _T_3501; // @[MemPrimitives.scala 110:228:@47000.4]
  wire  _T_3506; // @[MemPrimitives.scala 110:210:@47003.4]
  wire  _T_3507; // @[MemPrimitives.scala 110:228:@47004.4]
  wire  _T_3512; // @[MemPrimitives.scala 110:210:@47007.4]
  wire  _T_3513; // @[MemPrimitives.scala 110:228:@47008.4]
  wire  _T_3518; // @[MemPrimitives.scala 110:210:@47011.4]
  wire  _T_3519; // @[MemPrimitives.scala 110:228:@47012.4]
  wire  _T_3524; // @[MemPrimitives.scala 110:210:@47015.4]
  wire  _T_3525; // @[MemPrimitives.scala 110:228:@47016.4]
  wire  _T_3530; // @[MemPrimitives.scala 110:210:@47019.4]
  wire  _T_3531; // @[MemPrimitives.scala 110:228:@47020.4]
  wire  _T_3536; // @[MemPrimitives.scala 110:210:@47023.4]
  wire  _T_3537; // @[MemPrimitives.scala 110:228:@47024.4]
  wire  _T_3542; // @[MemPrimitives.scala 110:210:@47027.4]
  wire  _T_3543; // @[MemPrimitives.scala 110:228:@47028.4]
  wire  _T_3548; // @[MemPrimitives.scala 110:210:@47031.4]
  wire  _T_3549; // @[MemPrimitives.scala 110:228:@47032.4]
  wire  _T_3554; // @[MemPrimitives.scala 110:210:@47035.4]
  wire  _T_3555; // @[MemPrimitives.scala 110:228:@47036.4]
  wire  _T_3560; // @[MemPrimitives.scala 110:210:@47039.4]
  wire  _T_3561; // @[MemPrimitives.scala 110:228:@47040.4]
  wire  _T_3566; // @[MemPrimitives.scala 110:210:@47043.4]
  wire  _T_3567; // @[MemPrimitives.scala 110:228:@47044.4]
  wire  _T_3572; // @[MemPrimitives.scala 110:210:@47047.4]
  wire  _T_3573; // @[MemPrimitives.scala 110:228:@47048.4]
  wire  _T_3578; // @[MemPrimitives.scala 110:210:@47051.4]
  wire  _T_3579; // @[MemPrimitives.scala 110:228:@47052.4]
  wire  _T_3581; // @[MemPrimitives.scala 123:41:@47072.4]
  wire  _T_3582; // @[MemPrimitives.scala 123:41:@47073.4]
  wire  _T_3583; // @[MemPrimitives.scala 123:41:@47074.4]
  wire  _T_3584; // @[MemPrimitives.scala 123:41:@47075.4]
  wire  _T_3585; // @[MemPrimitives.scala 123:41:@47076.4]
  wire  _T_3586; // @[MemPrimitives.scala 123:41:@47077.4]
  wire  _T_3587; // @[MemPrimitives.scala 123:41:@47078.4]
  wire  _T_3588; // @[MemPrimitives.scala 123:41:@47079.4]
  wire  _T_3589; // @[MemPrimitives.scala 123:41:@47080.4]
  wire  _T_3590; // @[MemPrimitives.scala 123:41:@47081.4]
  wire  _T_3591; // @[MemPrimitives.scala 123:41:@47082.4]
  wire  _T_3592; // @[MemPrimitives.scala 123:41:@47083.4]
  wire  _T_3593; // @[MemPrimitives.scala 123:41:@47084.4]
  wire  _T_3594; // @[MemPrimitives.scala 123:41:@47085.4]
  wire  _T_3595; // @[MemPrimitives.scala 123:41:@47086.4]
  wire [9:0] _T_3597; // @[Cat.scala 30:58:@47088.4]
  wire [9:0] _T_3599; // @[Cat.scala 30:58:@47090.4]
  wire [9:0] _T_3601; // @[Cat.scala 30:58:@47092.4]
  wire [9:0] _T_3603; // @[Cat.scala 30:58:@47094.4]
  wire [9:0] _T_3605; // @[Cat.scala 30:58:@47096.4]
  wire [9:0] _T_3607; // @[Cat.scala 30:58:@47098.4]
  wire [9:0] _T_3609; // @[Cat.scala 30:58:@47100.4]
  wire [9:0] _T_3611; // @[Cat.scala 30:58:@47102.4]
  wire [9:0] _T_3613; // @[Cat.scala 30:58:@47104.4]
  wire [9:0] _T_3615; // @[Cat.scala 30:58:@47106.4]
  wire [9:0] _T_3617; // @[Cat.scala 30:58:@47108.4]
  wire [9:0] _T_3619; // @[Cat.scala 30:58:@47110.4]
  wire [9:0] _T_3621; // @[Cat.scala 30:58:@47112.4]
  wire [9:0] _T_3623; // @[Cat.scala 30:58:@47114.4]
  wire [9:0] _T_3625; // @[Cat.scala 30:58:@47116.4]
  wire [9:0] _T_3626; // @[Mux.scala 31:69:@47117.4]
  wire [9:0] _T_3627; // @[Mux.scala 31:69:@47118.4]
  wire [9:0] _T_3628; // @[Mux.scala 31:69:@47119.4]
  wire [9:0] _T_3629; // @[Mux.scala 31:69:@47120.4]
  wire [9:0] _T_3630; // @[Mux.scala 31:69:@47121.4]
  wire [9:0] _T_3631; // @[Mux.scala 31:69:@47122.4]
  wire [9:0] _T_3632; // @[Mux.scala 31:69:@47123.4]
  wire [9:0] _T_3633; // @[Mux.scala 31:69:@47124.4]
  wire [9:0] _T_3634; // @[Mux.scala 31:69:@47125.4]
  wire [9:0] _T_3635; // @[Mux.scala 31:69:@47126.4]
  wire [9:0] _T_3636; // @[Mux.scala 31:69:@47127.4]
  wire [9:0] _T_3637; // @[Mux.scala 31:69:@47128.4]
  wire [9:0] _T_3638; // @[Mux.scala 31:69:@47129.4]
  wire [9:0] _T_3639; // @[Mux.scala 31:69:@47130.4]
  wire  _T_3646; // @[MemPrimitives.scala 110:210:@47138.4]
  wire  _T_3647; // @[MemPrimitives.scala 110:228:@47139.4]
  wire  _T_3652; // @[MemPrimitives.scala 110:210:@47142.4]
  wire  _T_3653; // @[MemPrimitives.scala 110:228:@47143.4]
  wire  _T_3658; // @[MemPrimitives.scala 110:210:@47146.4]
  wire  _T_3659; // @[MemPrimitives.scala 110:228:@47147.4]
  wire  _T_3664; // @[MemPrimitives.scala 110:210:@47150.4]
  wire  _T_3665; // @[MemPrimitives.scala 110:228:@47151.4]
  wire  _T_3670; // @[MemPrimitives.scala 110:210:@47154.4]
  wire  _T_3671; // @[MemPrimitives.scala 110:228:@47155.4]
  wire  _T_3676; // @[MemPrimitives.scala 110:210:@47158.4]
  wire  _T_3677; // @[MemPrimitives.scala 110:228:@47159.4]
  wire  _T_3682; // @[MemPrimitives.scala 110:210:@47162.4]
  wire  _T_3683; // @[MemPrimitives.scala 110:228:@47163.4]
  wire  _T_3688; // @[MemPrimitives.scala 110:210:@47166.4]
  wire  _T_3689; // @[MemPrimitives.scala 110:228:@47167.4]
  wire  _T_3694; // @[MemPrimitives.scala 110:210:@47170.4]
  wire  _T_3695; // @[MemPrimitives.scala 110:228:@47171.4]
  wire  _T_3700; // @[MemPrimitives.scala 110:210:@47174.4]
  wire  _T_3701; // @[MemPrimitives.scala 110:228:@47175.4]
  wire  _T_3706; // @[MemPrimitives.scala 110:210:@47178.4]
  wire  _T_3707; // @[MemPrimitives.scala 110:228:@47179.4]
  wire  _T_3712; // @[MemPrimitives.scala 110:210:@47182.4]
  wire  _T_3713; // @[MemPrimitives.scala 110:228:@47183.4]
  wire  _T_3718; // @[MemPrimitives.scala 110:210:@47186.4]
  wire  _T_3719; // @[MemPrimitives.scala 110:228:@47187.4]
  wire  _T_3724; // @[MemPrimitives.scala 110:210:@47190.4]
  wire  _T_3725; // @[MemPrimitives.scala 110:228:@47191.4]
  wire  _T_3730; // @[MemPrimitives.scala 110:210:@47194.4]
  wire  _T_3731; // @[MemPrimitives.scala 110:228:@47195.4]
  wire  _T_3733; // @[MemPrimitives.scala 123:41:@47215.4]
  wire  _T_3734; // @[MemPrimitives.scala 123:41:@47216.4]
  wire  _T_3735; // @[MemPrimitives.scala 123:41:@47217.4]
  wire  _T_3736; // @[MemPrimitives.scala 123:41:@47218.4]
  wire  _T_3737; // @[MemPrimitives.scala 123:41:@47219.4]
  wire  _T_3738; // @[MemPrimitives.scala 123:41:@47220.4]
  wire  _T_3739; // @[MemPrimitives.scala 123:41:@47221.4]
  wire  _T_3740; // @[MemPrimitives.scala 123:41:@47222.4]
  wire  _T_3741; // @[MemPrimitives.scala 123:41:@47223.4]
  wire  _T_3742; // @[MemPrimitives.scala 123:41:@47224.4]
  wire  _T_3743; // @[MemPrimitives.scala 123:41:@47225.4]
  wire  _T_3744; // @[MemPrimitives.scala 123:41:@47226.4]
  wire  _T_3745; // @[MemPrimitives.scala 123:41:@47227.4]
  wire  _T_3746; // @[MemPrimitives.scala 123:41:@47228.4]
  wire  _T_3747; // @[MemPrimitives.scala 123:41:@47229.4]
  wire [9:0] _T_3749; // @[Cat.scala 30:58:@47231.4]
  wire [9:0] _T_3751; // @[Cat.scala 30:58:@47233.4]
  wire [9:0] _T_3753; // @[Cat.scala 30:58:@47235.4]
  wire [9:0] _T_3755; // @[Cat.scala 30:58:@47237.4]
  wire [9:0] _T_3757; // @[Cat.scala 30:58:@47239.4]
  wire [9:0] _T_3759; // @[Cat.scala 30:58:@47241.4]
  wire [9:0] _T_3761; // @[Cat.scala 30:58:@47243.4]
  wire [9:0] _T_3763; // @[Cat.scala 30:58:@47245.4]
  wire [9:0] _T_3765; // @[Cat.scala 30:58:@47247.4]
  wire [9:0] _T_3767; // @[Cat.scala 30:58:@47249.4]
  wire [9:0] _T_3769; // @[Cat.scala 30:58:@47251.4]
  wire [9:0] _T_3771; // @[Cat.scala 30:58:@47253.4]
  wire [9:0] _T_3773; // @[Cat.scala 30:58:@47255.4]
  wire [9:0] _T_3775; // @[Cat.scala 30:58:@47257.4]
  wire [9:0] _T_3777; // @[Cat.scala 30:58:@47259.4]
  wire [9:0] _T_3778; // @[Mux.scala 31:69:@47260.4]
  wire [9:0] _T_3779; // @[Mux.scala 31:69:@47261.4]
  wire [9:0] _T_3780; // @[Mux.scala 31:69:@47262.4]
  wire [9:0] _T_3781; // @[Mux.scala 31:69:@47263.4]
  wire [9:0] _T_3782; // @[Mux.scala 31:69:@47264.4]
  wire [9:0] _T_3783; // @[Mux.scala 31:69:@47265.4]
  wire [9:0] _T_3784; // @[Mux.scala 31:69:@47266.4]
  wire [9:0] _T_3785; // @[Mux.scala 31:69:@47267.4]
  wire [9:0] _T_3786; // @[Mux.scala 31:69:@47268.4]
  wire [9:0] _T_3787; // @[Mux.scala 31:69:@47269.4]
  wire [9:0] _T_3788; // @[Mux.scala 31:69:@47270.4]
  wire [9:0] _T_3789; // @[Mux.scala 31:69:@47271.4]
  wire [9:0] _T_3790; // @[Mux.scala 31:69:@47272.4]
  wire [9:0] _T_3791; // @[Mux.scala 31:69:@47273.4]
  wire  _T_3798; // @[MemPrimitives.scala 110:210:@47281.4]
  wire  _T_3799; // @[MemPrimitives.scala 110:228:@47282.4]
  wire  _T_3804; // @[MemPrimitives.scala 110:210:@47285.4]
  wire  _T_3805; // @[MemPrimitives.scala 110:228:@47286.4]
  wire  _T_3810; // @[MemPrimitives.scala 110:210:@47289.4]
  wire  _T_3811; // @[MemPrimitives.scala 110:228:@47290.4]
  wire  _T_3816; // @[MemPrimitives.scala 110:210:@47293.4]
  wire  _T_3817; // @[MemPrimitives.scala 110:228:@47294.4]
  wire  _T_3822; // @[MemPrimitives.scala 110:210:@47297.4]
  wire  _T_3823; // @[MemPrimitives.scala 110:228:@47298.4]
  wire  _T_3828; // @[MemPrimitives.scala 110:210:@47301.4]
  wire  _T_3829; // @[MemPrimitives.scala 110:228:@47302.4]
  wire  _T_3834; // @[MemPrimitives.scala 110:210:@47305.4]
  wire  _T_3835; // @[MemPrimitives.scala 110:228:@47306.4]
  wire  _T_3840; // @[MemPrimitives.scala 110:210:@47309.4]
  wire  _T_3841; // @[MemPrimitives.scala 110:228:@47310.4]
  wire  _T_3846; // @[MemPrimitives.scala 110:210:@47313.4]
  wire  _T_3847; // @[MemPrimitives.scala 110:228:@47314.4]
  wire  _T_3852; // @[MemPrimitives.scala 110:210:@47317.4]
  wire  _T_3853; // @[MemPrimitives.scala 110:228:@47318.4]
  wire  _T_3858; // @[MemPrimitives.scala 110:210:@47321.4]
  wire  _T_3859; // @[MemPrimitives.scala 110:228:@47322.4]
  wire  _T_3864; // @[MemPrimitives.scala 110:210:@47325.4]
  wire  _T_3865; // @[MemPrimitives.scala 110:228:@47326.4]
  wire  _T_3870; // @[MemPrimitives.scala 110:210:@47329.4]
  wire  _T_3871; // @[MemPrimitives.scala 110:228:@47330.4]
  wire  _T_3876; // @[MemPrimitives.scala 110:210:@47333.4]
  wire  _T_3877; // @[MemPrimitives.scala 110:228:@47334.4]
  wire  _T_3882; // @[MemPrimitives.scala 110:210:@47337.4]
  wire  _T_3883; // @[MemPrimitives.scala 110:228:@47338.4]
  wire  _T_3885; // @[MemPrimitives.scala 123:41:@47358.4]
  wire  _T_3886; // @[MemPrimitives.scala 123:41:@47359.4]
  wire  _T_3887; // @[MemPrimitives.scala 123:41:@47360.4]
  wire  _T_3888; // @[MemPrimitives.scala 123:41:@47361.4]
  wire  _T_3889; // @[MemPrimitives.scala 123:41:@47362.4]
  wire  _T_3890; // @[MemPrimitives.scala 123:41:@47363.4]
  wire  _T_3891; // @[MemPrimitives.scala 123:41:@47364.4]
  wire  _T_3892; // @[MemPrimitives.scala 123:41:@47365.4]
  wire  _T_3893; // @[MemPrimitives.scala 123:41:@47366.4]
  wire  _T_3894; // @[MemPrimitives.scala 123:41:@47367.4]
  wire  _T_3895; // @[MemPrimitives.scala 123:41:@47368.4]
  wire  _T_3896; // @[MemPrimitives.scala 123:41:@47369.4]
  wire  _T_3897; // @[MemPrimitives.scala 123:41:@47370.4]
  wire  _T_3898; // @[MemPrimitives.scala 123:41:@47371.4]
  wire  _T_3899; // @[MemPrimitives.scala 123:41:@47372.4]
  wire [9:0] _T_3901; // @[Cat.scala 30:58:@47374.4]
  wire [9:0] _T_3903; // @[Cat.scala 30:58:@47376.4]
  wire [9:0] _T_3905; // @[Cat.scala 30:58:@47378.4]
  wire [9:0] _T_3907; // @[Cat.scala 30:58:@47380.4]
  wire [9:0] _T_3909; // @[Cat.scala 30:58:@47382.4]
  wire [9:0] _T_3911; // @[Cat.scala 30:58:@47384.4]
  wire [9:0] _T_3913; // @[Cat.scala 30:58:@47386.4]
  wire [9:0] _T_3915; // @[Cat.scala 30:58:@47388.4]
  wire [9:0] _T_3917; // @[Cat.scala 30:58:@47390.4]
  wire [9:0] _T_3919; // @[Cat.scala 30:58:@47392.4]
  wire [9:0] _T_3921; // @[Cat.scala 30:58:@47394.4]
  wire [9:0] _T_3923; // @[Cat.scala 30:58:@47396.4]
  wire [9:0] _T_3925; // @[Cat.scala 30:58:@47398.4]
  wire [9:0] _T_3927; // @[Cat.scala 30:58:@47400.4]
  wire [9:0] _T_3929; // @[Cat.scala 30:58:@47402.4]
  wire [9:0] _T_3930; // @[Mux.scala 31:69:@47403.4]
  wire [9:0] _T_3931; // @[Mux.scala 31:69:@47404.4]
  wire [9:0] _T_3932; // @[Mux.scala 31:69:@47405.4]
  wire [9:0] _T_3933; // @[Mux.scala 31:69:@47406.4]
  wire [9:0] _T_3934; // @[Mux.scala 31:69:@47407.4]
  wire [9:0] _T_3935; // @[Mux.scala 31:69:@47408.4]
  wire [9:0] _T_3936; // @[Mux.scala 31:69:@47409.4]
  wire [9:0] _T_3937; // @[Mux.scala 31:69:@47410.4]
  wire [9:0] _T_3938; // @[Mux.scala 31:69:@47411.4]
  wire [9:0] _T_3939; // @[Mux.scala 31:69:@47412.4]
  wire [9:0] _T_3940; // @[Mux.scala 31:69:@47413.4]
  wire [9:0] _T_3941; // @[Mux.scala 31:69:@47414.4]
  wire [9:0] _T_3942; // @[Mux.scala 31:69:@47415.4]
  wire [9:0] _T_3943; // @[Mux.scala 31:69:@47416.4]
  wire  _T_3950; // @[MemPrimitives.scala 110:210:@47424.4]
  wire  _T_3951; // @[MemPrimitives.scala 110:228:@47425.4]
  wire  _T_3956; // @[MemPrimitives.scala 110:210:@47428.4]
  wire  _T_3957; // @[MemPrimitives.scala 110:228:@47429.4]
  wire  _T_3962; // @[MemPrimitives.scala 110:210:@47432.4]
  wire  _T_3963; // @[MemPrimitives.scala 110:228:@47433.4]
  wire  _T_3968; // @[MemPrimitives.scala 110:210:@47436.4]
  wire  _T_3969; // @[MemPrimitives.scala 110:228:@47437.4]
  wire  _T_3974; // @[MemPrimitives.scala 110:210:@47440.4]
  wire  _T_3975; // @[MemPrimitives.scala 110:228:@47441.4]
  wire  _T_3980; // @[MemPrimitives.scala 110:210:@47444.4]
  wire  _T_3981; // @[MemPrimitives.scala 110:228:@47445.4]
  wire  _T_3986; // @[MemPrimitives.scala 110:210:@47448.4]
  wire  _T_3987; // @[MemPrimitives.scala 110:228:@47449.4]
  wire  _T_3992; // @[MemPrimitives.scala 110:210:@47452.4]
  wire  _T_3993; // @[MemPrimitives.scala 110:228:@47453.4]
  wire  _T_3998; // @[MemPrimitives.scala 110:210:@47456.4]
  wire  _T_3999; // @[MemPrimitives.scala 110:228:@47457.4]
  wire  _T_4004; // @[MemPrimitives.scala 110:210:@47460.4]
  wire  _T_4005; // @[MemPrimitives.scala 110:228:@47461.4]
  wire  _T_4010; // @[MemPrimitives.scala 110:210:@47464.4]
  wire  _T_4011; // @[MemPrimitives.scala 110:228:@47465.4]
  wire  _T_4016; // @[MemPrimitives.scala 110:210:@47468.4]
  wire  _T_4017; // @[MemPrimitives.scala 110:228:@47469.4]
  wire  _T_4022; // @[MemPrimitives.scala 110:210:@47472.4]
  wire  _T_4023; // @[MemPrimitives.scala 110:228:@47473.4]
  wire  _T_4028; // @[MemPrimitives.scala 110:210:@47476.4]
  wire  _T_4029; // @[MemPrimitives.scala 110:228:@47477.4]
  wire  _T_4034; // @[MemPrimitives.scala 110:210:@47480.4]
  wire  _T_4035; // @[MemPrimitives.scala 110:228:@47481.4]
  wire  _T_4037; // @[MemPrimitives.scala 123:41:@47501.4]
  wire  _T_4038; // @[MemPrimitives.scala 123:41:@47502.4]
  wire  _T_4039; // @[MemPrimitives.scala 123:41:@47503.4]
  wire  _T_4040; // @[MemPrimitives.scala 123:41:@47504.4]
  wire  _T_4041; // @[MemPrimitives.scala 123:41:@47505.4]
  wire  _T_4042; // @[MemPrimitives.scala 123:41:@47506.4]
  wire  _T_4043; // @[MemPrimitives.scala 123:41:@47507.4]
  wire  _T_4044; // @[MemPrimitives.scala 123:41:@47508.4]
  wire  _T_4045; // @[MemPrimitives.scala 123:41:@47509.4]
  wire  _T_4046; // @[MemPrimitives.scala 123:41:@47510.4]
  wire  _T_4047; // @[MemPrimitives.scala 123:41:@47511.4]
  wire  _T_4048; // @[MemPrimitives.scala 123:41:@47512.4]
  wire  _T_4049; // @[MemPrimitives.scala 123:41:@47513.4]
  wire  _T_4050; // @[MemPrimitives.scala 123:41:@47514.4]
  wire  _T_4051; // @[MemPrimitives.scala 123:41:@47515.4]
  wire [9:0] _T_4053; // @[Cat.scala 30:58:@47517.4]
  wire [9:0] _T_4055; // @[Cat.scala 30:58:@47519.4]
  wire [9:0] _T_4057; // @[Cat.scala 30:58:@47521.4]
  wire [9:0] _T_4059; // @[Cat.scala 30:58:@47523.4]
  wire [9:0] _T_4061; // @[Cat.scala 30:58:@47525.4]
  wire [9:0] _T_4063; // @[Cat.scala 30:58:@47527.4]
  wire [9:0] _T_4065; // @[Cat.scala 30:58:@47529.4]
  wire [9:0] _T_4067; // @[Cat.scala 30:58:@47531.4]
  wire [9:0] _T_4069; // @[Cat.scala 30:58:@47533.4]
  wire [9:0] _T_4071; // @[Cat.scala 30:58:@47535.4]
  wire [9:0] _T_4073; // @[Cat.scala 30:58:@47537.4]
  wire [9:0] _T_4075; // @[Cat.scala 30:58:@47539.4]
  wire [9:0] _T_4077; // @[Cat.scala 30:58:@47541.4]
  wire [9:0] _T_4079; // @[Cat.scala 30:58:@47543.4]
  wire [9:0] _T_4081; // @[Cat.scala 30:58:@47545.4]
  wire [9:0] _T_4082; // @[Mux.scala 31:69:@47546.4]
  wire [9:0] _T_4083; // @[Mux.scala 31:69:@47547.4]
  wire [9:0] _T_4084; // @[Mux.scala 31:69:@47548.4]
  wire [9:0] _T_4085; // @[Mux.scala 31:69:@47549.4]
  wire [9:0] _T_4086; // @[Mux.scala 31:69:@47550.4]
  wire [9:0] _T_4087; // @[Mux.scala 31:69:@47551.4]
  wire [9:0] _T_4088; // @[Mux.scala 31:69:@47552.4]
  wire [9:0] _T_4089; // @[Mux.scala 31:69:@47553.4]
  wire [9:0] _T_4090; // @[Mux.scala 31:69:@47554.4]
  wire [9:0] _T_4091; // @[Mux.scala 31:69:@47555.4]
  wire [9:0] _T_4092; // @[Mux.scala 31:69:@47556.4]
  wire [9:0] _T_4093; // @[Mux.scala 31:69:@47557.4]
  wire [9:0] _T_4094; // @[Mux.scala 31:69:@47558.4]
  wire [9:0] _T_4095; // @[Mux.scala 31:69:@47559.4]
  wire  _T_4102; // @[MemPrimitives.scala 110:210:@47567.4]
  wire  _T_4103; // @[MemPrimitives.scala 110:228:@47568.4]
  wire  _T_4108; // @[MemPrimitives.scala 110:210:@47571.4]
  wire  _T_4109; // @[MemPrimitives.scala 110:228:@47572.4]
  wire  _T_4114; // @[MemPrimitives.scala 110:210:@47575.4]
  wire  _T_4115; // @[MemPrimitives.scala 110:228:@47576.4]
  wire  _T_4120; // @[MemPrimitives.scala 110:210:@47579.4]
  wire  _T_4121; // @[MemPrimitives.scala 110:228:@47580.4]
  wire  _T_4126; // @[MemPrimitives.scala 110:210:@47583.4]
  wire  _T_4127; // @[MemPrimitives.scala 110:228:@47584.4]
  wire  _T_4132; // @[MemPrimitives.scala 110:210:@47587.4]
  wire  _T_4133; // @[MemPrimitives.scala 110:228:@47588.4]
  wire  _T_4138; // @[MemPrimitives.scala 110:210:@47591.4]
  wire  _T_4139; // @[MemPrimitives.scala 110:228:@47592.4]
  wire  _T_4144; // @[MemPrimitives.scala 110:210:@47595.4]
  wire  _T_4145; // @[MemPrimitives.scala 110:228:@47596.4]
  wire  _T_4150; // @[MemPrimitives.scala 110:210:@47599.4]
  wire  _T_4151; // @[MemPrimitives.scala 110:228:@47600.4]
  wire  _T_4156; // @[MemPrimitives.scala 110:210:@47603.4]
  wire  _T_4157; // @[MemPrimitives.scala 110:228:@47604.4]
  wire  _T_4162; // @[MemPrimitives.scala 110:210:@47607.4]
  wire  _T_4163; // @[MemPrimitives.scala 110:228:@47608.4]
  wire  _T_4168; // @[MemPrimitives.scala 110:210:@47611.4]
  wire  _T_4169; // @[MemPrimitives.scala 110:228:@47612.4]
  wire  _T_4174; // @[MemPrimitives.scala 110:210:@47615.4]
  wire  _T_4175; // @[MemPrimitives.scala 110:228:@47616.4]
  wire  _T_4180; // @[MemPrimitives.scala 110:210:@47619.4]
  wire  _T_4181; // @[MemPrimitives.scala 110:228:@47620.4]
  wire  _T_4186; // @[MemPrimitives.scala 110:210:@47623.4]
  wire  _T_4187; // @[MemPrimitives.scala 110:228:@47624.4]
  wire  _T_4189; // @[MemPrimitives.scala 123:41:@47644.4]
  wire  _T_4190; // @[MemPrimitives.scala 123:41:@47645.4]
  wire  _T_4191; // @[MemPrimitives.scala 123:41:@47646.4]
  wire  _T_4192; // @[MemPrimitives.scala 123:41:@47647.4]
  wire  _T_4193; // @[MemPrimitives.scala 123:41:@47648.4]
  wire  _T_4194; // @[MemPrimitives.scala 123:41:@47649.4]
  wire  _T_4195; // @[MemPrimitives.scala 123:41:@47650.4]
  wire  _T_4196; // @[MemPrimitives.scala 123:41:@47651.4]
  wire  _T_4197; // @[MemPrimitives.scala 123:41:@47652.4]
  wire  _T_4198; // @[MemPrimitives.scala 123:41:@47653.4]
  wire  _T_4199; // @[MemPrimitives.scala 123:41:@47654.4]
  wire  _T_4200; // @[MemPrimitives.scala 123:41:@47655.4]
  wire  _T_4201; // @[MemPrimitives.scala 123:41:@47656.4]
  wire  _T_4202; // @[MemPrimitives.scala 123:41:@47657.4]
  wire  _T_4203; // @[MemPrimitives.scala 123:41:@47658.4]
  wire [9:0] _T_4205; // @[Cat.scala 30:58:@47660.4]
  wire [9:0] _T_4207; // @[Cat.scala 30:58:@47662.4]
  wire [9:0] _T_4209; // @[Cat.scala 30:58:@47664.4]
  wire [9:0] _T_4211; // @[Cat.scala 30:58:@47666.4]
  wire [9:0] _T_4213; // @[Cat.scala 30:58:@47668.4]
  wire [9:0] _T_4215; // @[Cat.scala 30:58:@47670.4]
  wire [9:0] _T_4217; // @[Cat.scala 30:58:@47672.4]
  wire [9:0] _T_4219; // @[Cat.scala 30:58:@47674.4]
  wire [9:0] _T_4221; // @[Cat.scala 30:58:@47676.4]
  wire [9:0] _T_4223; // @[Cat.scala 30:58:@47678.4]
  wire [9:0] _T_4225; // @[Cat.scala 30:58:@47680.4]
  wire [9:0] _T_4227; // @[Cat.scala 30:58:@47682.4]
  wire [9:0] _T_4229; // @[Cat.scala 30:58:@47684.4]
  wire [9:0] _T_4231; // @[Cat.scala 30:58:@47686.4]
  wire [9:0] _T_4233; // @[Cat.scala 30:58:@47688.4]
  wire [9:0] _T_4234; // @[Mux.scala 31:69:@47689.4]
  wire [9:0] _T_4235; // @[Mux.scala 31:69:@47690.4]
  wire [9:0] _T_4236; // @[Mux.scala 31:69:@47691.4]
  wire [9:0] _T_4237; // @[Mux.scala 31:69:@47692.4]
  wire [9:0] _T_4238; // @[Mux.scala 31:69:@47693.4]
  wire [9:0] _T_4239; // @[Mux.scala 31:69:@47694.4]
  wire [9:0] _T_4240; // @[Mux.scala 31:69:@47695.4]
  wire [9:0] _T_4241; // @[Mux.scala 31:69:@47696.4]
  wire [9:0] _T_4242; // @[Mux.scala 31:69:@47697.4]
  wire [9:0] _T_4243; // @[Mux.scala 31:69:@47698.4]
  wire [9:0] _T_4244; // @[Mux.scala 31:69:@47699.4]
  wire [9:0] _T_4245; // @[Mux.scala 31:69:@47700.4]
  wire [9:0] _T_4246; // @[Mux.scala 31:69:@47701.4]
  wire [9:0] _T_4247; // @[Mux.scala 31:69:@47702.4]
  wire  _T_4252; // @[MemPrimitives.scala 110:210:@47709.4]
  wire  _T_4255; // @[MemPrimitives.scala 110:228:@47711.4]
  wire  _T_4258; // @[MemPrimitives.scala 110:210:@47713.4]
  wire  _T_4261; // @[MemPrimitives.scala 110:228:@47715.4]
  wire  _T_4264; // @[MemPrimitives.scala 110:210:@47717.4]
  wire  _T_4267; // @[MemPrimitives.scala 110:228:@47719.4]
  wire  _T_4270; // @[MemPrimitives.scala 110:210:@47721.4]
  wire  _T_4273; // @[MemPrimitives.scala 110:228:@47723.4]
  wire  _T_4276; // @[MemPrimitives.scala 110:210:@47725.4]
  wire  _T_4279; // @[MemPrimitives.scala 110:228:@47727.4]
  wire  _T_4282; // @[MemPrimitives.scala 110:210:@47729.4]
  wire  _T_4285; // @[MemPrimitives.scala 110:228:@47731.4]
  wire  _T_4288; // @[MemPrimitives.scala 110:210:@47733.4]
  wire  _T_4291; // @[MemPrimitives.scala 110:228:@47735.4]
  wire  _T_4294; // @[MemPrimitives.scala 110:210:@47737.4]
  wire  _T_4297; // @[MemPrimitives.scala 110:228:@47739.4]
  wire  _T_4300; // @[MemPrimitives.scala 110:210:@47741.4]
  wire  _T_4303; // @[MemPrimitives.scala 110:228:@47743.4]
  wire  _T_4306; // @[MemPrimitives.scala 110:210:@47745.4]
  wire  _T_4309; // @[MemPrimitives.scala 110:228:@47747.4]
  wire  _T_4312; // @[MemPrimitives.scala 110:210:@47749.4]
  wire  _T_4315; // @[MemPrimitives.scala 110:228:@47751.4]
  wire  _T_4318; // @[MemPrimitives.scala 110:210:@47753.4]
  wire  _T_4321; // @[MemPrimitives.scala 110:228:@47755.4]
  wire  _T_4324; // @[MemPrimitives.scala 110:210:@47757.4]
  wire  _T_4327; // @[MemPrimitives.scala 110:228:@47759.4]
  wire  _T_4330; // @[MemPrimitives.scala 110:210:@47761.4]
  wire  _T_4333; // @[MemPrimitives.scala 110:228:@47763.4]
  wire  _T_4336; // @[MemPrimitives.scala 110:210:@47765.4]
  wire  _T_4339; // @[MemPrimitives.scala 110:228:@47767.4]
  wire  _T_4341; // @[MemPrimitives.scala 123:41:@47787.4]
  wire  _T_4342; // @[MemPrimitives.scala 123:41:@47788.4]
  wire  _T_4343; // @[MemPrimitives.scala 123:41:@47789.4]
  wire  _T_4344; // @[MemPrimitives.scala 123:41:@47790.4]
  wire  _T_4345; // @[MemPrimitives.scala 123:41:@47791.4]
  wire  _T_4346; // @[MemPrimitives.scala 123:41:@47792.4]
  wire  _T_4347; // @[MemPrimitives.scala 123:41:@47793.4]
  wire  _T_4348; // @[MemPrimitives.scala 123:41:@47794.4]
  wire  _T_4349; // @[MemPrimitives.scala 123:41:@47795.4]
  wire  _T_4350; // @[MemPrimitives.scala 123:41:@47796.4]
  wire  _T_4351; // @[MemPrimitives.scala 123:41:@47797.4]
  wire  _T_4352; // @[MemPrimitives.scala 123:41:@47798.4]
  wire  _T_4353; // @[MemPrimitives.scala 123:41:@47799.4]
  wire  _T_4354; // @[MemPrimitives.scala 123:41:@47800.4]
  wire  _T_4355; // @[MemPrimitives.scala 123:41:@47801.4]
  wire [9:0] _T_4357; // @[Cat.scala 30:58:@47803.4]
  wire [9:0] _T_4359; // @[Cat.scala 30:58:@47805.4]
  wire [9:0] _T_4361; // @[Cat.scala 30:58:@47807.4]
  wire [9:0] _T_4363; // @[Cat.scala 30:58:@47809.4]
  wire [9:0] _T_4365; // @[Cat.scala 30:58:@47811.4]
  wire [9:0] _T_4367; // @[Cat.scala 30:58:@47813.4]
  wire [9:0] _T_4369; // @[Cat.scala 30:58:@47815.4]
  wire [9:0] _T_4371; // @[Cat.scala 30:58:@47817.4]
  wire [9:0] _T_4373; // @[Cat.scala 30:58:@47819.4]
  wire [9:0] _T_4375; // @[Cat.scala 30:58:@47821.4]
  wire [9:0] _T_4377; // @[Cat.scala 30:58:@47823.4]
  wire [9:0] _T_4379; // @[Cat.scala 30:58:@47825.4]
  wire [9:0] _T_4381; // @[Cat.scala 30:58:@47827.4]
  wire [9:0] _T_4383; // @[Cat.scala 30:58:@47829.4]
  wire [9:0] _T_4385; // @[Cat.scala 30:58:@47831.4]
  wire [9:0] _T_4386; // @[Mux.scala 31:69:@47832.4]
  wire [9:0] _T_4387; // @[Mux.scala 31:69:@47833.4]
  wire [9:0] _T_4388; // @[Mux.scala 31:69:@47834.4]
  wire [9:0] _T_4389; // @[Mux.scala 31:69:@47835.4]
  wire [9:0] _T_4390; // @[Mux.scala 31:69:@47836.4]
  wire [9:0] _T_4391; // @[Mux.scala 31:69:@47837.4]
  wire [9:0] _T_4392; // @[Mux.scala 31:69:@47838.4]
  wire [9:0] _T_4393; // @[Mux.scala 31:69:@47839.4]
  wire [9:0] _T_4394; // @[Mux.scala 31:69:@47840.4]
  wire [9:0] _T_4395; // @[Mux.scala 31:69:@47841.4]
  wire [9:0] _T_4396; // @[Mux.scala 31:69:@47842.4]
  wire [9:0] _T_4397; // @[Mux.scala 31:69:@47843.4]
  wire [9:0] _T_4398; // @[Mux.scala 31:69:@47844.4]
  wire [9:0] _T_4399; // @[Mux.scala 31:69:@47845.4]
  wire  _T_4404; // @[MemPrimitives.scala 110:210:@47852.4]
  wire  _T_4407; // @[MemPrimitives.scala 110:228:@47854.4]
  wire  _T_4410; // @[MemPrimitives.scala 110:210:@47856.4]
  wire  _T_4413; // @[MemPrimitives.scala 110:228:@47858.4]
  wire  _T_4416; // @[MemPrimitives.scala 110:210:@47860.4]
  wire  _T_4419; // @[MemPrimitives.scala 110:228:@47862.4]
  wire  _T_4422; // @[MemPrimitives.scala 110:210:@47864.4]
  wire  _T_4425; // @[MemPrimitives.scala 110:228:@47866.4]
  wire  _T_4428; // @[MemPrimitives.scala 110:210:@47868.4]
  wire  _T_4431; // @[MemPrimitives.scala 110:228:@47870.4]
  wire  _T_4434; // @[MemPrimitives.scala 110:210:@47872.4]
  wire  _T_4437; // @[MemPrimitives.scala 110:228:@47874.4]
  wire  _T_4440; // @[MemPrimitives.scala 110:210:@47876.4]
  wire  _T_4443; // @[MemPrimitives.scala 110:228:@47878.4]
  wire  _T_4446; // @[MemPrimitives.scala 110:210:@47880.4]
  wire  _T_4449; // @[MemPrimitives.scala 110:228:@47882.4]
  wire  _T_4452; // @[MemPrimitives.scala 110:210:@47884.4]
  wire  _T_4455; // @[MemPrimitives.scala 110:228:@47886.4]
  wire  _T_4458; // @[MemPrimitives.scala 110:210:@47888.4]
  wire  _T_4461; // @[MemPrimitives.scala 110:228:@47890.4]
  wire  _T_4464; // @[MemPrimitives.scala 110:210:@47892.4]
  wire  _T_4467; // @[MemPrimitives.scala 110:228:@47894.4]
  wire  _T_4470; // @[MemPrimitives.scala 110:210:@47896.4]
  wire  _T_4473; // @[MemPrimitives.scala 110:228:@47898.4]
  wire  _T_4476; // @[MemPrimitives.scala 110:210:@47900.4]
  wire  _T_4479; // @[MemPrimitives.scala 110:228:@47902.4]
  wire  _T_4482; // @[MemPrimitives.scala 110:210:@47904.4]
  wire  _T_4485; // @[MemPrimitives.scala 110:228:@47906.4]
  wire  _T_4488; // @[MemPrimitives.scala 110:210:@47908.4]
  wire  _T_4491; // @[MemPrimitives.scala 110:228:@47910.4]
  wire  _T_4493; // @[MemPrimitives.scala 123:41:@47930.4]
  wire  _T_4494; // @[MemPrimitives.scala 123:41:@47931.4]
  wire  _T_4495; // @[MemPrimitives.scala 123:41:@47932.4]
  wire  _T_4496; // @[MemPrimitives.scala 123:41:@47933.4]
  wire  _T_4497; // @[MemPrimitives.scala 123:41:@47934.4]
  wire  _T_4498; // @[MemPrimitives.scala 123:41:@47935.4]
  wire  _T_4499; // @[MemPrimitives.scala 123:41:@47936.4]
  wire  _T_4500; // @[MemPrimitives.scala 123:41:@47937.4]
  wire  _T_4501; // @[MemPrimitives.scala 123:41:@47938.4]
  wire  _T_4502; // @[MemPrimitives.scala 123:41:@47939.4]
  wire  _T_4503; // @[MemPrimitives.scala 123:41:@47940.4]
  wire  _T_4504; // @[MemPrimitives.scala 123:41:@47941.4]
  wire  _T_4505; // @[MemPrimitives.scala 123:41:@47942.4]
  wire  _T_4506; // @[MemPrimitives.scala 123:41:@47943.4]
  wire  _T_4507; // @[MemPrimitives.scala 123:41:@47944.4]
  wire [9:0] _T_4509; // @[Cat.scala 30:58:@47946.4]
  wire [9:0] _T_4511; // @[Cat.scala 30:58:@47948.4]
  wire [9:0] _T_4513; // @[Cat.scala 30:58:@47950.4]
  wire [9:0] _T_4515; // @[Cat.scala 30:58:@47952.4]
  wire [9:0] _T_4517; // @[Cat.scala 30:58:@47954.4]
  wire [9:0] _T_4519; // @[Cat.scala 30:58:@47956.4]
  wire [9:0] _T_4521; // @[Cat.scala 30:58:@47958.4]
  wire [9:0] _T_4523; // @[Cat.scala 30:58:@47960.4]
  wire [9:0] _T_4525; // @[Cat.scala 30:58:@47962.4]
  wire [9:0] _T_4527; // @[Cat.scala 30:58:@47964.4]
  wire [9:0] _T_4529; // @[Cat.scala 30:58:@47966.4]
  wire [9:0] _T_4531; // @[Cat.scala 30:58:@47968.4]
  wire [9:0] _T_4533; // @[Cat.scala 30:58:@47970.4]
  wire [9:0] _T_4535; // @[Cat.scala 30:58:@47972.4]
  wire [9:0] _T_4537; // @[Cat.scala 30:58:@47974.4]
  wire [9:0] _T_4538; // @[Mux.scala 31:69:@47975.4]
  wire [9:0] _T_4539; // @[Mux.scala 31:69:@47976.4]
  wire [9:0] _T_4540; // @[Mux.scala 31:69:@47977.4]
  wire [9:0] _T_4541; // @[Mux.scala 31:69:@47978.4]
  wire [9:0] _T_4542; // @[Mux.scala 31:69:@47979.4]
  wire [9:0] _T_4543; // @[Mux.scala 31:69:@47980.4]
  wire [9:0] _T_4544; // @[Mux.scala 31:69:@47981.4]
  wire [9:0] _T_4545; // @[Mux.scala 31:69:@47982.4]
  wire [9:0] _T_4546; // @[Mux.scala 31:69:@47983.4]
  wire [9:0] _T_4547; // @[Mux.scala 31:69:@47984.4]
  wire [9:0] _T_4548; // @[Mux.scala 31:69:@47985.4]
  wire [9:0] _T_4549; // @[Mux.scala 31:69:@47986.4]
  wire [9:0] _T_4550; // @[Mux.scala 31:69:@47987.4]
  wire [9:0] _T_4551; // @[Mux.scala 31:69:@47988.4]
  wire  _T_4559; // @[MemPrimitives.scala 110:228:@47997.4]
  wire  _T_4565; // @[MemPrimitives.scala 110:228:@48001.4]
  wire  _T_4571; // @[MemPrimitives.scala 110:228:@48005.4]
  wire  _T_4577; // @[MemPrimitives.scala 110:228:@48009.4]
  wire  _T_4583; // @[MemPrimitives.scala 110:228:@48013.4]
  wire  _T_4589; // @[MemPrimitives.scala 110:228:@48017.4]
  wire  _T_4595; // @[MemPrimitives.scala 110:228:@48021.4]
  wire  _T_4601; // @[MemPrimitives.scala 110:228:@48025.4]
  wire  _T_4607; // @[MemPrimitives.scala 110:228:@48029.4]
  wire  _T_4613; // @[MemPrimitives.scala 110:228:@48033.4]
  wire  _T_4619; // @[MemPrimitives.scala 110:228:@48037.4]
  wire  _T_4625; // @[MemPrimitives.scala 110:228:@48041.4]
  wire  _T_4631; // @[MemPrimitives.scala 110:228:@48045.4]
  wire  _T_4637; // @[MemPrimitives.scala 110:228:@48049.4]
  wire  _T_4643; // @[MemPrimitives.scala 110:228:@48053.4]
  wire  _T_4645; // @[MemPrimitives.scala 123:41:@48073.4]
  wire  _T_4646; // @[MemPrimitives.scala 123:41:@48074.4]
  wire  _T_4647; // @[MemPrimitives.scala 123:41:@48075.4]
  wire  _T_4648; // @[MemPrimitives.scala 123:41:@48076.4]
  wire  _T_4649; // @[MemPrimitives.scala 123:41:@48077.4]
  wire  _T_4650; // @[MemPrimitives.scala 123:41:@48078.4]
  wire  _T_4651; // @[MemPrimitives.scala 123:41:@48079.4]
  wire  _T_4652; // @[MemPrimitives.scala 123:41:@48080.4]
  wire  _T_4653; // @[MemPrimitives.scala 123:41:@48081.4]
  wire  _T_4654; // @[MemPrimitives.scala 123:41:@48082.4]
  wire  _T_4655; // @[MemPrimitives.scala 123:41:@48083.4]
  wire  _T_4656; // @[MemPrimitives.scala 123:41:@48084.4]
  wire  _T_4657; // @[MemPrimitives.scala 123:41:@48085.4]
  wire  _T_4658; // @[MemPrimitives.scala 123:41:@48086.4]
  wire  _T_4659; // @[MemPrimitives.scala 123:41:@48087.4]
  wire [9:0] _T_4661; // @[Cat.scala 30:58:@48089.4]
  wire [9:0] _T_4663; // @[Cat.scala 30:58:@48091.4]
  wire [9:0] _T_4665; // @[Cat.scala 30:58:@48093.4]
  wire [9:0] _T_4667; // @[Cat.scala 30:58:@48095.4]
  wire [9:0] _T_4669; // @[Cat.scala 30:58:@48097.4]
  wire [9:0] _T_4671; // @[Cat.scala 30:58:@48099.4]
  wire [9:0] _T_4673; // @[Cat.scala 30:58:@48101.4]
  wire [9:0] _T_4675; // @[Cat.scala 30:58:@48103.4]
  wire [9:0] _T_4677; // @[Cat.scala 30:58:@48105.4]
  wire [9:0] _T_4679; // @[Cat.scala 30:58:@48107.4]
  wire [9:0] _T_4681; // @[Cat.scala 30:58:@48109.4]
  wire [9:0] _T_4683; // @[Cat.scala 30:58:@48111.4]
  wire [9:0] _T_4685; // @[Cat.scala 30:58:@48113.4]
  wire [9:0] _T_4687; // @[Cat.scala 30:58:@48115.4]
  wire [9:0] _T_4689; // @[Cat.scala 30:58:@48117.4]
  wire [9:0] _T_4690; // @[Mux.scala 31:69:@48118.4]
  wire [9:0] _T_4691; // @[Mux.scala 31:69:@48119.4]
  wire [9:0] _T_4692; // @[Mux.scala 31:69:@48120.4]
  wire [9:0] _T_4693; // @[Mux.scala 31:69:@48121.4]
  wire [9:0] _T_4694; // @[Mux.scala 31:69:@48122.4]
  wire [9:0] _T_4695; // @[Mux.scala 31:69:@48123.4]
  wire [9:0] _T_4696; // @[Mux.scala 31:69:@48124.4]
  wire [9:0] _T_4697; // @[Mux.scala 31:69:@48125.4]
  wire [9:0] _T_4698; // @[Mux.scala 31:69:@48126.4]
  wire [9:0] _T_4699; // @[Mux.scala 31:69:@48127.4]
  wire [9:0] _T_4700; // @[Mux.scala 31:69:@48128.4]
  wire [9:0] _T_4701; // @[Mux.scala 31:69:@48129.4]
  wire [9:0] _T_4702; // @[Mux.scala 31:69:@48130.4]
  wire [9:0] _T_4703; // @[Mux.scala 31:69:@48131.4]
  wire  _T_4711; // @[MemPrimitives.scala 110:228:@48140.4]
  wire  _T_4717; // @[MemPrimitives.scala 110:228:@48144.4]
  wire  _T_4723; // @[MemPrimitives.scala 110:228:@48148.4]
  wire  _T_4729; // @[MemPrimitives.scala 110:228:@48152.4]
  wire  _T_4735; // @[MemPrimitives.scala 110:228:@48156.4]
  wire  _T_4741; // @[MemPrimitives.scala 110:228:@48160.4]
  wire  _T_4747; // @[MemPrimitives.scala 110:228:@48164.4]
  wire  _T_4753; // @[MemPrimitives.scala 110:228:@48168.4]
  wire  _T_4759; // @[MemPrimitives.scala 110:228:@48172.4]
  wire  _T_4765; // @[MemPrimitives.scala 110:228:@48176.4]
  wire  _T_4771; // @[MemPrimitives.scala 110:228:@48180.4]
  wire  _T_4777; // @[MemPrimitives.scala 110:228:@48184.4]
  wire  _T_4783; // @[MemPrimitives.scala 110:228:@48188.4]
  wire  _T_4789; // @[MemPrimitives.scala 110:228:@48192.4]
  wire  _T_4795; // @[MemPrimitives.scala 110:228:@48196.4]
  wire  _T_4797; // @[MemPrimitives.scala 123:41:@48216.4]
  wire  _T_4798; // @[MemPrimitives.scala 123:41:@48217.4]
  wire  _T_4799; // @[MemPrimitives.scala 123:41:@48218.4]
  wire  _T_4800; // @[MemPrimitives.scala 123:41:@48219.4]
  wire  _T_4801; // @[MemPrimitives.scala 123:41:@48220.4]
  wire  _T_4802; // @[MemPrimitives.scala 123:41:@48221.4]
  wire  _T_4803; // @[MemPrimitives.scala 123:41:@48222.4]
  wire  _T_4804; // @[MemPrimitives.scala 123:41:@48223.4]
  wire  _T_4805; // @[MemPrimitives.scala 123:41:@48224.4]
  wire  _T_4806; // @[MemPrimitives.scala 123:41:@48225.4]
  wire  _T_4807; // @[MemPrimitives.scala 123:41:@48226.4]
  wire  _T_4808; // @[MemPrimitives.scala 123:41:@48227.4]
  wire  _T_4809; // @[MemPrimitives.scala 123:41:@48228.4]
  wire  _T_4810; // @[MemPrimitives.scala 123:41:@48229.4]
  wire  _T_4811; // @[MemPrimitives.scala 123:41:@48230.4]
  wire [9:0] _T_4813; // @[Cat.scala 30:58:@48232.4]
  wire [9:0] _T_4815; // @[Cat.scala 30:58:@48234.4]
  wire [9:0] _T_4817; // @[Cat.scala 30:58:@48236.4]
  wire [9:0] _T_4819; // @[Cat.scala 30:58:@48238.4]
  wire [9:0] _T_4821; // @[Cat.scala 30:58:@48240.4]
  wire [9:0] _T_4823; // @[Cat.scala 30:58:@48242.4]
  wire [9:0] _T_4825; // @[Cat.scala 30:58:@48244.4]
  wire [9:0] _T_4827; // @[Cat.scala 30:58:@48246.4]
  wire [9:0] _T_4829; // @[Cat.scala 30:58:@48248.4]
  wire [9:0] _T_4831; // @[Cat.scala 30:58:@48250.4]
  wire [9:0] _T_4833; // @[Cat.scala 30:58:@48252.4]
  wire [9:0] _T_4835; // @[Cat.scala 30:58:@48254.4]
  wire [9:0] _T_4837; // @[Cat.scala 30:58:@48256.4]
  wire [9:0] _T_4839; // @[Cat.scala 30:58:@48258.4]
  wire [9:0] _T_4841; // @[Cat.scala 30:58:@48260.4]
  wire [9:0] _T_4842; // @[Mux.scala 31:69:@48261.4]
  wire [9:0] _T_4843; // @[Mux.scala 31:69:@48262.4]
  wire [9:0] _T_4844; // @[Mux.scala 31:69:@48263.4]
  wire [9:0] _T_4845; // @[Mux.scala 31:69:@48264.4]
  wire [9:0] _T_4846; // @[Mux.scala 31:69:@48265.4]
  wire [9:0] _T_4847; // @[Mux.scala 31:69:@48266.4]
  wire [9:0] _T_4848; // @[Mux.scala 31:69:@48267.4]
  wire [9:0] _T_4849; // @[Mux.scala 31:69:@48268.4]
  wire [9:0] _T_4850; // @[Mux.scala 31:69:@48269.4]
  wire [9:0] _T_4851; // @[Mux.scala 31:69:@48270.4]
  wire [9:0] _T_4852; // @[Mux.scala 31:69:@48271.4]
  wire [9:0] _T_4853; // @[Mux.scala 31:69:@48272.4]
  wire [9:0] _T_4854; // @[Mux.scala 31:69:@48273.4]
  wire [9:0] _T_4855; // @[Mux.scala 31:69:@48274.4]
  wire  _T_4863; // @[MemPrimitives.scala 110:228:@48283.4]
  wire  _T_4869; // @[MemPrimitives.scala 110:228:@48287.4]
  wire  _T_4875; // @[MemPrimitives.scala 110:228:@48291.4]
  wire  _T_4881; // @[MemPrimitives.scala 110:228:@48295.4]
  wire  _T_4887; // @[MemPrimitives.scala 110:228:@48299.4]
  wire  _T_4893; // @[MemPrimitives.scala 110:228:@48303.4]
  wire  _T_4899; // @[MemPrimitives.scala 110:228:@48307.4]
  wire  _T_4905; // @[MemPrimitives.scala 110:228:@48311.4]
  wire  _T_4911; // @[MemPrimitives.scala 110:228:@48315.4]
  wire  _T_4917; // @[MemPrimitives.scala 110:228:@48319.4]
  wire  _T_4923; // @[MemPrimitives.scala 110:228:@48323.4]
  wire  _T_4929; // @[MemPrimitives.scala 110:228:@48327.4]
  wire  _T_4935; // @[MemPrimitives.scala 110:228:@48331.4]
  wire  _T_4941; // @[MemPrimitives.scala 110:228:@48335.4]
  wire  _T_4947; // @[MemPrimitives.scala 110:228:@48339.4]
  wire  _T_4949; // @[MemPrimitives.scala 123:41:@48359.4]
  wire  _T_4950; // @[MemPrimitives.scala 123:41:@48360.4]
  wire  _T_4951; // @[MemPrimitives.scala 123:41:@48361.4]
  wire  _T_4952; // @[MemPrimitives.scala 123:41:@48362.4]
  wire  _T_4953; // @[MemPrimitives.scala 123:41:@48363.4]
  wire  _T_4954; // @[MemPrimitives.scala 123:41:@48364.4]
  wire  _T_4955; // @[MemPrimitives.scala 123:41:@48365.4]
  wire  _T_4956; // @[MemPrimitives.scala 123:41:@48366.4]
  wire  _T_4957; // @[MemPrimitives.scala 123:41:@48367.4]
  wire  _T_4958; // @[MemPrimitives.scala 123:41:@48368.4]
  wire  _T_4959; // @[MemPrimitives.scala 123:41:@48369.4]
  wire  _T_4960; // @[MemPrimitives.scala 123:41:@48370.4]
  wire  _T_4961; // @[MemPrimitives.scala 123:41:@48371.4]
  wire  _T_4962; // @[MemPrimitives.scala 123:41:@48372.4]
  wire  _T_4963; // @[MemPrimitives.scala 123:41:@48373.4]
  wire [9:0] _T_4965; // @[Cat.scala 30:58:@48375.4]
  wire [9:0] _T_4967; // @[Cat.scala 30:58:@48377.4]
  wire [9:0] _T_4969; // @[Cat.scala 30:58:@48379.4]
  wire [9:0] _T_4971; // @[Cat.scala 30:58:@48381.4]
  wire [9:0] _T_4973; // @[Cat.scala 30:58:@48383.4]
  wire [9:0] _T_4975; // @[Cat.scala 30:58:@48385.4]
  wire [9:0] _T_4977; // @[Cat.scala 30:58:@48387.4]
  wire [9:0] _T_4979; // @[Cat.scala 30:58:@48389.4]
  wire [9:0] _T_4981; // @[Cat.scala 30:58:@48391.4]
  wire [9:0] _T_4983; // @[Cat.scala 30:58:@48393.4]
  wire [9:0] _T_4985; // @[Cat.scala 30:58:@48395.4]
  wire [9:0] _T_4987; // @[Cat.scala 30:58:@48397.4]
  wire [9:0] _T_4989; // @[Cat.scala 30:58:@48399.4]
  wire [9:0] _T_4991; // @[Cat.scala 30:58:@48401.4]
  wire [9:0] _T_4993; // @[Cat.scala 30:58:@48403.4]
  wire [9:0] _T_4994; // @[Mux.scala 31:69:@48404.4]
  wire [9:0] _T_4995; // @[Mux.scala 31:69:@48405.4]
  wire [9:0] _T_4996; // @[Mux.scala 31:69:@48406.4]
  wire [9:0] _T_4997; // @[Mux.scala 31:69:@48407.4]
  wire [9:0] _T_4998; // @[Mux.scala 31:69:@48408.4]
  wire [9:0] _T_4999; // @[Mux.scala 31:69:@48409.4]
  wire [9:0] _T_5000; // @[Mux.scala 31:69:@48410.4]
  wire [9:0] _T_5001; // @[Mux.scala 31:69:@48411.4]
  wire [9:0] _T_5002; // @[Mux.scala 31:69:@48412.4]
  wire [9:0] _T_5003; // @[Mux.scala 31:69:@48413.4]
  wire [9:0] _T_5004; // @[Mux.scala 31:69:@48414.4]
  wire [9:0] _T_5005; // @[Mux.scala 31:69:@48415.4]
  wire [9:0] _T_5006; // @[Mux.scala 31:69:@48416.4]
  wire [9:0] _T_5007; // @[Mux.scala 31:69:@48417.4]
  wire  _T_5015; // @[MemPrimitives.scala 110:228:@48426.4]
  wire  _T_5021; // @[MemPrimitives.scala 110:228:@48430.4]
  wire  _T_5027; // @[MemPrimitives.scala 110:228:@48434.4]
  wire  _T_5033; // @[MemPrimitives.scala 110:228:@48438.4]
  wire  _T_5039; // @[MemPrimitives.scala 110:228:@48442.4]
  wire  _T_5045; // @[MemPrimitives.scala 110:228:@48446.4]
  wire  _T_5051; // @[MemPrimitives.scala 110:228:@48450.4]
  wire  _T_5057; // @[MemPrimitives.scala 110:228:@48454.4]
  wire  _T_5063; // @[MemPrimitives.scala 110:228:@48458.4]
  wire  _T_5069; // @[MemPrimitives.scala 110:228:@48462.4]
  wire  _T_5075; // @[MemPrimitives.scala 110:228:@48466.4]
  wire  _T_5081; // @[MemPrimitives.scala 110:228:@48470.4]
  wire  _T_5087; // @[MemPrimitives.scala 110:228:@48474.4]
  wire  _T_5093; // @[MemPrimitives.scala 110:228:@48478.4]
  wire  _T_5099; // @[MemPrimitives.scala 110:228:@48482.4]
  wire  _T_5101; // @[MemPrimitives.scala 123:41:@48502.4]
  wire  _T_5102; // @[MemPrimitives.scala 123:41:@48503.4]
  wire  _T_5103; // @[MemPrimitives.scala 123:41:@48504.4]
  wire  _T_5104; // @[MemPrimitives.scala 123:41:@48505.4]
  wire  _T_5105; // @[MemPrimitives.scala 123:41:@48506.4]
  wire  _T_5106; // @[MemPrimitives.scala 123:41:@48507.4]
  wire  _T_5107; // @[MemPrimitives.scala 123:41:@48508.4]
  wire  _T_5108; // @[MemPrimitives.scala 123:41:@48509.4]
  wire  _T_5109; // @[MemPrimitives.scala 123:41:@48510.4]
  wire  _T_5110; // @[MemPrimitives.scala 123:41:@48511.4]
  wire  _T_5111; // @[MemPrimitives.scala 123:41:@48512.4]
  wire  _T_5112; // @[MemPrimitives.scala 123:41:@48513.4]
  wire  _T_5113; // @[MemPrimitives.scala 123:41:@48514.4]
  wire  _T_5114; // @[MemPrimitives.scala 123:41:@48515.4]
  wire  _T_5115; // @[MemPrimitives.scala 123:41:@48516.4]
  wire [9:0] _T_5117; // @[Cat.scala 30:58:@48518.4]
  wire [9:0] _T_5119; // @[Cat.scala 30:58:@48520.4]
  wire [9:0] _T_5121; // @[Cat.scala 30:58:@48522.4]
  wire [9:0] _T_5123; // @[Cat.scala 30:58:@48524.4]
  wire [9:0] _T_5125; // @[Cat.scala 30:58:@48526.4]
  wire [9:0] _T_5127; // @[Cat.scala 30:58:@48528.4]
  wire [9:0] _T_5129; // @[Cat.scala 30:58:@48530.4]
  wire [9:0] _T_5131; // @[Cat.scala 30:58:@48532.4]
  wire [9:0] _T_5133; // @[Cat.scala 30:58:@48534.4]
  wire [9:0] _T_5135; // @[Cat.scala 30:58:@48536.4]
  wire [9:0] _T_5137; // @[Cat.scala 30:58:@48538.4]
  wire [9:0] _T_5139; // @[Cat.scala 30:58:@48540.4]
  wire [9:0] _T_5141; // @[Cat.scala 30:58:@48542.4]
  wire [9:0] _T_5143; // @[Cat.scala 30:58:@48544.4]
  wire [9:0] _T_5145; // @[Cat.scala 30:58:@48546.4]
  wire [9:0] _T_5146; // @[Mux.scala 31:69:@48547.4]
  wire [9:0] _T_5147; // @[Mux.scala 31:69:@48548.4]
  wire [9:0] _T_5148; // @[Mux.scala 31:69:@48549.4]
  wire [9:0] _T_5149; // @[Mux.scala 31:69:@48550.4]
  wire [9:0] _T_5150; // @[Mux.scala 31:69:@48551.4]
  wire [9:0] _T_5151; // @[Mux.scala 31:69:@48552.4]
  wire [9:0] _T_5152; // @[Mux.scala 31:69:@48553.4]
  wire [9:0] _T_5153; // @[Mux.scala 31:69:@48554.4]
  wire [9:0] _T_5154; // @[Mux.scala 31:69:@48555.4]
  wire [9:0] _T_5155; // @[Mux.scala 31:69:@48556.4]
  wire [9:0] _T_5156; // @[Mux.scala 31:69:@48557.4]
  wire [9:0] _T_5157; // @[Mux.scala 31:69:@48558.4]
  wire [9:0] _T_5158; // @[Mux.scala 31:69:@48559.4]
  wire [9:0] _T_5159; // @[Mux.scala 31:69:@48560.4]
  wire  _T_5167; // @[MemPrimitives.scala 110:228:@48569.4]
  wire  _T_5173; // @[MemPrimitives.scala 110:228:@48573.4]
  wire  _T_5179; // @[MemPrimitives.scala 110:228:@48577.4]
  wire  _T_5185; // @[MemPrimitives.scala 110:228:@48581.4]
  wire  _T_5191; // @[MemPrimitives.scala 110:228:@48585.4]
  wire  _T_5197; // @[MemPrimitives.scala 110:228:@48589.4]
  wire  _T_5203; // @[MemPrimitives.scala 110:228:@48593.4]
  wire  _T_5209; // @[MemPrimitives.scala 110:228:@48597.4]
  wire  _T_5215; // @[MemPrimitives.scala 110:228:@48601.4]
  wire  _T_5221; // @[MemPrimitives.scala 110:228:@48605.4]
  wire  _T_5227; // @[MemPrimitives.scala 110:228:@48609.4]
  wire  _T_5233; // @[MemPrimitives.scala 110:228:@48613.4]
  wire  _T_5239; // @[MemPrimitives.scala 110:228:@48617.4]
  wire  _T_5245; // @[MemPrimitives.scala 110:228:@48621.4]
  wire  _T_5251; // @[MemPrimitives.scala 110:228:@48625.4]
  wire  _T_5253; // @[MemPrimitives.scala 123:41:@48645.4]
  wire  _T_5254; // @[MemPrimitives.scala 123:41:@48646.4]
  wire  _T_5255; // @[MemPrimitives.scala 123:41:@48647.4]
  wire  _T_5256; // @[MemPrimitives.scala 123:41:@48648.4]
  wire  _T_5257; // @[MemPrimitives.scala 123:41:@48649.4]
  wire  _T_5258; // @[MemPrimitives.scala 123:41:@48650.4]
  wire  _T_5259; // @[MemPrimitives.scala 123:41:@48651.4]
  wire  _T_5260; // @[MemPrimitives.scala 123:41:@48652.4]
  wire  _T_5261; // @[MemPrimitives.scala 123:41:@48653.4]
  wire  _T_5262; // @[MemPrimitives.scala 123:41:@48654.4]
  wire  _T_5263; // @[MemPrimitives.scala 123:41:@48655.4]
  wire  _T_5264; // @[MemPrimitives.scala 123:41:@48656.4]
  wire  _T_5265; // @[MemPrimitives.scala 123:41:@48657.4]
  wire  _T_5266; // @[MemPrimitives.scala 123:41:@48658.4]
  wire  _T_5267; // @[MemPrimitives.scala 123:41:@48659.4]
  wire [9:0] _T_5269; // @[Cat.scala 30:58:@48661.4]
  wire [9:0] _T_5271; // @[Cat.scala 30:58:@48663.4]
  wire [9:0] _T_5273; // @[Cat.scala 30:58:@48665.4]
  wire [9:0] _T_5275; // @[Cat.scala 30:58:@48667.4]
  wire [9:0] _T_5277; // @[Cat.scala 30:58:@48669.4]
  wire [9:0] _T_5279; // @[Cat.scala 30:58:@48671.4]
  wire [9:0] _T_5281; // @[Cat.scala 30:58:@48673.4]
  wire [9:0] _T_5283; // @[Cat.scala 30:58:@48675.4]
  wire [9:0] _T_5285; // @[Cat.scala 30:58:@48677.4]
  wire [9:0] _T_5287; // @[Cat.scala 30:58:@48679.4]
  wire [9:0] _T_5289; // @[Cat.scala 30:58:@48681.4]
  wire [9:0] _T_5291; // @[Cat.scala 30:58:@48683.4]
  wire [9:0] _T_5293; // @[Cat.scala 30:58:@48685.4]
  wire [9:0] _T_5295; // @[Cat.scala 30:58:@48687.4]
  wire [9:0] _T_5297; // @[Cat.scala 30:58:@48689.4]
  wire [9:0] _T_5298; // @[Mux.scala 31:69:@48690.4]
  wire [9:0] _T_5299; // @[Mux.scala 31:69:@48691.4]
  wire [9:0] _T_5300; // @[Mux.scala 31:69:@48692.4]
  wire [9:0] _T_5301; // @[Mux.scala 31:69:@48693.4]
  wire [9:0] _T_5302; // @[Mux.scala 31:69:@48694.4]
  wire [9:0] _T_5303; // @[Mux.scala 31:69:@48695.4]
  wire [9:0] _T_5304; // @[Mux.scala 31:69:@48696.4]
  wire [9:0] _T_5305; // @[Mux.scala 31:69:@48697.4]
  wire [9:0] _T_5306; // @[Mux.scala 31:69:@48698.4]
  wire [9:0] _T_5307; // @[Mux.scala 31:69:@48699.4]
  wire [9:0] _T_5308; // @[Mux.scala 31:69:@48700.4]
  wire [9:0] _T_5309; // @[Mux.scala 31:69:@48701.4]
  wire [9:0] _T_5310; // @[Mux.scala 31:69:@48702.4]
  wire [9:0] _T_5311; // @[Mux.scala 31:69:@48703.4]
  wire  _T_5319; // @[MemPrimitives.scala 110:228:@48712.4]
  wire  _T_5325; // @[MemPrimitives.scala 110:228:@48716.4]
  wire  _T_5331; // @[MemPrimitives.scala 110:228:@48720.4]
  wire  _T_5337; // @[MemPrimitives.scala 110:228:@48724.4]
  wire  _T_5343; // @[MemPrimitives.scala 110:228:@48728.4]
  wire  _T_5349; // @[MemPrimitives.scala 110:228:@48732.4]
  wire  _T_5355; // @[MemPrimitives.scala 110:228:@48736.4]
  wire  _T_5361; // @[MemPrimitives.scala 110:228:@48740.4]
  wire  _T_5367; // @[MemPrimitives.scala 110:228:@48744.4]
  wire  _T_5373; // @[MemPrimitives.scala 110:228:@48748.4]
  wire  _T_5379; // @[MemPrimitives.scala 110:228:@48752.4]
  wire  _T_5385; // @[MemPrimitives.scala 110:228:@48756.4]
  wire  _T_5391; // @[MemPrimitives.scala 110:228:@48760.4]
  wire  _T_5397; // @[MemPrimitives.scala 110:228:@48764.4]
  wire  _T_5403; // @[MemPrimitives.scala 110:228:@48768.4]
  wire  _T_5405; // @[MemPrimitives.scala 123:41:@48788.4]
  wire  _T_5406; // @[MemPrimitives.scala 123:41:@48789.4]
  wire  _T_5407; // @[MemPrimitives.scala 123:41:@48790.4]
  wire  _T_5408; // @[MemPrimitives.scala 123:41:@48791.4]
  wire  _T_5409; // @[MemPrimitives.scala 123:41:@48792.4]
  wire  _T_5410; // @[MemPrimitives.scala 123:41:@48793.4]
  wire  _T_5411; // @[MemPrimitives.scala 123:41:@48794.4]
  wire  _T_5412; // @[MemPrimitives.scala 123:41:@48795.4]
  wire  _T_5413; // @[MemPrimitives.scala 123:41:@48796.4]
  wire  _T_5414; // @[MemPrimitives.scala 123:41:@48797.4]
  wire  _T_5415; // @[MemPrimitives.scala 123:41:@48798.4]
  wire  _T_5416; // @[MemPrimitives.scala 123:41:@48799.4]
  wire  _T_5417; // @[MemPrimitives.scala 123:41:@48800.4]
  wire  _T_5418; // @[MemPrimitives.scala 123:41:@48801.4]
  wire  _T_5419; // @[MemPrimitives.scala 123:41:@48802.4]
  wire [9:0] _T_5421; // @[Cat.scala 30:58:@48804.4]
  wire [9:0] _T_5423; // @[Cat.scala 30:58:@48806.4]
  wire [9:0] _T_5425; // @[Cat.scala 30:58:@48808.4]
  wire [9:0] _T_5427; // @[Cat.scala 30:58:@48810.4]
  wire [9:0] _T_5429; // @[Cat.scala 30:58:@48812.4]
  wire [9:0] _T_5431; // @[Cat.scala 30:58:@48814.4]
  wire [9:0] _T_5433; // @[Cat.scala 30:58:@48816.4]
  wire [9:0] _T_5435; // @[Cat.scala 30:58:@48818.4]
  wire [9:0] _T_5437; // @[Cat.scala 30:58:@48820.4]
  wire [9:0] _T_5439; // @[Cat.scala 30:58:@48822.4]
  wire [9:0] _T_5441; // @[Cat.scala 30:58:@48824.4]
  wire [9:0] _T_5443; // @[Cat.scala 30:58:@48826.4]
  wire [9:0] _T_5445; // @[Cat.scala 30:58:@48828.4]
  wire [9:0] _T_5447; // @[Cat.scala 30:58:@48830.4]
  wire [9:0] _T_5449; // @[Cat.scala 30:58:@48832.4]
  wire [9:0] _T_5450; // @[Mux.scala 31:69:@48833.4]
  wire [9:0] _T_5451; // @[Mux.scala 31:69:@48834.4]
  wire [9:0] _T_5452; // @[Mux.scala 31:69:@48835.4]
  wire [9:0] _T_5453; // @[Mux.scala 31:69:@48836.4]
  wire [9:0] _T_5454; // @[Mux.scala 31:69:@48837.4]
  wire [9:0] _T_5455; // @[Mux.scala 31:69:@48838.4]
  wire [9:0] _T_5456; // @[Mux.scala 31:69:@48839.4]
  wire [9:0] _T_5457; // @[Mux.scala 31:69:@48840.4]
  wire [9:0] _T_5458; // @[Mux.scala 31:69:@48841.4]
  wire [9:0] _T_5459; // @[Mux.scala 31:69:@48842.4]
  wire [9:0] _T_5460; // @[Mux.scala 31:69:@48843.4]
  wire [9:0] _T_5461; // @[Mux.scala 31:69:@48844.4]
  wire [9:0] _T_5462; // @[Mux.scala 31:69:@48845.4]
  wire [9:0] _T_5463; // @[Mux.scala 31:69:@48846.4]
  wire  _T_5471; // @[MemPrimitives.scala 110:228:@48855.4]
  wire  _T_5477; // @[MemPrimitives.scala 110:228:@48859.4]
  wire  _T_5483; // @[MemPrimitives.scala 110:228:@48863.4]
  wire  _T_5489; // @[MemPrimitives.scala 110:228:@48867.4]
  wire  _T_5495; // @[MemPrimitives.scala 110:228:@48871.4]
  wire  _T_5501; // @[MemPrimitives.scala 110:228:@48875.4]
  wire  _T_5507; // @[MemPrimitives.scala 110:228:@48879.4]
  wire  _T_5513; // @[MemPrimitives.scala 110:228:@48883.4]
  wire  _T_5519; // @[MemPrimitives.scala 110:228:@48887.4]
  wire  _T_5525; // @[MemPrimitives.scala 110:228:@48891.4]
  wire  _T_5531; // @[MemPrimitives.scala 110:228:@48895.4]
  wire  _T_5537; // @[MemPrimitives.scala 110:228:@48899.4]
  wire  _T_5543; // @[MemPrimitives.scala 110:228:@48903.4]
  wire  _T_5549; // @[MemPrimitives.scala 110:228:@48907.4]
  wire  _T_5555; // @[MemPrimitives.scala 110:228:@48911.4]
  wire  _T_5557; // @[MemPrimitives.scala 123:41:@48931.4]
  wire  _T_5558; // @[MemPrimitives.scala 123:41:@48932.4]
  wire  _T_5559; // @[MemPrimitives.scala 123:41:@48933.4]
  wire  _T_5560; // @[MemPrimitives.scala 123:41:@48934.4]
  wire  _T_5561; // @[MemPrimitives.scala 123:41:@48935.4]
  wire  _T_5562; // @[MemPrimitives.scala 123:41:@48936.4]
  wire  _T_5563; // @[MemPrimitives.scala 123:41:@48937.4]
  wire  _T_5564; // @[MemPrimitives.scala 123:41:@48938.4]
  wire  _T_5565; // @[MemPrimitives.scala 123:41:@48939.4]
  wire  _T_5566; // @[MemPrimitives.scala 123:41:@48940.4]
  wire  _T_5567; // @[MemPrimitives.scala 123:41:@48941.4]
  wire  _T_5568; // @[MemPrimitives.scala 123:41:@48942.4]
  wire  _T_5569; // @[MemPrimitives.scala 123:41:@48943.4]
  wire  _T_5570; // @[MemPrimitives.scala 123:41:@48944.4]
  wire  _T_5571; // @[MemPrimitives.scala 123:41:@48945.4]
  wire [9:0] _T_5573; // @[Cat.scala 30:58:@48947.4]
  wire [9:0] _T_5575; // @[Cat.scala 30:58:@48949.4]
  wire [9:0] _T_5577; // @[Cat.scala 30:58:@48951.4]
  wire [9:0] _T_5579; // @[Cat.scala 30:58:@48953.4]
  wire [9:0] _T_5581; // @[Cat.scala 30:58:@48955.4]
  wire [9:0] _T_5583; // @[Cat.scala 30:58:@48957.4]
  wire [9:0] _T_5585; // @[Cat.scala 30:58:@48959.4]
  wire [9:0] _T_5587; // @[Cat.scala 30:58:@48961.4]
  wire [9:0] _T_5589; // @[Cat.scala 30:58:@48963.4]
  wire [9:0] _T_5591; // @[Cat.scala 30:58:@48965.4]
  wire [9:0] _T_5593; // @[Cat.scala 30:58:@48967.4]
  wire [9:0] _T_5595; // @[Cat.scala 30:58:@48969.4]
  wire [9:0] _T_5597; // @[Cat.scala 30:58:@48971.4]
  wire [9:0] _T_5599; // @[Cat.scala 30:58:@48973.4]
  wire [9:0] _T_5601; // @[Cat.scala 30:58:@48975.4]
  wire [9:0] _T_5602; // @[Mux.scala 31:69:@48976.4]
  wire [9:0] _T_5603; // @[Mux.scala 31:69:@48977.4]
  wire [9:0] _T_5604; // @[Mux.scala 31:69:@48978.4]
  wire [9:0] _T_5605; // @[Mux.scala 31:69:@48979.4]
  wire [9:0] _T_5606; // @[Mux.scala 31:69:@48980.4]
  wire [9:0] _T_5607; // @[Mux.scala 31:69:@48981.4]
  wire [9:0] _T_5608; // @[Mux.scala 31:69:@48982.4]
  wire [9:0] _T_5609; // @[Mux.scala 31:69:@48983.4]
  wire [9:0] _T_5610; // @[Mux.scala 31:69:@48984.4]
  wire [9:0] _T_5611; // @[Mux.scala 31:69:@48985.4]
  wire [9:0] _T_5612; // @[Mux.scala 31:69:@48986.4]
  wire [9:0] _T_5613; // @[Mux.scala 31:69:@48987.4]
  wire [9:0] _T_5614; // @[Mux.scala 31:69:@48988.4]
  wire [9:0] _T_5615; // @[Mux.scala 31:69:@48989.4]
  wire  _T_5623; // @[MemPrimitives.scala 110:228:@48998.4]
  wire  _T_5629; // @[MemPrimitives.scala 110:228:@49002.4]
  wire  _T_5635; // @[MemPrimitives.scala 110:228:@49006.4]
  wire  _T_5641; // @[MemPrimitives.scala 110:228:@49010.4]
  wire  _T_5647; // @[MemPrimitives.scala 110:228:@49014.4]
  wire  _T_5653; // @[MemPrimitives.scala 110:228:@49018.4]
  wire  _T_5659; // @[MemPrimitives.scala 110:228:@49022.4]
  wire  _T_5665; // @[MemPrimitives.scala 110:228:@49026.4]
  wire  _T_5671; // @[MemPrimitives.scala 110:228:@49030.4]
  wire  _T_5677; // @[MemPrimitives.scala 110:228:@49034.4]
  wire  _T_5683; // @[MemPrimitives.scala 110:228:@49038.4]
  wire  _T_5689; // @[MemPrimitives.scala 110:228:@49042.4]
  wire  _T_5695; // @[MemPrimitives.scala 110:228:@49046.4]
  wire  _T_5701; // @[MemPrimitives.scala 110:228:@49050.4]
  wire  _T_5707; // @[MemPrimitives.scala 110:228:@49054.4]
  wire  _T_5709; // @[MemPrimitives.scala 123:41:@49074.4]
  wire  _T_5710; // @[MemPrimitives.scala 123:41:@49075.4]
  wire  _T_5711; // @[MemPrimitives.scala 123:41:@49076.4]
  wire  _T_5712; // @[MemPrimitives.scala 123:41:@49077.4]
  wire  _T_5713; // @[MemPrimitives.scala 123:41:@49078.4]
  wire  _T_5714; // @[MemPrimitives.scala 123:41:@49079.4]
  wire  _T_5715; // @[MemPrimitives.scala 123:41:@49080.4]
  wire  _T_5716; // @[MemPrimitives.scala 123:41:@49081.4]
  wire  _T_5717; // @[MemPrimitives.scala 123:41:@49082.4]
  wire  _T_5718; // @[MemPrimitives.scala 123:41:@49083.4]
  wire  _T_5719; // @[MemPrimitives.scala 123:41:@49084.4]
  wire  _T_5720; // @[MemPrimitives.scala 123:41:@49085.4]
  wire  _T_5721; // @[MemPrimitives.scala 123:41:@49086.4]
  wire  _T_5722; // @[MemPrimitives.scala 123:41:@49087.4]
  wire  _T_5723; // @[MemPrimitives.scala 123:41:@49088.4]
  wire [9:0] _T_5725; // @[Cat.scala 30:58:@49090.4]
  wire [9:0] _T_5727; // @[Cat.scala 30:58:@49092.4]
  wire [9:0] _T_5729; // @[Cat.scala 30:58:@49094.4]
  wire [9:0] _T_5731; // @[Cat.scala 30:58:@49096.4]
  wire [9:0] _T_5733; // @[Cat.scala 30:58:@49098.4]
  wire [9:0] _T_5735; // @[Cat.scala 30:58:@49100.4]
  wire [9:0] _T_5737; // @[Cat.scala 30:58:@49102.4]
  wire [9:0] _T_5739; // @[Cat.scala 30:58:@49104.4]
  wire [9:0] _T_5741; // @[Cat.scala 30:58:@49106.4]
  wire [9:0] _T_5743; // @[Cat.scala 30:58:@49108.4]
  wire [9:0] _T_5745; // @[Cat.scala 30:58:@49110.4]
  wire [9:0] _T_5747; // @[Cat.scala 30:58:@49112.4]
  wire [9:0] _T_5749; // @[Cat.scala 30:58:@49114.4]
  wire [9:0] _T_5751; // @[Cat.scala 30:58:@49116.4]
  wire [9:0] _T_5753; // @[Cat.scala 30:58:@49118.4]
  wire [9:0] _T_5754; // @[Mux.scala 31:69:@49119.4]
  wire [9:0] _T_5755; // @[Mux.scala 31:69:@49120.4]
  wire [9:0] _T_5756; // @[Mux.scala 31:69:@49121.4]
  wire [9:0] _T_5757; // @[Mux.scala 31:69:@49122.4]
  wire [9:0] _T_5758; // @[Mux.scala 31:69:@49123.4]
  wire [9:0] _T_5759; // @[Mux.scala 31:69:@49124.4]
  wire [9:0] _T_5760; // @[Mux.scala 31:69:@49125.4]
  wire [9:0] _T_5761; // @[Mux.scala 31:69:@49126.4]
  wire [9:0] _T_5762; // @[Mux.scala 31:69:@49127.4]
  wire [9:0] _T_5763; // @[Mux.scala 31:69:@49128.4]
  wire [9:0] _T_5764; // @[Mux.scala 31:69:@49129.4]
  wire [9:0] _T_5765; // @[Mux.scala 31:69:@49130.4]
  wire [9:0] _T_5766; // @[Mux.scala 31:69:@49131.4]
  wire [9:0] _T_5767; // @[Mux.scala 31:69:@49132.4]
  wire  _T_5772; // @[MemPrimitives.scala 110:210:@49139.4]
  wire  _T_5775; // @[MemPrimitives.scala 110:228:@49141.4]
  wire  _T_5778; // @[MemPrimitives.scala 110:210:@49143.4]
  wire  _T_5781; // @[MemPrimitives.scala 110:228:@49145.4]
  wire  _T_5784; // @[MemPrimitives.scala 110:210:@49147.4]
  wire  _T_5787; // @[MemPrimitives.scala 110:228:@49149.4]
  wire  _T_5790; // @[MemPrimitives.scala 110:210:@49151.4]
  wire  _T_5793; // @[MemPrimitives.scala 110:228:@49153.4]
  wire  _T_5796; // @[MemPrimitives.scala 110:210:@49155.4]
  wire  _T_5799; // @[MemPrimitives.scala 110:228:@49157.4]
  wire  _T_5802; // @[MemPrimitives.scala 110:210:@49159.4]
  wire  _T_5805; // @[MemPrimitives.scala 110:228:@49161.4]
  wire  _T_5808; // @[MemPrimitives.scala 110:210:@49163.4]
  wire  _T_5811; // @[MemPrimitives.scala 110:228:@49165.4]
  wire  _T_5814; // @[MemPrimitives.scala 110:210:@49167.4]
  wire  _T_5817; // @[MemPrimitives.scala 110:228:@49169.4]
  wire  _T_5820; // @[MemPrimitives.scala 110:210:@49171.4]
  wire  _T_5823; // @[MemPrimitives.scala 110:228:@49173.4]
  wire  _T_5826; // @[MemPrimitives.scala 110:210:@49175.4]
  wire  _T_5829; // @[MemPrimitives.scala 110:228:@49177.4]
  wire  _T_5832; // @[MemPrimitives.scala 110:210:@49179.4]
  wire  _T_5835; // @[MemPrimitives.scala 110:228:@49181.4]
  wire  _T_5838; // @[MemPrimitives.scala 110:210:@49183.4]
  wire  _T_5841; // @[MemPrimitives.scala 110:228:@49185.4]
  wire  _T_5844; // @[MemPrimitives.scala 110:210:@49187.4]
  wire  _T_5847; // @[MemPrimitives.scala 110:228:@49189.4]
  wire  _T_5850; // @[MemPrimitives.scala 110:210:@49191.4]
  wire  _T_5853; // @[MemPrimitives.scala 110:228:@49193.4]
  wire  _T_5856; // @[MemPrimitives.scala 110:210:@49195.4]
  wire  _T_5859; // @[MemPrimitives.scala 110:228:@49197.4]
  wire  _T_5861; // @[MemPrimitives.scala 123:41:@49217.4]
  wire  _T_5862; // @[MemPrimitives.scala 123:41:@49218.4]
  wire  _T_5863; // @[MemPrimitives.scala 123:41:@49219.4]
  wire  _T_5864; // @[MemPrimitives.scala 123:41:@49220.4]
  wire  _T_5865; // @[MemPrimitives.scala 123:41:@49221.4]
  wire  _T_5866; // @[MemPrimitives.scala 123:41:@49222.4]
  wire  _T_5867; // @[MemPrimitives.scala 123:41:@49223.4]
  wire  _T_5868; // @[MemPrimitives.scala 123:41:@49224.4]
  wire  _T_5869; // @[MemPrimitives.scala 123:41:@49225.4]
  wire  _T_5870; // @[MemPrimitives.scala 123:41:@49226.4]
  wire  _T_5871; // @[MemPrimitives.scala 123:41:@49227.4]
  wire  _T_5872; // @[MemPrimitives.scala 123:41:@49228.4]
  wire  _T_5873; // @[MemPrimitives.scala 123:41:@49229.4]
  wire  _T_5874; // @[MemPrimitives.scala 123:41:@49230.4]
  wire  _T_5875; // @[MemPrimitives.scala 123:41:@49231.4]
  wire [9:0] _T_5877; // @[Cat.scala 30:58:@49233.4]
  wire [9:0] _T_5879; // @[Cat.scala 30:58:@49235.4]
  wire [9:0] _T_5881; // @[Cat.scala 30:58:@49237.4]
  wire [9:0] _T_5883; // @[Cat.scala 30:58:@49239.4]
  wire [9:0] _T_5885; // @[Cat.scala 30:58:@49241.4]
  wire [9:0] _T_5887; // @[Cat.scala 30:58:@49243.4]
  wire [9:0] _T_5889; // @[Cat.scala 30:58:@49245.4]
  wire [9:0] _T_5891; // @[Cat.scala 30:58:@49247.4]
  wire [9:0] _T_5893; // @[Cat.scala 30:58:@49249.4]
  wire [9:0] _T_5895; // @[Cat.scala 30:58:@49251.4]
  wire [9:0] _T_5897; // @[Cat.scala 30:58:@49253.4]
  wire [9:0] _T_5899; // @[Cat.scala 30:58:@49255.4]
  wire [9:0] _T_5901; // @[Cat.scala 30:58:@49257.4]
  wire [9:0] _T_5903; // @[Cat.scala 30:58:@49259.4]
  wire [9:0] _T_5905; // @[Cat.scala 30:58:@49261.4]
  wire [9:0] _T_5906; // @[Mux.scala 31:69:@49262.4]
  wire [9:0] _T_5907; // @[Mux.scala 31:69:@49263.4]
  wire [9:0] _T_5908; // @[Mux.scala 31:69:@49264.4]
  wire [9:0] _T_5909; // @[Mux.scala 31:69:@49265.4]
  wire [9:0] _T_5910; // @[Mux.scala 31:69:@49266.4]
  wire [9:0] _T_5911; // @[Mux.scala 31:69:@49267.4]
  wire [9:0] _T_5912; // @[Mux.scala 31:69:@49268.4]
  wire [9:0] _T_5913; // @[Mux.scala 31:69:@49269.4]
  wire [9:0] _T_5914; // @[Mux.scala 31:69:@49270.4]
  wire [9:0] _T_5915; // @[Mux.scala 31:69:@49271.4]
  wire [9:0] _T_5916; // @[Mux.scala 31:69:@49272.4]
  wire [9:0] _T_5917; // @[Mux.scala 31:69:@49273.4]
  wire [9:0] _T_5918; // @[Mux.scala 31:69:@49274.4]
  wire [9:0] _T_5919; // @[Mux.scala 31:69:@49275.4]
  wire  _T_5924; // @[MemPrimitives.scala 110:210:@49282.4]
  wire  _T_5927; // @[MemPrimitives.scala 110:228:@49284.4]
  wire  _T_5930; // @[MemPrimitives.scala 110:210:@49286.4]
  wire  _T_5933; // @[MemPrimitives.scala 110:228:@49288.4]
  wire  _T_5936; // @[MemPrimitives.scala 110:210:@49290.4]
  wire  _T_5939; // @[MemPrimitives.scala 110:228:@49292.4]
  wire  _T_5942; // @[MemPrimitives.scala 110:210:@49294.4]
  wire  _T_5945; // @[MemPrimitives.scala 110:228:@49296.4]
  wire  _T_5948; // @[MemPrimitives.scala 110:210:@49298.4]
  wire  _T_5951; // @[MemPrimitives.scala 110:228:@49300.4]
  wire  _T_5954; // @[MemPrimitives.scala 110:210:@49302.4]
  wire  _T_5957; // @[MemPrimitives.scala 110:228:@49304.4]
  wire  _T_5960; // @[MemPrimitives.scala 110:210:@49306.4]
  wire  _T_5963; // @[MemPrimitives.scala 110:228:@49308.4]
  wire  _T_5966; // @[MemPrimitives.scala 110:210:@49310.4]
  wire  _T_5969; // @[MemPrimitives.scala 110:228:@49312.4]
  wire  _T_5972; // @[MemPrimitives.scala 110:210:@49314.4]
  wire  _T_5975; // @[MemPrimitives.scala 110:228:@49316.4]
  wire  _T_5978; // @[MemPrimitives.scala 110:210:@49318.4]
  wire  _T_5981; // @[MemPrimitives.scala 110:228:@49320.4]
  wire  _T_5984; // @[MemPrimitives.scala 110:210:@49322.4]
  wire  _T_5987; // @[MemPrimitives.scala 110:228:@49324.4]
  wire  _T_5990; // @[MemPrimitives.scala 110:210:@49326.4]
  wire  _T_5993; // @[MemPrimitives.scala 110:228:@49328.4]
  wire  _T_5996; // @[MemPrimitives.scala 110:210:@49330.4]
  wire  _T_5999; // @[MemPrimitives.scala 110:228:@49332.4]
  wire  _T_6002; // @[MemPrimitives.scala 110:210:@49334.4]
  wire  _T_6005; // @[MemPrimitives.scala 110:228:@49336.4]
  wire  _T_6008; // @[MemPrimitives.scala 110:210:@49338.4]
  wire  _T_6011; // @[MemPrimitives.scala 110:228:@49340.4]
  wire  _T_6013; // @[MemPrimitives.scala 123:41:@49360.4]
  wire  _T_6014; // @[MemPrimitives.scala 123:41:@49361.4]
  wire  _T_6015; // @[MemPrimitives.scala 123:41:@49362.4]
  wire  _T_6016; // @[MemPrimitives.scala 123:41:@49363.4]
  wire  _T_6017; // @[MemPrimitives.scala 123:41:@49364.4]
  wire  _T_6018; // @[MemPrimitives.scala 123:41:@49365.4]
  wire  _T_6019; // @[MemPrimitives.scala 123:41:@49366.4]
  wire  _T_6020; // @[MemPrimitives.scala 123:41:@49367.4]
  wire  _T_6021; // @[MemPrimitives.scala 123:41:@49368.4]
  wire  _T_6022; // @[MemPrimitives.scala 123:41:@49369.4]
  wire  _T_6023; // @[MemPrimitives.scala 123:41:@49370.4]
  wire  _T_6024; // @[MemPrimitives.scala 123:41:@49371.4]
  wire  _T_6025; // @[MemPrimitives.scala 123:41:@49372.4]
  wire  _T_6026; // @[MemPrimitives.scala 123:41:@49373.4]
  wire  _T_6027; // @[MemPrimitives.scala 123:41:@49374.4]
  wire [9:0] _T_6029; // @[Cat.scala 30:58:@49376.4]
  wire [9:0] _T_6031; // @[Cat.scala 30:58:@49378.4]
  wire [9:0] _T_6033; // @[Cat.scala 30:58:@49380.4]
  wire [9:0] _T_6035; // @[Cat.scala 30:58:@49382.4]
  wire [9:0] _T_6037; // @[Cat.scala 30:58:@49384.4]
  wire [9:0] _T_6039; // @[Cat.scala 30:58:@49386.4]
  wire [9:0] _T_6041; // @[Cat.scala 30:58:@49388.4]
  wire [9:0] _T_6043; // @[Cat.scala 30:58:@49390.4]
  wire [9:0] _T_6045; // @[Cat.scala 30:58:@49392.4]
  wire [9:0] _T_6047; // @[Cat.scala 30:58:@49394.4]
  wire [9:0] _T_6049; // @[Cat.scala 30:58:@49396.4]
  wire [9:0] _T_6051; // @[Cat.scala 30:58:@49398.4]
  wire [9:0] _T_6053; // @[Cat.scala 30:58:@49400.4]
  wire [9:0] _T_6055; // @[Cat.scala 30:58:@49402.4]
  wire [9:0] _T_6057; // @[Cat.scala 30:58:@49404.4]
  wire [9:0] _T_6058; // @[Mux.scala 31:69:@49405.4]
  wire [9:0] _T_6059; // @[Mux.scala 31:69:@49406.4]
  wire [9:0] _T_6060; // @[Mux.scala 31:69:@49407.4]
  wire [9:0] _T_6061; // @[Mux.scala 31:69:@49408.4]
  wire [9:0] _T_6062; // @[Mux.scala 31:69:@49409.4]
  wire [9:0] _T_6063; // @[Mux.scala 31:69:@49410.4]
  wire [9:0] _T_6064; // @[Mux.scala 31:69:@49411.4]
  wire [9:0] _T_6065; // @[Mux.scala 31:69:@49412.4]
  wire [9:0] _T_6066; // @[Mux.scala 31:69:@49413.4]
  wire [9:0] _T_6067; // @[Mux.scala 31:69:@49414.4]
  wire [9:0] _T_6068; // @[Mux.scala 31:69:@49415.4]
  wire [9:0] _T_6069; // @[Mux.scala 31:69:@49416.4]
  wire [9:0] _T_6070; // @[Mux.scala 31:69:@49417.4]
  wire [9:0] _T_6071; // @[Mux.scala 31:69:@49418.4]
  wire  _T_6079; // @[MemPrimitives.scala 110:228:@49427.4]
  wire  _T_6085; // @[MemPrimitives.scala 110:228:@49431.4]
  wire  _T_6091; // @[MemPrimitives.scala 110:228:@49435.4]
  wire  _T_6097; // @[MemPrimitives.scala 110:228:@49439.4]
  wire  _T_6103; // @[MemPrimitives.scala 110:228:@49443.4]
  wire  _T_6109; // @[MemPrimitives.scala 110:228:@49447.4]
  wire  _T_6115; // @[MemPrimitives.scala 110:228:@49451.4]
  wire  _T_6121; // @[MemPrimitives.scala 110:228:@49455.4]
  wire  _T_6127; // @[MemPrimitives.scala 110:228:@49459.4]
  wire  _T_6133; // @[MemPrimitives.scala 110:228:@49463.4]
  wire  _T_6139; // @[MemPrimitives.scala 110:228:@49467.4]
  wire  _T_6145; // @[MemPrimitives.scala 110:228:@49471.4]
  wire  _T_6151; // @[MemPrimitives.scala 110:228:@49475.4]
  wire  _T_6157; // @[MemPrimitives.scala 110:228:@49479.4]
  wire  _T_6163; // @[MemPrimitives.scala 110:228:@49483.4]
  wire  _T_6165; // @[MemPrimitives.scala 123:41:@49503.4]
  wire  _T_6166; // @[MemPrimitives.scala 123:41:@49504.4]
  wire  _T_6167; // @[MemPrimitives.scala 123:41:@49505.4]
  wire  _T_6168; // @[MemPrimitives.scala 123:41:@49506.4]
  wire  _T_6169; // @[MemPrimitives.scala 123:41:@49507.4]
  wire  _T_6170; // @[MemPrimitives.scala 123:41:@49508.4]
  wire  _T_6171; // @[MemPrimitives.scala 123:41:@49509.4]
  wire  _T_6172; // @[MemPrimitives.scala 123:41:@49510.4]
  wire  _T_6173; // @[MemPrimitives.scala 123:41:@49511.4]
  wire  _T_6174; // @[MemPrimitives.scala 123:41:@49512.4]
  wire  _T_6175; // @[MemPrimitives.scala 123:41:@49513.4]
  wire  _T_6176; // @[MemPrimitives.scala 123:41:@49514.4]
  wire  _T_6177; // @[MemPrimitives.scala 123:41:@49515.4]
  wire  _T_6178; // @[MemPrimitives.scala 123:41:@49516.4]
  wire  _T_6179; // @[MemPrimitives.scala 123:41:@49517.4]
  wire [9:0] _T_6181; // @[Cat.scala 30:58:@49519.4]
  wire [9:0] _T_6183; // @[Cat.scala 30:58:@49521.4]
  wire [9:0] _T_6185; // @[Cat.scala 30:58:@49523.4]
  wire [9:0] _T_6187; // @[Cat.scala 30:58:@49525.4]
  wire [9:0] _T_6189; // @[Cat.scala 30:58:@49527.4]
  wire [9:0] _T_6191; // @[Cat.scala 30:58:@49529.4]
  wire [9:0] _T_6193; // @[Cat.scala 30:58:@49531.4]
  wire [9:0] _T_6195; // @[Cat.scala 30:58:@49533.4]
  wire [9:0] _T_6197; // @[Cat.scala 30:58:@49535.4]
  wire [9:0] _T_6199; // @[Cat.scala 30:58:@49537.4]
  wire [9:0] _T_6201; // @[Cat.scala 30:58:@49539.4]
  wire [9:0] _T_6203; // @[Cat.scala 30:58:@49541.4]
  wire [9:0] _T_6205; // @[Cat.scala 30:58:@49543.4]
  wire [9:0] _T_6207; // @[Cat.scala 30:58:@49545.4]
  wire [9:0] _T_6209; // @[Cat.scala 30:58:@49547.4]
  wire [9:0] _T_6210; // @[Mux.scala 31:69:@49548.4]
  wire [9:0] _T_6211; // @[Mux.scala 31:69:@49549.4]
  wire [9:0] _T_6212; // @[Mux.scala 31:69:@49550.4]
  wire [9:0] _T_6213; // @[Mux.scala 31:69:@49551.4]
  wire [9:0] _T_6214; // @[Mux.scala 31:69:@49552.4]
  wire [9:0] _T_6215; // @[Mux.scala 31:69:@49553.4]
  wire [9:0] _T_6216; // @[Mux.scala 31:69:@49554.4]
  wire [9:0] _T_6217; // @[Mux.scala 31:69:@49555.4]
  wire [9:0] _T_6218; // @[Mux.scala 31:69:@49556.4]
  wire [9:0] _T_6219; // @[Mux.scala 31:69:@49557.4]
  wire [9:0] _T_6220; // @[Mux.scala 31:69:@49558.4]
  wire [9:0] _T_6221; // @[Mux.scala 31:69:@49559.4]
  wire [9:0] _T_6222; // @[Mux.scala 31:69:@49560.4]
  wire [9:0] _T_6223; // @[Mux.scala 31:69:@49561.4]
  wire  _T_6231; // @[MemPrimitives.scala 110:228:@49570.4]
  wire  _T_6237; // @[MemPrimitives.scala 110:228:@49574.4]
  wire  _T_6243; // @[MemPrimitives.scala 110:228:@49578.4]
  wire  _T_6249; // @[MemPrimitives.scala 110:228:@49582.4]
  wire  _T_6255; // @[MemPrimitives.scala 110:228:@49586.4]
  wire  _T_6261; // @[MemPrimitives.scala 110:228:@49590.4]
  wire  _T_6267; // @[MemPrimitives.scala 110:228:@49594.4]
  wire  _T_6273; // @[MemPrimitives.scala 110:228:@49598.4]
  wire  _T_6279; // @[MemPrimitives.scala 110:228:@49602.4]
  wire  _T_6285; // @[MemPrimitives.scala 110:228:@49606.4]
  wire  _T_6291; // @[MemPrimitives.scala 110:228:@49610.4]
  wire  _T_6297; // @[MemPrimitives.scala 110:228:@49614.4]
  wire  _T_6303; // @[MemPrimitives.scala 110:228:@49618.4]
  wire  _T_6309; // @[MemPrimitives.scala 110:228:@49622.4]
  wire  _T_6315; // @[MemPrimitives.scala 110:228:@49626.4]
  wire  _T_6317; // @[MemPrimitives.scala 123:41:@49646.4]
  wire  _T_6318; // @[MemPrimitives.scala 123:41:@49647.4]
  wire  _T_6319; // @[MemPrimitives.scala 123:41:@49648.4]
  wire  _T_6320; // @[MemPrimitives.scala 123:41:@49649.4]
  wire  _T_6321; // @[MemPrimitives.scala 123:41:@49650.4]
  wire  _T_6322; // @[MemPrimitives.scala 123:41:@49651.4]
  wire  _T_6323; // @[MemPrimitives.scala 123:41:@49652.4]
  wire  _T_6324; // @[MemPrimitives.scala 123:41:@49653.4]
  wire  _T_6325; // @[MemPrimitives.scala 123:41:@49654.4]
  wire  _T_6326; // @[MemPrimitives.scala 123:41:@49655.4]
  wire  _T_6327; // @[MemPrimitives.scala 123:41:@49656.4]
  wire  _T_6328; // @[MemPrimitives.scala 123:41:@49657.4]
  wire  _T_6329; // @[MemPrimitives.scala 123:41:@49658.4]
  wire  _T_6330; // @[MemPrimitives.scala 123:41:@49659.4]
  wire  _T_6331; // @[MemPrimitives.scala 123:41:@49660.4]
  wire [9:0] _T_6333; // @[Cat.scala 30:58:@49662.4]
  wire [9:0] _T_6335; // @[Cat.scala 30:58:@49664.4]
  wire [9:0] _T_6337; // @[Cat.scala 30:58:@49666.4]
  wire [9:0] _T_6339; // @[Cat.scala 30:58:@49668.4]
  wire [9:0] _T_6341; // @[Cat.scala 30:58:@49670.4]
  wire [9:0] _T_6343; // @[Cat.scala 30:58:@49672.4]
  wire [9:0] _T_6345; // @[Cat.scala 30:58:@49674.4]
  wire [9:0] _T_6347; // @[Cat.scala 30:58:@49676.4]
  wire [9:0] _T_6349; // @[Cat.scala 30:58:@49678.4]
  wire [9:0] _T_6351; // @[Cat.scala 30:58:@49680.4]
  wire [9:0] _T_6353; // @[Cat.scala 30:58:@49682.4]
  wire [9:0] _T_6355; // @[Cat.scala 30:58:@49684.4]
  wire [9:0] _T_6357; // @[Cat.scala 30:58:@49686.4]
  wire [9:0] _T_6359; // @[Cat.scala 30:58:@49688.4]
  wire [9:0] _T_6361; // @[Cat.scala 30:58:@49690.4]
  wire [9:0] _T_6362; // @[Mux.scala 31:69:@49691.4]
  wire [9:0] _T_6363; // @[Mux.scala 31:69:@49692.4]
  wire [9:0] _T_6364; // @[Mux.scala 31:69:@49693.4]
  wire [9:0] _T_6365; // @[Mux.scala 31:69:@49694.4]
  wire [9:0] _T_6366; // @[Mux.scala 31:69:@49695.4]
  wire [9:0] _T_6367; // @[Mux.scala 31:69:@49696.4]
  wire [9:0] _T_6368; // @[Mux.scala 31:69:@49697.4]
  wire [9:0] _T_6369; // @[Mux.scala 31:69:@49698.4]
  wire [9:0] _T_6370; // @[Mux.scala 31:69:@49699.4]
  wire [9:0] _T_6371; // @[Mux.scala 31:69:@49700.4]
  wire [9:0] _T_6372; // @[Mux.scala 31:69:@49701.4]
  wire [9:0] _T_6373; // @[Mux.scala 31:69:@49702.4]
  wire [9:0] _T_6374; // @[Mux.scala 31:69:@49703.4]
  wire [9:0] _T_6375; // @[Mux.scala 31:69:@49704.4]
  wire  _T_6383; // @[MemPrimitives.scala 110:228:@49713.4]
  wire  _T_6389; // @[MemPrimitives.scala 110:228:@49717.4]
  wire  _T_6395; // @[MemPrimitives.scala 110:228:@49721.4]
  wire  _T_6401; // @[MemPrimitives.scala 110:228:@49725.4]
  wire  _T_6407; // @[MemPrimitives.scala 110:228:@49729.4]
  wire  _T_6413; // @[MemPrimitives.scala 110:228:@49733.4]
  wire  _T_6419; // @[MemPrimitives.scala 110:228:@49737.4]
  wire  _T_6425; // @[MemPrimitives.scala 110:228:@49741.4]
  wire  _T_6431; // @[MemPrimitives.scala 110:228:@49745.4]
  wire  _T_6437; // @[MemPrimitives.scala 110:228:@49749.4]
  wire  _T_6443; // @[MemPrimitives.scala 110:228:@49753.4]
  wire  _T_6449; // @[MemPrimitives.scala 110:228:@49757.4]
  wire  _T_6455; // @[MemPrimitives.scala 110:228:@49761.4]
  wire  _T_6461; // @[MemPrimitives.scala 110:228:@49765.4]
  wire  _T_6467; // @[MemPrimitives.scala 110:228:@49769.4]
  wire  _T_6469; // @[MemPrimitives.scala 123:41:@49789.4]
  wire  _T_6470; // @[MemPrimitives.scala 123:41:@49790.4]
  wire  _T_6471; // @[MemPrimitives.scala 123:41:@49791.4]
  wire  _T_6472; // @[MemPrimitives.scala 123:41:@49792.4]
  wire  _T_6473; // @[MemPrimitives.scala 123:41:@49793.4]
  wire  _T_6474; // @[MemPrimitives.scala 123:41:@49794.4]
  wire  _T_6475; // @[MemPrimitives.scala 123:41:@49795.4]
  wire  _T_6476; // @[MemPrimitives.scala 123:41:@49796.4]
  wire  _T_6477; // @[MemPrimitives.scala 123:41:@49797.4]
  wire  _T_6478; // @[MemPrimitives.scala 123:41:@49798.4]
  wire  _T_6479; // @[MemPrimitives.scala 123:41:@49799.4]
  wire  _T_6480; // @[MemPrimitives.scala 123:41:@49800.4]
  wire  _T_6481; // @[MemPrimitives.scala 123:41:@49801.4]
  wire  _T_6482; // @[MemPrimitives.scala 123:41:@49802.4]
  wire  _T_6483; // @[MemPrimitives.scala 123:41:@49803.4]
  wire [9:0] _T_6485; // @[Cat.scala 30:58:@49805.4]
  wire [9:0] _T_6487; // @[Cat.scala 30:58:@49807.4]
  wire [9:0] _T_6489; // @[Cat.scala 30:58:@49809.4]
  wire [9:0] _T_6491; // @[Cat.scala 30:58:@49811.4]
  wire [9:0] _T_6493; // @[Cat.scala 30:58:@49813.4]
  wire [9:0] _T_6495; // @[Cat.scala 30:58:@49815.4]
  wire [9:0] _T_6497; // @[Cat.scala 30:58:@49817.4]
  wire [9:0] _T_6499; // @[Cat.scala 30:58:@49819.4]
  wire [9:0] _T_6501; // @[Cat.scala 30:58:@49821.4]
  wire [9:0] _T_6503; // @[Cat.scala 30:58:@49823.4]
  wire [9:0] _T_6505; // @[Cat.scala 30:58:@49825.4]
  wire [9:0] _T_6507; // @[Cat.scala 30:58:@49827.4]
  wire [9:0] _T_6509; // @[Cat.scala 30:58:@49829.4]
  wire [9:0] _T_6511; // @[Cat.scala 30:58:@49831.4]
  wire [9:0] _T_6513; // @[Cat.scala 30:58:@49833.4]
  wire [9:0] _T_6514; // @[Mux.scala 31:69:@49834.4]
  wire [9:0] _T_6515; // @[Mux.scala 31:69:@49835.4]
  wire [9:0] _T_6516; // @[Mux.scala 31:69:@49836.4]
  wire [9:0] _T_6517; // @[Mux.scala 31:69:@49837.4]
  wire [9:0] _T_6518; // @[Mux.scala 31:69:@49838.4]
  wire [9:0] _T_6519; // @[Mux.scala 31:69:@49839.4]
  wire [9:0] _T_6520; // @[Mux.scala 31:69:@49840.4]
  wire [9:0] _T_6521; // @[Mux.scala 31:69:@49841.4]
  wire [9:0] _T_6522; // @[Mux.scala 31:69:@49842.4]
  wire [9:0] _T_6523; // @[Mux.scala 31:69:@49843.4]
  wire [9:0] _T_6524; // @[Mux.scala 31:69:@49844.4]
  wire [9:0] _T_6525; // @[Mux.scala 31:69:@49845.4]
  wire [9:0] _T_6526; // @[Mux.scala 31:69:@49846.4]
  wire [9:0] _T_6527; // @[Mux.scala 31:69:@49847.4]
  wire  _T_6535; // @[MemPrimitives.scala 110:228:@49856.4]
  wire  _T_6541; // @[MemPrimitives.scala 110:228:@49860.4]
  wire  _T_6547; // @[MemPrimitives.scala 110:228:@49864.4]
  wire  _T_6553; // @[MemPrimitives.scala 110:228:@49868.4]
  wire  _T_6559; // @[MemPrimitives.scala 110:228:@49872.4]
  wire  _T_6565; // @[MemPrimitives.scala 110:228:@49876.4]
  wire  _T_6571; // @[MemPrimitives.scala 110:228:@49880.4]
  wire  _T_6577; // @[MemPrimitives.scala 110:228:@49884.4]
  wire  _T_6583; // @[MemPrimitives.scala 110:228:@49888.4]
  wire  _T_6589; // @[MemPrimitives.scala 110:228:@49892.4]
  wire  _T_6595; // @[MemPrimitives.scala 110:228:@49896.4]
  wire  _T_6601; // @[MemPrimitives.scala 110:228:@49900.4]
  wire  _T_6607; // @[MemPrimitives.scala 110:228:@49904.4]
  wire  _T_6613; // @[MemPrimitives.scala 110:228:@49908.4]
  wire  _T_6619; // @[MemPrimitives.scala 110:228:@49912.4]
  wire  _T_6621; // @[MemPrimitives.scala 123:41:@49932.4]
  wire  _T_6622; // @[MemPrimitives.scala 123:41:@49933.4]
  wire  _T_6623; // @[MemPrimitives.scala 123:41:@49934.4]
  wire  _T_6624; // @[MemPrimitives.scala 123:41:@49935.4]
  wire  _T_6625; // @[MemPrimitives.scala 123:41:@49936.4]
  wire  _T_6626; // @[MemPrimitives.scala 123:41:@49937.4]
  wire  _T_6627; // @[MemPrimitives.scala 123:41:@49938.4]
  wire  _T_6628; // @[MemPrimitives.scala 123:41:@49939.4]
  wire  _T_6629; // @[MemPrimitives.scala 123:41:@49940.4]
  wire  _T_6630; // @[MemPrimitives.scala 123:41:@49941.4]
  wire  _T_6631; // @[MemPrimitives.scala 123:41:@49942.4]
  wire  _T_6632; // @[MemPrimitives.scala 123:41:@49943.4]
  wire  _T_6633; // @[MemPrimitives.scala 123:41:@49944.4]
  wire  _T_6634; // @[MemPrimitives.scala 123:41:@49945.4]
  wire  _T_6635; // @[MemPrimitives.scala 123:41:@49946.4]
  wire [9:0] _T_6637; // @[Cat.scala 30:58:@49948.4]
  wire [9:0] _T_6639; // @[Cat.scala 30:58:@49950.4]
  wire [9:0] _T_6641; // @[Cat.scala 30:58:@49952.4]
  wire [9:0] _T_6643; // @[Cat.scala 30:58:@49954.4]
  wire [9:0] _T_6645; // @[Cat.scala 30:58:@49956.4]
  wire [9:0] _T_6647; // @[Cat.scala 30:58:@49958.4]
  wire [9:0] _T_6649; // @[Cat.scala 30:58:@49960.4]
  wire [9:0] _T_6651; // @[Cat.scala 30:58:@49962.4]
  wire [9:0] _T_6653; // @[Cat.scala 30:58:@49964.4]
  wire [9:0] _T_6655; // @[Cat.scala 30:58:@49966.4]
  wire [9:0] _T_6657; // @[Cat.scala 30:58:@49968.4]
  wire [9:0] _T_6659; // @[Cat.scala 30:58:@49970.4]
  wire [9:0] _T_6661; // @[Cat.scala 30:58:@49972.4]
  wire [9:0] _T_6663; // @[Cat.scala 30:58:@49974.4]
  wire [9:0] _T_6665; // @[Cat.scala 30:58:@49976.4]
  wire [9:0] _T_6666; // @[Mux.scala 31:69:@49977.4]
  wire [9:0] _T_6667; // @[Mux.scala 31:69:@49978.4]
  wire [9:0] _T_6668; // @[Mux.scala 31:69:@49979.4]
  wire [9:0] _T_6669; // @[Mux.scala 31:69:@49980.4]
  wire [9:0] _T_6670; // @[Mux.scala 31:69:@49981.4]
  wire [9:0] _T_6671; // @[Mux.scala 31:69:@49982.4]
  wire [9:0] _T_6672; // @[Mux.scala 31:69:@49983.4]
  wire [9:0] _T_6673; // @[Mux.scala 31:69:@49984.4]
  wire [9:0] _T_6674; // @[Mux.scala 31:69:@49985.4]
  wire [9:0] _T_6675; // @[Mux.scala 31:69:@49986.4]
  wire [9:0] _T_6676; // @[Mux.scala 31:69:@49987.4]
  wire [9:0] _T_6677; // @[Mux.scala 31:69:@49988.4]
  wire [9:0] _T_6678; // @[Mux.scala 31:69:@49989.4]
  wire [9:0] _T_6679; // @[Mux.scala 31:69:@49990.4]
  wire  _T_6687; // @[MemPrimitives.scala 110:228:@49999.4]
  wire  _T_6693; // @[MemPrimitives.scala 110:228:@50003.4]
  wire  _T_6699; // @[MemPrimitives.scala 110:228:@50007.4]
  wire  _T_6705; // @[MemPrimitives.scala 110:228:@50011.4]
  wire  _T_6711; // @[MemPrimitives.scala 110:228:@50015.4]
  wire  _T_6717; // @[MemPrimitives.scala 110:228:@50019.4]
  wire  _T_6723; // @[MemPrimitives.scala 110:228:@50023.4]
  wire  _T_6729; // @[MemPrimitives.scala 110:228:@50027.4]
  wire  _T_6735; // @[MemPrimitives.scala 110:228:@50031.4]
  wire  _T_6741; // @[MemPrimitives.scala 110:228:@50035.4]
  wire  _T_6747; // @[MemPrimitives.scala 110:228:@50039.4]
  wire  _T_6753; // @[MemPrimitives.scala 110:228:@50043.4]
  wire  _T_6759; // @[MemPrimitives.scala 110:228:@50047.4]
  wire  _T_6765; // @[MemPrimitives.scala 110:228:@50051.4]
  wire  _T_6771; // @[MemPrimitives.scala 110:228:@50055.4]
  wire  _T_6773; // @[MemPrimitives.scala 123:41:@50075.4]
  wire  _T_6774; // @[MemPrimitives.scala 123:41:@50076.4]
  wire  _T_6775; // @[MemPrimitives.scala 123:41:@50077.4]
  wire  _T_6776; // @[MemPrimitives.scala 123:41:@50078.4]
  wire  _T_6777; // @[MemPrimitives.scala 123:41:@50079.4]
  wire  _T_6778; // @[MemPrimitives.scala 123:41:@50080.4]
  wire  _T_6779; // @[MemPrimitives.scala 123:41:@50081.4]
  wire  _T_6780; // @[MemPrimitives.scala 123:41:@50082.4]
  wire  _T_6781; // @[MemPrimitives.scala 123:41:@50083.4]
  wire  _T_6782; // @[MemPrimitives.scala 123:41:@50084.4]
  wire  _T_6783; // @[MemPrimitives.scala 123:41:@50085.4]
  wire  _T_6784; // @[MemPrimitives.scala 123:41:@50086.4]
  wire  _T_6785; // @[MemPrimitives.scala 123:41:@50087.4]
  wire  _T_6786; // @[MemPrimitives.scala 123:41:@50088.4]
  wire  _T_6787; // @[MemPrimitives.scala 123:41:@50089.4]
  wire [9:0] _T_6789; // @[Cat.scala 30:58:@50091.4]
  wire [9:0] _T_6791; // @[Cat.scala 30:58:@50093.4]
  wire [9:0] _T_6793; // @[Cat.scala 30:58:@50095.4]
  wire [9:0] _T_6795; // @[Cat.scala 30:58:@50097.4]
  wire [9:0] _T_6797; // @[Cat.scala 30:58:@50099.4]
  wire [9:0] _T_6799; // @[Cat.scala 30:58:@50101.4]
  wire [9:0] _T_6801; // @[Cat.scala 30:58:@50103.4]
  wire [9:0] _T_6803; // @[Cat.scala 30:58:@50105.4]
  wire [9:0] _T_6805; // @[Cat.scala 30:58:@50107.4]
  wire [9:0] _T_6807; // @[Cat.scala 30:58:@50109.4]
  wire [9:0] _T_6809; // @[Cat.scala 30:58:@50111.4]
  wire [9:0] _T_6811; // @[Cat.scala 30:58:@50113.4]
  wire [9:0] _T_6813; // @[Cat.scala 30:58:@50115.4]
  wire [9:0] _T_6815; // @[Cat.scala 30:58:@50117.4]
  wire [9:0] _T_6817; // @[Cat.scala 30:58:@50119.4]
  wire [9:0] _T_6818; // @[Mux.scala 31:69:@50120.4]
  wire [9:0] _T_6819; // @[Mux.scala 31:69:@50121.4]
  wire [9:0] _T_6820; // @[Mux.scala 31:69:@50122.4]
  wire [9:0] _T_6821; // @[Mux.scala 31:69:@50123.4]
  wire [9:0] _T_6822; // @[Mux.scala 31:69:@50124.4]
  wire [9:0] _T_6823; // @[Mux.scala 31:69:@50125.4]
  wire [9:0] _T_6824; // @[Mux.scala 31:69:@50126.4]
  wire [9:0] _T_6825; // @[Mux.scala 31:69:@50127.4]
  wire [9:0] _T_6826; // @[Mux.scala 31:69:@50128.4]
  wire [9:0] _T_6827; // @[Mux.scala 31:69:@50129.4]
  wire [9:0] _T_6828; // @[Mux.scala 31:69:@50130.4]
  wire [9:0] _T_6829; // @[Mux.scala 31:69:@50131.4]
  wire [9:0] _T_6830; // @[Mux.scala 31:69:@50132.4]
  wire [9:0] _T_6831; // @[Mux.scala 31:69:@50133.4]
  wire  _T_6839; // @[MemPrimitives.scala 110:228:@50142.4]
  wire  _T_6845; // @[MemPrimitives.scala 110:228:@50146.4]
  wire  _T_6851; // @[MemPrimitives.scala 110:228:@50150.4]
  wire  _T_6857; // @[MemPrimitives.scala 110:228:@50154.4]
  wire  _T_6863; // @[MemPrimitives.scala 110:228:@50158.4]
  wire  _T_6869; // @[MemPrimitives.scala 110:228:@50162.4]
  wire  _T_6875; // @[MemPrimitives.scala 110:228:@50166.4]
  wire  _T_6881; // @[MemPrimitives.scala 110:228:@50170.4]
  wire  _T_6887; // @[MemPrimitives.scala 110:228:@50174.4]
  wire  _T_6893; // @[MemPrimitives.scala 110:228:@50178.4]
  wire  _T_6899; // @[MemPrimitives.scala 110:228:@50182.4]
  wire  _T_6905; // @[MemPrimitives.scala 110:228:@50186.4]
  wire  _T_6911; // @[MemPrimitives.scala 110:228:@50190.4]
  wire  _T_6917; // @[MemPrimitives.scala 110:228:@50194.4]
  wire  _T_6923; // @[MemPrimitives.scala 110:228:@50198.4]
  wire  _T_6925; // @[MemPrimitives.scala 123:41:@50218.4]
  wire  _T_6926; // @[MemPrimitives.scala 123:41:@50219.4]
  wire  _T_6927; // @[MemPrimitives.scala 123:41:@50220.4]
  wire  _T_6928; // @[MemPrimitives.scala 123:41:@50221.4]
  wire  _T_6929; // @[MemPrimitives.scala 123:41:@50222.4]
  wire  _T_6930; // @[MemPrimitives.scala 123:41:@50223.4]
  wire  _T_6931; // @[MemPrimitives.scala 123:41:@50224.4]
  wire  _T_6932; // @[MemPrimitives.scala 123:41:@50225.4]
  wire  _T_6933; // @[MemPrimitives.scala 123:41:@50226.4]
  wire  _T_6934; // @[MemPrimitives.scala 123:41:@50227.4]
  wire  _T_6935; // @[MemPrimitives.scala 123:41:@50228.4]
  wire  _T_6936; // @[MemPrimitives.scala 123:41:@50229.4]
  wire  _T_6937; // @[MemPrimitives.scala 123:41:@50230.4]
  wire  _T_6938; // @[MemPrimitives.scala 123:41:@50231.4]
  wire  _T_6939; // @[MemPrimitives.scala 123:41:@50232.4]
  wire [9:0] _T_6941; // @[Cat.scala 30:58:@50234.4]
  wire [9:0] _T_6943; // @[Cat.scala 30:58:@50236.4]
  wire [9:0] _T_6945; // @[Cat.scala 30:58:@50238.4]
  wire [9:0] _T_6947; // @[Cat.scala 30:58:@50240.4]
  wire [9:0] _T_6949; // @[Cat.scala 30:58:@50242.4]
  wire [9:0] _T_6951; // @[Cat.scala 30:58:@50244.4]
  wire [9:0] _T_6953; // @[Cat.scala 30:58:@50246.4]
  wire [9:0] _T_6955; // @[Cat.scala 30:58:@50248.4]
  wire [9:0] _T_6957; // @[Cat.scala 30:58:@50250.4]
  wire [9:0] _T_6959; // @[Cat.scala 30:58:@50252.4]
  wire [9:0] _T_6961; // @[Cat.scala 30:58:@50254.4]
  wire [9:0] _T_6963; // @[Cat.scala 30:58:@50256.4]
  wire [9:0] _T_6965; // @[Cat.scala 30:58:@50258.4]
  wire [9:0] _T_6967; // @[Cat.scala 30:58:@50260.4]
  wire [9:0] _T_6969; // @[Cat.scala 30:58:@50262.4]
  wire [9:0] _T_6970; // @[Mux.scala 31:69:@50263.4]
  wire [9:0] _T_6971; // @[Mux.scala 31:69:@50264.4]
  wire [9:0] _T_6972; // @[Mux.scala 31:69:@50265.4]
  wire [9:0] _T_6973; // @[Mux.scala 31:69:@50266.4]
  wire [9:0] _T_6974; // @[Mux.scala 31:69:@50267.4]
  wire [9:0] _T_6975; // @[Mux.scala 31:69:@50268.4]
  wire [9:0] _T_6976; // @[Mux.scala 31:69:@50269.4]
  wire [9:0] _T_6977; // @[Mux.scala 31:69:@50270.4]
  wire [9:0] _T_6978; // @[Mux.scala 31:69:@50271.4]
  wire [9:0] _T_6979; // @[Mux.scala 31:69:@50272.4]
  wire [9:0] _T_6980; // @[Mux.scala 31:69:@50273.4]
  wire [9:0] _T_6981; // @[Mux.scala 31:69:@50274.4]
  wire [9:0] _T_6982; // @[Mux.scala 31:69:@50275.4]
  wire [9:0] _T_6983; // @[Mux.scala 31:69:@50276.4]
  wire  _T_6991; // @[MemPrimitives.scala 110:228:@50285.4]
  wire  _T_6997; // @[MemPrimitives.scala 110:228:@50289.4]
  wire  _T_7003; // @[MemPrimitives.scala 110:228:@50293.4]
  wire  _T_7009; // @[MemPrimitives.scala 110:228:@50297.4]
  wire  _T_7015; // @[MemPrimitives.scala 110:228:@50301.4]
  wire  _T_7021; // @[MemPrimitives.scala 110:228:@50305.4]
  wire  _T_7027; // @[MemPrimitives.scala 110:228:@50309.4]
  wire  _T_7033; // @[MemPrimitives.scala 110:228:@50313.4]
  wire  _T_7039; // @[MemPrimitives.scala 110:228:@50317.4]
  wire  _T_7045; // @[MemPrimitives.scala 110:228:@50321.4]
  wire  _T_7051; // @[MemPrimitives.scala 110:228:@50325.4]
  wire  _T_7057; // @[MemPrimitives.scala 110:228:@50329.4]
  wire  _T_7063; // @[MemPrimitives.scala 110:228:@50333.4]
  wire  _T_7069; // @[MemPrimitives.scala 110:228:@50337.4]
  wire  _T_7075; // @[MemPrimitives.scala 110:228:@50341.4]
  wire  _T_7077; // @[MemPrimitives.scala 123:41:@50361.4]
  wire  _T_7078; // @[MemPrimitives.scala 123:41:@50362.4]
  wire  _T_7079; // @[MemPrimitives.scala 123:41:@50363.4]
  wire  _T_7080; // @[MemPrimitives.scala 123:41:@50364.4]
  wire  _T_7081; // @[MemPrimitives.scala 123:41:@50365.4]
  wire  _T_7082; // @[MemPrimitives.scala 123:41:@50366.4]
  wire  _T_7083; // @[MemPrimitives.scala 123:41:@50367.4]
  wire  _T_7084; // @[MemPrimitives.scala 123:41:@50368.4]
  wire  _T_7085; // @[MemPrimitives.scala 123:41:@50369.4]
  wire  _T_7086; // @[MemPrimitives.scala 123:41:@50370.4]
  wire  _T_7087; // @[MemPrimitives.scala 123:41:@50371.4]
  wire  _T_7088; // @[MemPrimitives.scala 123:41:@50372.4]
  wire  _T_7089; // @[MemPrimitives.scala 123:41:@50373.4]
  wire  _T_7090; // @[MemPrimitives.scala 123:41:@50374.4]
  wire  _T_7091; // @[MemPrimitives.scala 123:41:@50375.4]
  wire [9:0] _T_7093; // @[Cat.scala 30:58:@50377.4]
  wire [9:0] _T_7095; // @[Cat.scala 30:58:@50379.4]
  wire [9:0] _T_7097; // @[Cat.scala 30:58:@50381.4]
  wire [9:0] _T_7099; // @[Cat.scala 30:58:@50383.4]
  wire [9:0] _T_7101; // @[Cat.scala 30:58:@50385.4]
  wire [9:0] _T_7103; // @[Cat.scala 30:58:@50387.4]
  wire [9:0] _T_7105; // @[Cat.scala 30:58:@50389.4]
  wire [9:0] _T_7107; // @[Cat.scala 30:58:@50391.4]
  wire [9:0] _T_7109; // @[Cat.scala 30:58:@50393.4]
  wire [9:0] _T_7111; // @[Cat.scala 30:58:@50395.4]
  wire [9:0] _T_7113; // @[Cat.scala 30:58:@50397.4]
  wire [9:0] _T_7115; // @[Cat.scala 30:58:@50399.4]
  wire [9:0] _T_7117; // @[Cat.scala 30:58:@50401.4]
  wire [9:0] _T_7119; // @[Cat.scala 30:58:@50403.4]
  wire [9:0] _T_7121; // @[Cat.scala 30:58:@50405.4]
  wire [9:0] _T_7122; // @[Mux.scala 31:69:@50406.4]
  wire [9:0] _T_7123; // @[Mux.scala 31:69:@50407.4]
  wire [9:0] _T_7124; // @[Mux.scala 31:69:@50408.4]
  wire [9:0] _T_7125; // @[Mux.scala 31:69:@50409.4]
  wire [9:0] _T_7126; // @[Mux.scala 31:69:@50410.4]
  wire [9:0] _T_7127; // @[Mux.scala 31:69:@50411.4]
  wire [9:0] _T_7128; // @[Mux.scala 31:69:@50412.4]
  wire [9:0] _T_7129; // @[Mux.scala 31:69:@50413.4]
  wire [9:0] _T_7130; // @[Mux.scala 31:69:@50414.4]
  wire [9:0] _T_7131; // @[Mux.scala 31:69:@50415.4]
  wire [9:0] _T_7132; // @[Mux.scala 31:69:@50416.4]
  wire [9:0] _T_7133; // @[Mux.scala 31:69:@50417.4]
  wire [9:0] _T_7134; // @[Mux.scala 31:69:@50418.4]
  wire [9:0] _T_7135; // @[Mux.scala 31:69:@50419.4]
  wire  _T_7143; // @[MemPrimitives.scala 110:228:@50428.4]
  wire  _T_7149; // @[MemPrimitives.scala 110:228:@50432.4]
  wire  _T_7155; // @[MemPrimitives.scala 110:228:@50436.4]
  wire  _T_7161; // @[MemPrimitives.scala 110:228:@50440.4]
  wire  _T_7167; // @[MemPrimitives.scala 110:228:@50444.4]
  wire  _T_7173; // @[MemPrimitives.scala 110:228:@50448.4]
  wire  _T_7179; // @[MemPrimitives.scala 110:228:@50452.4]
  wire  _T_7185; // @[MemPrimitives.scala 110:228:@50456.4]
  wire  _T_7191; // @[MemPrimitives.scala 110:228:@50460.4]
  wire  _T_7197; // @[MemPrimitives.scala 110:228:@50464.4]
  wire  _T_7203; // @[MemPrimitives.scala 110:228:@50468.4]
  wire  _T_7209; // @[MemPrimitives.scala 110:228:@50472.4]
  wire  _T_7215; // @[MemPrimitives.scala 110:228:@50476.4]
  wire  _T_7221; // @[MemPrimitives.scala 110:228:@50480.4]
  wire  _T_7227; // @[MemPrimitives.scala 110:228:@50484.4]
  wire  _T_7229; // @[MemPrimitives.scala 123:41:@50504.4]
  wire  _T_7230; // @[MemPrimitives.scala 123:41:@50505.4]
  wire  _T_7231; // @[MemPrimitives.scala 123:41:@50506.4]
  wire  _T_7232; // @[MemPrimitives.scala 123:41:@50507.4]
  wire  _T_7233; // @[MemPrimitives.scala 123:41:@50508.4]
  wire  _T_7234; // @[MemPrimitives.scala 123:41:@50509.4]
  wire  _T_7235; // @[MemPrimitives.scala 123:41:@50510.4]
  wire  _T_7236; // @[MemPrimitives.scala 123:41:@50511.4]
  wire  _T_7237; // @[MemPrimitives.scala 123:41:@50512.4]
  wire  _T_7238; // @[MemPrimitives.scala 123:41:@50513.4]
  wire  _T_7239; // @[MemPrimitives.scala 123:41:@50514.4]
  wire  _T_7240; // @[MemPrimitives.scala 123:41:@50515.4]
  wire  _T_7241; // @[MemPrimitives.scala 123:41:@50516.4]
  wire  _T_7242; // @[MemPrimitives.scala 123:41:@50517.4]
  wire  _T_7243; // @[MemPrimitives.scala 123:41:@50518.4]
  wire [9:0] _T_7245; // @[Cat.scala 30:58:@50520.4]
  wire [9:0] _T_7247; // @[Cat.scala 30:58:@50522.4]
  wire [9:0] _T_7249; // @[Cat.scala 30:58:@50524.4]
  wire [9:0] _T_7251; // @[Cat.scala 30:58:@50526.4]
  wire [9:0] _T_7253; // @[Cat.scala 30:58:@50528.4]
  wire [9:0] _T_7255; // @[Cat.scala 30:58:@50530.4]
  wire [9:0] _T_7257; // @[Cat.scala 30:58:@50532.4]
  wire [9:0] _T_7259; // @[Cat.scala 30:58:@50534.4]
  wire [9:0] _T_7261; // @[Cat.scala 30:58:@50536.4]
  wire [9:0] _T_7263; // @[Cat.scala 30:58:@50538.4]
  wire [9:0] _T_7265; // @[Cat.scala 30:58:@50540.4]
  wire [9:0] _T_7267; // @[Cat.scala 30:58:@50542.4]
  wire [9:0] _T_7269; // @[Cat.scala 30:58:@50544.4]
  wire [9:0] _T_7271; // @[Cat.scala 30:58:@50546.4]
  wire [9:0] _T_7273; // @[Cat.scala 30:58:@50548.4]
  wire [9:0] _T_7274; // @[Mux.scala 31:69:@50549.4]
  wire [9:0] _T_7275; // @[Mux.scala 31:69:@50550.4]
  wire [9:0] _T_7276; // @[Mux.scala 31:69:@50551.4]
  wire [9:0] _T_7277; // @[Mux.scala 31:69:@50552.4]
  wire [9:0] _T_7278; // @[Mux.scala 31:69:@50553.4]
  wire [9:0] _T_7279; // @[Mux.scala 31:69:@50554.4]
  wire [9:0] _T_7280; // @[Mux.scala 31:69:@50555.4]
  wire [9:0] _T_7281; // @[Mux.scala 31:69:@50556.4]
  wire [9:0] _T_7282; // @[Mux.scala 31:69:@50557.4]
  wire [9:0] _T_7283; // @[Mux.scala 31:69:@50558.4]
  wire [9:0] _T_7284; // @[Mux.scala 31:69:@50559.4]
  wire [9:0] _T_7285; // @[Mux.scala 31:69:@50560.4]
  wire [9:0] _T_7286; // @[Mux.scala 31:69:@50561.4]
  wire [9:0] _T_7287; // @[Mux.scala 31:69:@50562.4]
  wire  _T_7292; // @[MemPrimitives.scala 110:210:@50569.4]
  wire  _T_7295; // @[MemPrimitives.scala 110:228:@50571.4]
  wire  _T_7298; // @[MemPrimitives.scala 110:210:@50573.4]
  wire  _T_7301; // @[MemPrimitives.scala 110:228:@50575.4]
  wire  _T_7304; // @[MemPrimitives.scala 110:210:@50577.4]
  wire  _T_7307; // @[MemPrimitives.scala 110:228:@50579.4]
  wire  _T_7310; // @[MemPrimitives.scala 110:210:@50581.4]
  wire  _T_7313; // @[MemPrimitives.scala 110:228:@50583.4]
  wire  _T_7316; // @[MemPrimitives.scala 110:210:@50585.4]
  wire  _T_7319; // @[MemPrimitives.scala 110:228:@50587.4]
  wire  _T_7322; // @[MemPrimitives.scala 110:210:@50589.4]
  wire  _T_7325; // @[MemPrimitives.scala 110:228:@50591.4]
  wire  _T_7328; // @[MemPrimitives.scala 110:210:@50593.4]
  wire  _T_7331; // @[MemPrimitives.scala 110:228:@50595.4]
  wire  _T_7334; // @[MemPrimitives.scala 110:210:@50597.4]
  wire  _T_7337; // @[MemPrimitives.scala 110:228:@50599.4]
  wire  _T_7340; // @[MemPrimitives.scala 110:210:@50601.4]
  wire  _T_7343; // @[MemPrimitives.scala 110:228:@50603.4]
  wire  _T_7346; // @[MemPrimitives.scala 110:210:@50605.4]
  wire  _T_7349; // @[MemPrimitives.scala 110:228:@50607.4]
  wire  _T_7352; // @[MemPrimitives.scala 110:210:@50609.4]
  wire  _T_7355; // @[MemPrimitives.scala 110:228:@50611.4]
  wire  _T_7358; // @[MemPrimitives.scala 110:210:@50613.4]
  wire  _T_7361; // @[MemPrimitives.scala 110:228:@50615.4]
  wire  _T_7364; // @[MemPrimitives.scala 110:210:@50617.4]
  wire  _T_7367; // @[MemPrimitives.scala 110:228:@50619.4]
  wire  _T_7370; // @[MemPrimitives.scala 110:210:@50621.4]
  wire  _T_7373; // @[MemPrimitives.scala 110:228:@50623.4]
  wire  _T_7376; // @[MemPrimitives.scala 110:210:@50625.4]
  wire  _T_7379; // @[MemPrimitives.scala 110:228:@50627.4]
  wire  _T_7381; // @[MemPrimitives.scala 123:41:@50647.4]
  wire  _T_7382; // @[MemPrimitives.scala 123:41:@50648.4]
  wire  _T_7383; // @[MemPrimitives.scala 123:41:@50649.4]
  wire  _T_7384; // @[MemPrimitives.scala 123:41:@50650.4]
  wire  _T_7385; // @[MemPrimitives.scala 123:41:@50651.4]
  wire  _T_7386; // @[MemPrimitives.scala 123:41:@50652.4]
  wire  _T_7387; // @[MemPrimitives.scala 123:41:@50653.4]
  wire  _T_7388; // @[MemPrimitives.scala 123:41:@50654.4]
  wire  _T_7389; // @[MemPrimitives.scala 123:41:@50655.4]
  wire  _T_7390; // @[MemPrimitives.scala 123:41:@50656.4]
  wire  _T_7391; // @[MemPrimitives.scala 123:41:@50657.4]
  wire  _T_7392; // @[MemPrimitives.scala 123:41:@50658.4]
  wire  _T_7393; // @[MemPrimitives.scala 123:41:@50659.4]
  wire  _T_7394; // @[MemPrimitives.scala 123:41:@50660.4]
  wire  _T_7395; // @[MemPrimitives.scala 123:41:@50661.4]
  wire [9:0] _T_7397; // @[Cat.scala 30:58:@50663.4]
  wire [9:0] _T_7399; // @[Cat.scala 30:58:@50665.4]
  wire [9:0] _T_7401; // @[Cat.scala 30:58:@50667.4]
  wire [9:0] _T_7403; // @[Cat.scala 30:58:@50669.4]
  wire [9:0] _T_7405; // @[Cat.scala 30:58:@50671.4]
  wire [9:0] _T_7407; // @[Cat.scala 30:58:@50673.4]
  wire [9:0] _T_7409; // @[Cat.scala 30:58:@50675.4]
  wire [9:0] _T_7411; // @[Cat.scala 30:58:@50677.4]
  wire [9:0] _T_7413; // @[Cat.scala 30:58:@50679.4]
  wire [9:0] _T_7415; // @[Cat.scala 30:58:@50681.4]
  wire [9:0] _T_7417; // @[Cat.scala 30:58:@50683.4]
  wire [9:0] _T_7419; // @[Cat.scala 30:58:@50685.4]
  wire [9:0] _T_7421; // @[Cat.scala 30:58:@50687.4]
  wire [9:0] _T_7423; // @[Cat.scala 30:58:@50689.4]
  wire [9:0] _T_7425; // @[Cat.scala 30:58:@50691.4]
  wire [9:0] _T_7426; // @[Mux.scala 31:69:@50692.4]
  wire [9:0] _T_7427; // @[Mux.scala 31:69:@50693.4]
  wire [9:0] _T_7428; // @[Mux.scala 31:69:@50694.4]
  wire [9:0] _T_7429; // @[Mux.scala 31:69:@50695.4]
  wire [9:0] _T_7430; // @[Mux.scala 31:69:@50696.4]
  wire [9:0] _T_7431; // @[Mux.scala 31:69:@50697.4]
  wire [9:0] _T_7432; // @[Mux.scala 31:69:@50698.4]
  wire [9:0] _T_7433; // @[Mux.scala 31:69:@50699.4]
  wire [9:0] _T_7434; // @[Mux.scala 31:69:@50700.4]
  wire [9:0] _T_7435; // @[Mux.scala 31:69:@50701.4]
  wire [9:0] _T_7436; // @[Mux.scala 31:69:@50702.4]
  wire [9:0] _T_7437; // @[Mux.scala 31:69:@50703.4]
  wire [9:0] _T_7438; // @[Mux.scala 31:69:@50704.4]
  wire [9:0] _T_7439; // @[Mux.scala 31:69:@50705.4]
  wire  _T_7444; // @[MemPrimitives.scala 110:210:@50712.4]
  wire  _T_7447; // @[MemPrimitives.scala 110:228:@50714.4]
  wire  _T_7450; // @[MemPrimitives.scala 110:210:@50716.4]
  wire  _T_7453; // @[MemPrimitives.scala 110:228:@50718.4]
  wire  _T_7456; // @[MemPrimitives.scala 110:210:@50720.4]
  wire  _T_7459; // @[MemPrimitives.scala 110:228:@50722.4]
  wire  _T_7462; // @[MemPrimitives.scala 110:210:@50724.4]
  wire  _T_7465; // @[MemPrimitives.scala 110:228:@50726.4]
  wire  _T_7468; // @[MemPrimitives.scala 110:210:@50728.4]
  wire  _T_7471; // @[MemPrimitives.scala 110:228:@50730.4]
  wire  _T_7474; // @[MemPrimitives.scala 110:210:@50732.4]
  wire  _T_7477; // @[MemPrimitives.scala 110:228:@50734.4]
  wire  _T_7480; // @[MemPrimitives.scala 110:210:@50736.4]
  wire  _T_7483; // @[MemPrimitives.scala 110:228:@50738.4]
  wire  _T_7486; // @[MemPrimitives.scala 110:210:@50740.4]
  wire  _T_7489; // @[MemPrimitives.scala 110:228:@50742.4]
  wire  _T_7492; // @[MemPrimitives.scala 110:210:@50744.4]
  wire  _T_7495; // @[MemPrimitives.scala 110:228:@50746.4]
  wire  _T_7498; // @[MemPrimitives.scala 110:210:@50748.4]
  wire  _T_7501; // @[MemPrimitives.scala 110:228:@50750.4]
  wire  _T_7504; // @[MemPrimitives.scala 110:210:@50752.4]
  wire  _T_7507; // @[MemPrimitives.scala 110:228:@50754.4]
  wire  _T_7510; // @[MemPrimitives.scala 110:210:@50756.4]
  wire  _T_7513; // @[MemPrimitives.scala 110:228:@50758.4]
  wire  _T_7516; // @[MemPrimitives.scala 110:210:@50760.4]
  wire  _T_7519; // @[MemPrimitives.scala 110:228:@50762.4]
  wire  _T_7522; // @[MemPrimitives.scala 110:210:@50764.4]
  wire  _T_7525; // @[MemPrimitives.scala 110:228:@50766.4]
  wire  _T_7528; // @[MemPrimitives.scala 110:210:@50768.4]
  wire  _T_7531; // @[MemPrimitives.scala 110:228:@50770.4]
  wire  _T_7533; // @[MemPrimitives.scala 123:41:@50790.4]
  wire  _T_7534; // @[MemPrimitives.scala 123:41:@50791.4]
  wire  _T_7535; // @[MemPrimitives.scala 123:41:@50792.4]
  wire  _T_7536; // @[MemPrimitives.scala 123:41:@50793.4]
  wire  _T_7537; // @[MemPrimitives.scala 123:41:@50794.4]
  wire  _T_7538; // @[MemPrimitives.scala 123:41:@50795.4]
  wire  _T_7539; // @[MemPrimitives.scala 123:41:@50796.4]
  wire  _T_7540; // @[MemPrimitives.scala 123:41:@50797.4]
  wire  _T_7541; // @[MemPrimitives.scala 123:41:@50798.4]
  wire  _T_7542; // @[MemPrimitives.scala 123:41:@50799.4]
  wire  _T_7543; // @[MemPrimitives.scala 123:41:@50800.4]
  wire  _T_7544; // @[MemPrimitives.scala 123:41:@50801.4]
  wire  _T_7545; // @[MemPrimitives.scala 123:41:@50802.4]
  wire  _T_7546; // @[MemPrimitives.scala 123:41:@50803.4]
  wire  _T_7547; // @[MemPrimitives.scala 123:41:@50804.4]
  wire [9:0] _T_7549; // @[Cat.scala 30:58:@50806.4]
  wire [9:0] _T_7551; // @[Cat.scala 30:58:@50808.4]
  wire [9:0] _T_7553; // @[Cat.scala 30:58:@50810.4]
  wire [9:0] _T_7555; // @[Cat.scala 30:58:@50812.4]
  wire [9:0] _T_7557; // @[Cat.scala 30:58:@50814.4]
  wire [9:0] _T_7559; // @[Cat.scala 30:58:@50816.4]
  wire [9:0] _T_7561; // @[Cat.scala 30:58:@50818.4]
  wire [9:0] _T_7563; // @[Cat.scala 30:58:@50820.4]
  wire [9:0] _T_7565; // @[Cat.scala 30:58:@50822.4]
  wire [9:0] _T_7567; // @[Cat.scala 30:58:@50824.4]
  wire [9:0] _T_7569; // @[Cat.scala 30:58:@50826.4]
  wire [9:0] _T_7571; // @[Cat.scala 30:58:@50828.4]
  wire [9:0] _T_7573; // @[Cat.scala 30:58:@50830.4]
  wire [9:0] _T_7575; // @[Cat.scala 30:58:@50832.4]
  wire [9:0] _T_7577; // @[Cat.scala 30:58:@50834.4]
  wire [9:0] _T_7578; // @[Mux.scala 31:69:@50835.4]
  wire [9:0] _T_7579; // @[Mux.scala 31:69:@50836.4]
  wire [9:0] _T_7580; // @[Mux.scala 31:69:@50837.4]
  wire [9:0] _T_7581; // @[Mux.scala 31:69:@50838.4]
  wire [9:0] _T_7582; // @[Mux.scala 31:69:@50839.4]
  wire [9:0] _T_7583; // @[Mux.scala 31:69:@50840.4]
  wire [9:0] _T_7584; // @[Mux.scala 31:69:@50841.4]
  wire [9:0] _T_7585; // @[Mux.scala 31:69:@50842.4]
  wire [9:0] _T_7586; // @[Mux.scala 31:69:@50843.4]
  wire [9:0] _T_7587; // @[Mux.scala 31:69:@50844.4]
  wire [9:0] _T_7588; // @[Mux.scala 31:69:@50845.4]
  wire [9:0] _T_7589; // @[Mux.scala 31:69:@50846.4]
  wire [9:0] _T_7590; // @[Mux.scala 31:69:@50847.4]
  wire [9:0] _T_7591; // @[Mux.scala 31:69:@50848.4]
  wire  _T_7599; // @[MemPrimitives.scala 110:228:@50857.4]
  wire  _T_7605; // @[MemPrimitives.scala 110:228:@50861.4]
  wire  _T_7611; // @[MemPrimitives.scala 110:228:@50865.4]
  wire  _T_7617; // @[MemPrimitives.scala 110:228:@50869.4]
  wire  _T_7623; // @[MemPrimitives.scala 110:228:@50873.4]
  wire  _T_7629; // @[MemPrimitives.scala 110:228:@50877.4]
  wire  _T_7635; // @[MemPrimitives.scala 110:228:@50881.4]
  wire  _T_7641; // @[MemPrimitives.scala 110:228:@50885.4]
  wire  _T_7647; // @[MemPrimitives.scala 110:228:@50889.4]
  wire  _T_7653; // @[MemPrimitives.scala 110:228:@50893.4]
  wire  _T_7659; // @[MemPrimitives.scala 110:228:@50897.4]
  wire  _T_7665; // @[MemPrimitives.scala 110:228:@50901.4]
  wire  _T_7671; // @[MemPrimitives.scala 110:228:@50905.4]
  wire  _T_7677; // @[MemPrimitives.scala 110:228:@50909.4]
  wire  _T_7683; // @[MemPrimitives.scala 110:228:@50913.4]
  wire  _T_7685; // @[MemPrimitives.scala 123:41:@50933.4]
  wire  _T_7686; // @[MemPrimitives.scala 123:41:@50934.4]
  wire  _T_7687; // @[MemPrimitives.scala 123:41:@50935.4]
  wire  _T_7688; // @[MemPrimitives.scala 123:41:@50936.4]
  wire  _T_7689; // @[MemPrimitives.scala 123:41:@50937.4]
  wire  _T_7690; // @[MemPrimitives.scala 123:41:@50938.4]
  wire  _T_7691; // @[MemPrimitives.scala 123:41:@50939.4]
  wire  _T_7692; // @[MemPrimitives.scala 123:41:@50940.4]
  wire  _T_7693; // @[MemPrimitives.scala 123:41:@50941.4]
  wire  _T_7694; // @[MemPrimitives.scala 123:41:@50942.4]
  wire  _T_7695; // @[MemPrimitives.scala 123:41:@50943.4]
  wire  _T_7696; // @[MemPrimitives.scala 123:41:@50944.4]
  wire  _T_7697; // @[MemPrimitives.scala 123:41:@50945.4]
  wire  _T_7698; // @[MemPrimitives.scala 123:41:@50946.4]
  wire  _T_7699; // @[MemPrimitives.scala 123:41:@50947.4]
  wire [9:0] _T_7701; // @[Cat.scala 30:58:@50949.4]
  wire [9:0] _T_7703; // @[Cat.scala 30:58:@50951.4]
  wire [9:0] _T_7705; // @[Cat.scala 30:58:@50953.4]
  wire [9:0] _T_7707; // @[Cat.scala 30:58:@50955.4]
  wire [9:0] _T_7709; // @[Cat.scala 30:58:@50957.4]
  wire [9:0] _T_7711; // @[Cat.scala 30:58:@50959.4]
  wire [9:0] _T_7713; // @[Cat.scala 30:58:@50961.4]
  wire [9:0] _T_7715; // @[Cat.scala 30:58:@50963.4]
  wire [9:0] _T_7717; // @[Cat.scala 30:58:@50965.4]
  wire [9:0] _T_7719; // @[Cat.scala 30:58:@50967.4]
  wire [9:0] _T_7721; // @[Cat.scala 30:58:@50969.4]
  wire [9:0] _T_7723; // @[Cat.scala 30:58:@50971.4]
  wire [9:0] _T_7725; // @[Cat.scala 30:58:@50973.4]
  wire [9:0] _T_7727; // @[Cat.scala 30:58:@50975.4]
  wire [9:0] _T_7729; // @[Cat.scala 30:58:@50977.4]
  wire [9:0] _T_7730; // @[Mux.scala 31:69:@50978.4]
  wire [9:0] _T_7731; // @[Mux.scala 31:69:@50979.4]
  wire [9:0] _T_7732; // @[Mux.scala 31:69:@50980.4]
  wire [9:0] _T_7733; // @[Mux.scala 31:69:@50981.4]
  wire [9:0] _T_7734; // @[Mux.scala 31:69:@50982.4]
  wire [9:0] _T_7735; // @[Mux.scala 31:69:@50983.4]
  wire [9:0] _T_7736; // @[Mux.scala 31:69:@50984.4]
  wire [9:0] _T_7737; // @[Mux.scala 31:69:@50985.4]
  wire [9:0] _T_7738; // @[Mux.scala 31:69:@50986.4]
  wire [9:0] _T_7739; // @[Mux.scala 31:69:@50987.4]
  wire [9:0] _T_7740; // @[Mux.scala 31:69:@50988.4]
  wire [9:0] _T_7741; // @[Mux.scala 31:69:@50989.4]
  wire [9:0] _T_7742; // @[Mux.scala 31:69:@50990.4]
  wire [9:0] _T_7743; // @[Mux.scala 31:69:@50991.4]
  wire  _T_7751; // @[MemPrimitives.scala 110:228:@51000.4]
  wire  _T_7757; // @[MemPrimitives.scala 110:228:@51004.4]
  wire  _T_7763; // @[MemPrimitives.scala 110:228:@51008.4]
  wire  _T_7769; // @[MemPrimitives.scala 110:228:@51012.4]
  wire  _T_7775; // @[MemPrimitives.scala 110:228:@51016.4]
  wire  _T_7781; // @[MemPrimitives.scala 110:228:@51020.4]
  wire  _T_7787; // @[MemPrimitives.scala 110:228:@51024.4]
  wire  _T_7793; // @[MemPrimitives.scala 110:228:@51028.4]
  wire  _T_7799; // @[MemPrimitives.scala 110:228:@51032.4]
  wire  _T_7805; // @[MemPrimitives.scala 110:228:@51036.4]
  wire  _T_7811; // @[MemPrimitives.scala 110:228:@51040.4]
  wire  _T_7817; // @[MemPrimitives.scala 110:228:@51044.4]
  wire  _T_7823; // @[MemPrimitives.scala 110:228:@51048.4]
  wire  _T_7829; // @[MemPrimitives.scala 110:228:@51052.4]
  wire  _T_7835; // @[MemPrimitives.scala 110:228:@51056.4]
  wire  _T_7837; // @[MemPrimitives.scala 123:41:@51076.4]
  wire  _T_7838; // @[MemPrimitives.scala 123:41:@51077.4]
  wire  _T_7839; // @[MemPrimitives.scala 123:41:@51078.4]
  wire  _T_7840; // @[MemPrimitives.scala 123:41:@51079.4]
  wire  _T_7841; // @[MemPrimitives.scala 123:41:@51080.4]
  wire  _T_7842; // @[MemPrimitives.scala 123:41:@51081.4]
  wire  _T_7843; // @[MemPrimitives.scala 123:41:@51082.4]
  wire  _T_7844; // @[MemPrimitives.scala 123:41:@51083.4]
  wire  _T_7845; // @[MemPrimitives.scala 123:41:@51084.4]
  wire  _T_7846; // @[MemPrimitives.scala 123:41:@51085.4]
  wire  _T_7847; // @[MemPrimitives.scala 123:41:@51086.4]
  wire  _T_7848; // @[MemPrimitives.scala 123:41:@51087.4]
  wire  _T_7849; // @[MemPrimitives.scala 123:41:@51088.4]
  wire  _T_7850; // @[MemPrimitives.scala 123:41:@51089.4]
  wire  _T_7851; // @[MemPrimitives.scala 123:41:@51090.4]
  wire [9:0] _T_7853; // @[Cat.scala 30:58:@51092.4]
  wire [9:0] _T_7855; // @[Cat.scala 30:58:@51094.4]
  wire [9:0] _T_7857; // @[Cat.scala 30:58:@51096.4]
  wire [9:0] _T_7859; // @[Cat.scala 30:58:@51098.4]
  wire [9:0] _T_7861; // @[Cat.scala 30:58:@51100.4]
  wire [9:0] _T_7863; // @[Cat.scala 30:58:@51102.4]
  wire [9:0] _T_7865; // @[Cat.scala 30:58:@51104.4]
  wire [9:0] _T_7867; // @[Cat.scala 30:58:@51106.4]
  wire [9:0] _T_7869; // @[Cat.scala 30:58:@51108.4]
  wire [9:0] _T_7871; // @[Cat.scala 30:58:@51110.4]
  wire [9:0] _T_7873; // @[Cat.scala 30:58:@51112.4]
  wire [9:0] _T_7875; // @[Cat.scala 30:58:@51114.4]
  wire [9:0] _T_7877; // @[Cat.scala 30:58:@51116.4]
  wire [9:0] _T_7879; // @[Cat.scala 30:58:@51118.4]
  wire [9:0] _T_7881; // @[Cat.scala 30:58:@51120.4]
  wire [9:0] _T_7882; // @[Mux.scala 31:69:@51121.4]
  wire [9:0] _T_7883; // @[Mux.scala 31:69:@51122.4]
  wire [9:0] _T_7884; // @[Mux.scala 31:69:@51123.4]
  wire [9:0] _T_7885; // @[Mux.scala 31:69:@51124.4]
  wire [9:0] _T_7886; // @[Mux.scala 31:69:@51125.4]
  wire [9:0] _T_7887; // @[Mux.scala 31:69:@51126.4]
  wire [9:0] _T_7888; // @[Mux.scala 31:69:@51127.4]
  wire [9:0] _T_7889; // @[Mux.scala 31:69:@51128.4]
  wire [9:0] _T_7890; // @[Mux.scala 31:69:@51129.4]
  wire [9:0] _T_7891; // @[Mux.scala 31:69:@51130.4]
  wire [9:0] _T_7892; // @[Mux.scala 31:69:@51131.4]
  wire [9:0] _T_7893; // @[Mux.scala 31:69:@51132.4]
  wire [9:0] _T_7894; // @[Mux.scala 31:69:@51133.4]
  wire [9:0] _T_7895; // @[Mux.scala 31:69:@51134.4]
  wire  _T_7903; // @[MemPrimitives.scala 110:228:@51143.4]
  wire  _T_7909; // @[MemPrimitives.scala 110:228:@51147.4]
  wire  _T_7915; // @[MemPrimitives.scala 110:228:@51151.4]
  wire  _T_7921; // @[MemPrimitives.scala 110:228:@51155.4]
  wire  _T_7927; // @[MemPrimitives.scala 110:228:@51159.4]
  wire  _T_7933; // @[MemPrimitives.scala 110:228:@51163.4]
  wire  _T_7939; // @[MemPrimitives.scala 110:228:@51167.4]
  wire  _T_7945; // @[MemPrimitives.scala 110:228:@51171.4]
  wire  _T_7951; // @[MemPrimitives.scala 110:228:@51175.4]
  wire  _T_7957; // @[MemPrimitives.scala 110:228:@51179.4]
  wire  _T_7963; // @[MemPrimitives.scala 110:228:@51183.4]
  wire  _T_7969; // @[MemPrimitives.scala 110:228:@51187.4]
  wire  _T_7975; // @[MemPrimitives.scala 110:228:@51191.4]
  wire  _T_7981; // @[MemPrimitives.scala 110:228:@51195.4]
  wire  _T_7987; // @[MemPrimitives.scala 110:228:@51199.4]
  wire  _T_7989; // @[MemPrimitives.scala 123:41:@51219.4]
  wire  _T_7990; // @[MemPrimitives.scala 123:41:@51220.4]
  wire  _T_7991; // @[MemPrimitives.scala 123:41:@51221.4]
  wire  _T_7992; // @[MemPrimitives.scala 123:41:@51222.4]
  wire  _T_7993; // @[MemPrimitives.scala 123:41:@51223.4]
  wire  _T_7994; // @[MemPrimitives.scala 123:41:@51224.4]
  wire  _T_7995; // @[MemPrimitives.scala 123:41:@51225.4]
  wire  _T_7996; // @[MemPrimitives.scala 123:41:@51226.4]
  wire  _T_7997; // @[MemPrimitives.scala 123:41:@51227.4]
  wire  _T_7998; // @[MemPrimitives.scala 123:41:@51228.4]
  wire  _T_7999; // @[MemPrimitives.scala 123:41:@51229.4]
  wire  _T_8000; // @[MemPrimitives.scala 123:41:@51230.4]
  wire  _T_8001; // @[MemPrimitives.scala 123:41:@51231.4]
  wire  _T_8002; // @[MemPrimitives.scala 123:41:@51232.4]
  wire  _T_8003; // @[MemPrimitives.scala 123:41:@51233.4]
  wire [9:0] _T_8005; // @[Cat.scala 30:58:@51235.4]
  wire [9:0] _T_8007; // @[Cat.scala 30:58:@51237.4]
  wire [9:0] _T_8009; // @[Cat.scala 30:58:@51239.4]
  wire [9:0] _T_8011; // @[Cat.scala 30:58:@51241.4]
  wire [9:0] _T_8013; // @[Cat.scala 30:58:@51243.4]
  wire [9:0] _T_8015; // @[Cat.scala 30:58:@51245.4]
  wire [9:0] _T_8017; // @[Cat.scala 30:58:@51247.4]
  wire [9:0] _T_8019; // @[Cat.scala 30:58:@51249.4]
  wire [9:0] _T_8021; // @[Cat.scala 30:58:@51251.4]
  wire [9:0] _T_8023; // @[Cat.scala 30:58:@51253.4]
  wire [9:0] _T_8025; // @[Cat.scala 30:58:@51255.4]
  wire [9:0] _T_8027; // @[Cat.scala 30:58:@51257.4]
  wire [9:0] _T_8029; // @[Cat.scala 30:58:@51259.4]
  wire [9:0] _T_8031; // @[Cat.scala 30:58:@51261.4]
  wire [9:0] _T_8033; // @[Cat.scala 30:58:@51263.4]
  wire [9:0] _T_8034; // @[Mux.scala 31:69:@51264.4]
  wire [9:0] _T_8035; // @[Mux.scala 31:69:@51265.4]
  wire [9:0] _T_8036; // @[Mux.scala 31:69:@51266.4]
  wire [9:0] _T_8037; // @[Mux.scala 31:69:@51267.4]
  wire [9:0] _T_8038; // @[Mux.scala 31:69:@51268.4]
  wire [9:0] _T_8039; // @[Mux.scala 31:69:@51269.4]
  wire [9:0] _T_8040; // @[Mux.scala 31:69:@51270.4]
  wire [9:0] _T_8041; // @[Mux.scala 31:69:@51271.4]
  wire [9:0] _T_8042; // @[Mux.scala 31:69:@51272.4]
  wire [9:0] _T_8043; // @[Mux.scala 31:69:@51273.4]
  wire [9:0] _T_8044; // @[Mux.scala 31:69:@51274.4]
  wire [9:0] _T_8045; // @[Mux.scala 31:69:@51275.4]
  wire [9:0] _T_8046; // @[Mux.scala 31:69:@51276.4]
  wire [9:0] _T_8047; // @[Mux.scala 31:69:@51277.4]
  wire  _T_8055; // @[MemPrimitives.scala 110:228:@51286.4]
  wire  _T_8061; // @[MemPrimitives.scala 110:228:@51290.4]
  wire  _T_8067; // @[MemPrimitives.scala 110:228:@51294.4]
  wire  _T_8073; // @[MemPrimitives.scala 110:228:@51298.4]
  wire  _T_8079; // @[MemPrimitives.scala 110:228:@51302.4]
  wire  _T_8085; // @[MemPrimitives.scala 110:228:@51306.4]
  wire  _T_8091; // @[MemPrimitives.scala 110:228:@51310.4]
  wire  _T_8097; // @[MemPrimitives.scala 110:228:@51314.4]
  wire  _T_8103; // @[MemPrimitives.scala 110:228:@51318.4]
  wire  _T_8109; // @[MemPrimitives.scala 110:228:@51322.4]
  wire  _T_8115; // @[MemPrimitives.scala 110:228:@51326.4]
  wire  _T_8121; // @[MemPrimitives.scala 110:228:@51330.4]
  wire  _T_8127; // @[MemPrimitives.scala 110:228:@51334.4]
  wire  _T_8133; // @[MemPrimitives.scala 110:228:@51338.4]
  wire  _T_8139; // @[MemPrimitives.scala 110:228:@51342.4]
  wire  _T_8141; // @[MemPrimitives.scala 123:41:@51362.4]
  wire  _T_8142; // @[MemPrimitives.scala 123:41:@51363.4]
  wire  _T_8143; // @[MemPrimitives.scala 123:41:@51364.4]
  wire  _T_8144; // @[MemPrimitives.scala 123:41:@51365.4]
  wire  _T_8145; // @[MemPrimitives.scala 123:41:@51366.4]
  wire  _T_8146; // @[MemPrimitives.scala 123:41:@51367.4]
  wire  _T_8147; // @[MemPrimitives.scala 123:41:@51368.4]
  wire  _T_8148; // @[MemPrimitives.scala 123:41:@51369.4]
  wire  _T_8149; // @[MemPrimitives.scala 123:41:@51370.4]
  wire  _T_8150; // @[MemPrimitives.scala 123:41:@51371.4]
  wire  _T_8151; // @[MemPrimitives.scala 123:41:@51372.4]
  wire  _T_8152; // @[MemPrimitives.scala 123:41:@51373.4]
  wire  _T_8153; // @[MemPrimitives.scala 123:41:@51374.4]
  wire  _T_8154; // @[MemPrimitives.scala 123:41:@51375.4]
  wire  _T_8155; // @[MemPrimitives.scala 123:41:@51376.4]
  wire [9:0] _T_8157; // @[Cat.scala 30:58:@51378.4]
  wire [9:0] _T_8159; // @[Cat.scala 30:58:@51380.4]
  wire [9:0] _T_8161; // @[Cat.scala 30:58:@51382.4]
  wire [9:0] _T_8163; // @[Cat.scala 30:58:@51384.4]
  wire [9:0] _T_8165; // @[Cat.scala 30:58:@51386.4]
  wire [9:0] _T_8167; // @[Cat.scala 30:58:@51388.4]
  wire [9:0] _T_8169; // @[Cat.scala 30:58:@51390.4]
  wire [9:0] _T_8171; // @[Cat.scala 30:58:@51392.4]
  wire [9:0] _T_8173; // @[Cat.scala 30:58:@51394.4]
  wire [9:0] _T_8175; // @[Cat.scala 30:58:@51396.4]
  wire [9:0] _T_8177; // @[Cat.scala 30:58:@51398.4]
  wire [9:0] _T_8179; // @[Cat.scala 30:58:@51400.4]
  wire [9:0] _T_8181; // @[Cat.scala 30:58:@51402.4]
  wire [9:0] _T_8183; // @[Cat.scala 30:58:@51404.4]
  wire [9:0] _T_8185; // @[Cat.scala 30:58:@51406.4]
  wire [9:0] _T_8186; // @[Mux.scala 31:69:@51407.4]
  wire [9:0] _T_8187; // @[Mux.scala 31:69:@51408.4]
  wire [9:0] _T_8188; // @[Mux.scala 31:69:@51409.4]
  wire [9:0] _T_8189; // @[Mux.scala 31:69:@51410.4]
  wire [9:0] _T_8190; // @[Mux.scala 31:69:@51411.4]
  wire [9:0] _T_8191; // @[Mux.scala 31:69:@51412.4]
  wire [9:0] _T_8192; // @[Mux.scala 31:69:@51413.4]
  wire [9:0] _T_8193; // @[Mux.scala 31:69:@51414.4]
  wire [9:0] _T_8194; // @[Mux.scala 31:69:@51415.4]
  wire [9:0] _T_8195; // @[Mux.scala 31:69:@51416.4]
  wire [9:0] _T_8196; // @[Mux.scala 31:69:@51417.4]
  wire [9:0] _T_8197; // @[Mux.scala 31:69:@51418.4]
  wire [9:0] _T_8198; // @[Mux.scala 31:69:@51419.4]
  wire [9:0] _T_8199; // @[Mux.scala 31:69:@51420.4]
  wire  _T_8207; // @[MemPrimitives.scala 110:228:@51429.4]
  wire  _T_8213; // @[MemPrimitives.scala 110:228:@51433.4]
  wire  _T_8219; // @[MemPrimitives.scala 110:228:@51437.4]
  wire  _T_8225; // @[MemPrimitives.scala 110:228:@51441.4]
  wire  _T_8231; // @[MemPrimitives.scala 110:228:@51445.4]
  wire  _T_8237; // @[MemPrimitives.scala 110:228:@51449.4]
  wire  _T_8243; // @[MemPrimitives.scala 110:228:@51453.4]
  wire  _T_8249; // @[MemPrimitives.scala 110:228:@51457.4]
  wire  _T_8255; // @[MemPrimitives.scala 110:228:@51461.4]
  wire  _T_8261; // @[MemPrimitives.scala 110:228:@51465.4]
  wire  _T_8267; // @[MemPrimitives.scala 110:228:@51469.4]
  wire  _T_8273; // @[MemPrimitives.scala 110:228:@51473.4]
  wire  _T_8279; // @[MemPrimitives.scala 110:228:@51477.4]
  wire  _T_8285; // @[MemPrimitives.scala 110:228:@51481.4]
  wire  _T_8291; // @[MemPrimitives.scala 110:228:@51485.4]
  wire  _T_8293; // @[MemPrimitives.scala 123:41:@51505.4]
  wire  _T_8294; // @[MemPrimitives.scala 123:41:@51506.4]
  wire  _T_8295; // @[MemPrimitives.scala 123:41:@51507.4]
  wire  _T_8296; // @[MemPrimitives.scala 123:41:@51508.4]
  wire  _T_8297; // @[MemPrimitives.scala 123:41:@51509.4]
  wire  _T_8298; // @[MemPrimitives.scala 123:41:@51510.4]
  wire  _T_8299; // @[MemPrimitives.scala 123:41:@51511.4]
  wire  _T_8300; // @[MemPrimitives.scala 123:41:@51512.4]
  wire  _T_8301; // @[MemPrimitives.scala 123:41:@51513.4]
  wire  _T_8302; // @[MemPrimitives.scala 123:41:@51514.4]
  wire  _T_8303; // @[MemPrimitives.scala 123:41:@51515.4]
  wire  _T_8304; // @[MemPrimitives.scala 123:41:@51516.4]
  wire  _T_8305; // @[MemPrimitives.scala 123:41:@51517.4]
  wire  _T_8306; // @[MemPrimitives.scala 123:41:@51518.4]
  wire  _T_8307; // @[MemPrimitives.scala 123:41:@51519.4]
  wire [9:0] _T_8309; // @[Cat.scala 30:58:@51521.4]
  wire [9:0] _T_8311; // @[Cat.scala 30:58:@51523.4]
  wire [9:0] _T_8313; // @[Cat.scala 30:58:@51525.4]
  wire [9:0] _T_8315; // @[Cat.scala 30:58:@51527.4]
  wire [9:0] _T_8317; // @[Cat.scala 30:58:@51529.4]
  wire [9:0] _T_8319; // @[Cat.scala 30:58:@51531.4]
  wire [9:0] _T_8321; // @[Cat.scala 30:58:@51533.4]
  wire [9:0] _T_8323; // @[Cat.scala 30:58:@51535.4]
  wire [9:0] _T_8325; // @[Cat.scala 30:58:@51537.4]
  wire [9:0] _T_8327; // @[Cat.scala 30:58:@51539.4]
  wire [9:0] _T_8329; // @[Cat.scala 30:58:@51541.4]
  wire [9:0] _T_8331; // @[Cat.scala 30:58:@51543.4]
  wire [9:0] _T_8333; // @[Cat.scala 30:58:@51545.4]
  wire [9:0] _T_8335; // @[Cat.scala 30:58:@51547.4]
  wire [9:0] _T_8337; // @[Cat.scala 30:58:@51549.4]
  wire [9:0] _T_8338; // @[Mux.scala 31:69:@51550.4]
  wire [9:0] _T_8339; // @[Mux.scala 31:69:@51551.4]
  wire [9:0] _T_8340; // @[Mux.scala 31:69:@51552.4]
  wire [9:0] _T_8341; // @[Mux.scala 31:69:@51553.4]
  wire [9:0] _T_8342; // @[Mux.scala 31:69:@51554.4]
  wire [9:0] _T_8343; // @[Mux.scala 31:69:@51555.4]
  wire [9:0] _T_8344; // @[Mux.scala 31:69:@51556.4]
  wire [9:0] _T_8345; // @[Mux.scala 31:69:@51557.4]
  wire [9:0] _T_8346; // @[Mux.scala 31:69:@51558.4]
  wire [9:0] _T_8347; // @[Mux.scala 31:69:@51559.4]
  wire [9:0] _T_8348; // @[Mux.scala 31:69:@51560.4]
  wire [9:0] _T_8349; // @[Mux.scala 31:69:@51561.4]
  wire [9:0] _T_8350; // @[Mux.scala 31:69:@51562.4]
  wire [9:0] _T_8351; // @[Mux.scala 31:69:@51563.4]
  wire  _T_8359; // @[MemPrimitives.scala 110:228:@51572.4]
  wire  _T_8365; // @[MemPrimitives.scala 110:228:@51576.4]
  wire  _T_8371; // @[MemPrimitives.scala 110:228:@51580.4]
  wire  _T_8377; // @[MemPrimitives.scala 110:228:@51584.4]
  wire  _T_8383; // @[MemPrimitives.scala 110:228:@51588.4]
  wire  _T_8389; // @[MemPrimitives.scala 110:228:@51592.4]
  wire  _T_8395; // @[MemPrimitives.scala 110:228:@51596.4]
  wire  _T_8401; // @[MemPrimitives.scala 110:228:@51600.4]
  wire  _T_8407; // @[MemPrimitives.scala 110:228:@51604.4]
  wire  _T_8413; // @[MemPrimitives.scala 110:228:@51608.4]
  wire  _T_8419; // @[MemPrimitives.scala 110:228:@51612.4]
  wire  _T_8425; // @[MemPrimitives.scala 110:228:@51616.4]
  wire  _T_8431; // @[MemPrimitives.scala 110:228:@51620.4]
  wire  _T_8437; // @[MemPrimitives.scala 110:228:@51624.4]
  wire  _T_8443; // @[MemPrimitives.scala 110:228:@51628.4]
  wire  _T_8445; // @[MemPrimitives.scala 123:41:@51648.4]
  wire  _T_8446; // @[MemPrimitives.scala 123:41:@51649.4]
  wire  _T_8447; // @[MemPrimitives.scala 123:41:@51650.4]
  wire  _T_8448; // @[MemPrimitives.scala 123:41:@51651.4]
  wire  _T_8449; // @[MemPrimitives.scala 123:41:@51652.4]
  wire  _T_8450; // @[MemPrimitives.scala 123:41:@51653.4]
  wire  _T_8451; // @[MemPrimitives.scala 123:41:@51654.4]
  wire  _T_8452; // @[MemPrimitives.scala 123:41:@51655.4]
  wire  _T_8453; // @[MemPrimitives.scala 123:41:@51656.4]
  wire  _T_8454; // @[MemPrimitives.scala 123:41:@51657.4]
  wire  _T_8455; // @[MemPrimitives.scala 123:41:@51658.4]
  wire  _T_8456; // @[MemPrimitives.scala 123:41:@51659.4]
  wire  _T_8457; // @[MemPrimitives.scala 123:41:@51660.4]
  wire  _T_8458; // @[MemPrimitives.scala 123:41:@51661.4]
  wire  _T_8459; // @[MemPrimitives.scala 123:41:@51662.4]
  wire [9:0] _T_8461; // @[Cat.scala 30:58:@51664.4]
  wire [9:0] _T_8463; // @[Cat.scala 30:58:@51666.4]
  wire [9:0] _T_8465; // @[Cat.scala 30:58:@51668.4]
  wire [9:0] _T_8467; // @[Cat.scala 30:58:@51670.4]
  wire [9:0] _T_8469; // @[Cat.scala 30:58:@51672.4]
  wire [9:0] _T_8471; // @[Cat.scala 30:58:@51674.4]
  wire [9:0] _T_8473; // @[Cat.scala 30:58:@51676.4]
  wire [9:0] _T_8475; // @[Cat.scala 30:58:@51678.4]
  wire [9:0] _T_8477; // @[Cat.scala 30:58:@51680.4]
  wire [9:0] _T_8479; // @[Cat.scala 30:58:@51682.4]
  wire [9:0] _T_8481; // @[Cat.scala 30:58:@51684.4]
  wire [9:0] _T_8483; // @[Cat.scala 30:58:@51686.4]
  wire [9:0] _T_8485; // @[Cat.scala 30:58:@51688.4]
  wire [9:0] _T_8487; // @[Cat.scala 30:58:@51690.4]
  wire [9:0] _T_8489; // @[Cat.scala 30:58:@51692.4]
  wire [9:0] _T_8490; // @[Mux.scala 31:69:@51693.4]
  wire [9:0] _T_8491; // @[Mux.scala 31:69:@51694.4]
  wire [9:0] _T_8492; // @[Mux.scala 31:69:@51695.4]
  wire [9:0] _T_8493; // @[Mux.scala 31:69:@51696.4]
  wire [9:0] _T_8494; // @[Mux.scala 31:69:@51697.4]
  wire [9:0] _T_8495; // @[Mux.scala 31:69:@51698.4]
  wire [9:0] _T_8496; // @[Mux.scala 31:69:@51699.4]
  wire [9:0] _T_8497; // @[Mux.scala 31:69:@51700.4]
  wire [9:0] _T_8498; // @[Mux.scala 31:69:@51701.4]
  wire [9:0] _T_8499; // @[Mux.scala 31:69:@51702.4]
  wire [9:0] _T_8500; // @[Mux.scala 31:69:@51703.4]
  wire [9:0] _T_8501; // @[Mux.scala 31:69:@51704.4]
  wire [9:0] _T_8502; // @[Mux.scala 31:69:@51705.4]
  wire [9:0] _T_8503; // @[Mux.scala 31:69:@51706.4]
  wire  _T_8511; // @[MemPrimitives.scala 110:228:@51715.4]
  wire  _T_8517; // @[MemPrimitives.scala 110:228:@51719.4]
  wire  _T_8523; // @[MemPrimitives.scala 110:228:@51723.4]
  wire  _T_8529; // @[MemPrimitives.scala 110:228:@51727.4]
  wire  _T_8535; // @[MemPrimitives.scala 110:228:@51731.4]
  wire  _T_8541; // @[MemPrimitives.scala 110:228:@51735.4]
  wire  _T_8547; // @[MemPrimitives.scala 110:228:@51739.4]
  wire  _T_8553; // @[MemPrimitives.scala 110:228:@51743.4]
  wire  _T_8559; // @[MemPrimitives.scala 110:228:@51747.4]
  wire  _T_8565; // @[MemPrimitives.scala 110:228:@51751.4]
  wire  _T_8571; // @[MemPrimitives.scala 110:228:@51755.4]
  wire  _T_8577; // @[MemPrimitives.scala 110:228:@51759.4]
  wire  _T_8583; // @[MemPrimitives.scala 110:228:@51763.4]
  wire  _T_8589; // @[MemPrimitives.scala 110:228:@51767.4]
  wire  _T_8595; // @[MemPrimitives.scala 110:228:@51771.4]
  wire  _T_8597; // @[MemPrimitives.scala 123:41:@51791.4]
  wire  _T_8598; // @[MemPrimitives.scala 123:41:@51792.4]
  wire  _T_8599; // @[MemPrimitives.scala 123:41:@51793.4]
  wire  _T_8600; // @[MemPrimitives.scala 123:41:@51794.4]
  wire  _T_8601; // @[MemPrimitives.scala 123:41:@51795.4]
  wire  _T_8602; // @[MemPrimitives.scala 123:41:@51796.4]
  wire  _T_8603; // @[MemPrimitives.scala 123:41:@51797.4]
  wire  _T_8604; // @[MemPrimitives.scala 123:41:@51798.4]
  wire  _T_8605; // @[MemPrimitives.scala 123:41:@51799.4]
  wire  _T_8606; // @[MemPrimitives.scala 123:41:@51800.4]
  wire  _T_8607; // @[MemPrimitives.scala 123:41:@51801.4]
  wire  _T_8608; // @[MemPrimitives.scala 123:41:@51802.4]
  wire  _T_8609; // @[MemPrimitives.scala 123:41:@51803.4]
  wire  _T_8610; // @[MemPrimitives.scala 123:41:@51804.4]
  wire  _T_8611; // @[MemPrimitives.scala 123:41:@51805.4]
  wire [9:0] _T_8613; // @[Cat.scala 30:58:@51807.4]
  wire [9:0] _T_8615; // @[Cat.scala 30:58:@51809.4]
  wire [9:0] _T_8617; // @[Cat.scala 30:58:@51811.4]
  wire [9:0] _T_8619; // @[Cat.scala 30:58:@51813.4]
  wire [9:0] _T_8621; // @[Cat.scala 30:58:@51815.4]
  wire [9:0] _T_8623; // @[Cat.scala 30:58:@51817.4]
  wire [9:0] _T_8625; // @[Cat.scala 30:58:@51819.4]
  wire [9:0] _T_8627; // @[Cat.scala 30:58:@51821.4]
  wire [9:0] _T_8629; // @[Cat.scala 30:58:@51823.4]
  wire [9:0] _T_8631; // @[Cat.scala 30:58:@51825.4]
  wire [9:0] _T_8633; // @[Cat.scala 30:58:@51827.4]
  wire [9:0] _T_8635; // @[Cat.scala 30:58:@51829.4]
  wire [9:0] _T_8637; // @[Cat.scala 30:58:@51831.4]
  wire [9:0] _T_8639; // @[Cat.scala 30:58:@51833.4]
  wire [9:0] _T_8641; // @[Cat.scala 30:58:@51835.4]
  wire [9:0] _T_8642; // @[Mux.scala 31:69:@51836.4]
  wire [9:0] _T_8643; // @[Mux.scala 31:69:@51837.4]
  wire [9:0] _T_8644; // @[Mux.scala 31:69:@51838.4]
  wire [9:0] _T_8645; // @[Mux.scala 31:69:@51839.4]
  wire [9:0] _T_8646; // @[Mux.scala 31:69:@51840.4]
  wire [9:0] _T_8647; // @[Mux.scala 31:69:@51841.4]
  wire [9:0] _T_8648; // @[Mux.scala 31:69:@51842.4]
  wire [9:0] _T_8649; // @[Mux.scala 31:69:@51843.4]
  wire [9:0] _T_8650; // @[Mux.scala 31:69:@51844.4]
  wire [9:0] _T_8651; // @[Mux.scala 31:69:@51845.4]
  wire [9:0] _T_8652; // @[Mux.scala 31:69:@51846.4]
  wire [9:0] _T_8653; // @[Mux.scala 31:69:@51847.4]
  wire [9:0] _T_8654; // @[Mux.scala 31:69:@51848.4]
  wire [9:0] _T_8655; // @[Mux.scala 31:69:@51849.4]
  wire  _T_8663; // @[MemPrimitives.scala 110:228:@51858.4]
  wire  _T_8669; // @[MemPrimitives.scala 110:228:@51862.4]
  wire  _T_8675; // @[MemPrimitives.scala 110:228:@51866.4]
  wire  _T_8681; // @[MemPrimitives.scala 110:228:@51870.4]
  wire  _T_8687; // @[MemPrimitives.scala 110:228:@51874.4]
  wire  _T_8693; // @[MemPrimitives.scala 110:228:@51878.4]
  wire  _T_8699; // @[MemPrimitives.scala 110:228:@51882.4]
  wire  _T_8705; // @[MemPrimitives.scala 110:228:@51886.4]
  wire  _T_8711; // @[MemPrimitives.scala 110:228:@51890.4]
  wire  _T_8717; // @[MemPrimitives.scala 110:228:@51894.4]
  wire  _T_8723; // @[MemPrimitives.scala 110:228:@51898.4]
  wire  _T_8729; // @[MemPrimitives.scala 110:228:@51902.4]
  wire  _T_8735; // @[MemPrimitives.scala 110:228:@51906.4]
  wire  _T_8741; // @[MemPrimitives.scala 110:228:@51910.4]
  wire  _T_8747; // @[MemPrimitives.scala 110:228:@51914.4]
  wire  _T_8749; // @[MemPrimitives.scala 123:41:@51934.4]
  wire  _T_8750; // @[MemPrimitives.scala 123:41:@51935.4]
  wire  _T_8751; // @[MemPrimitives.scala 123:41:@51936.4]
  wire  _T_8752; // @[MemPrimitives.scala 123:41:@51937.4]
  wire  _T_8753; // @[MemPrimitives.scala 123:41:@51938.4]
  wire  _T_8754; // @[MemPrimitives.scala 123:41:@51939.4]
  wire  _T_8755; // @[MemPrimitives.scala 123:41:@51940.4]
  wire  _T_8756; // @[MemPrimitives.scala 123:41:@51941.4]
  wire  _T_8757; // @[MemPrimitives.scala 123:41:@51942.4]
  wire  _T_8758; // @[MemPrimitives.scala 123:41:@51943.4]
  wire  _T_8759; // @[MemPrimitives.scala 123:41:@51944.4]
  wire  _T_8760; // @[MemPrimitives.scala 123:41:@51945.4]
  wire  _T_8761; // @[MemPrimitives.scala 123:41:@51946.4]
  wire  _T_8762; // @[MemPrimitives.scala 123:41:@51947.4]
  wire  _T_8763; // @[MemPrimitives.scala 123:41:@51948.4]
  wire [9:0] _T_8765; // @[Cat.scala 30:58:@51950.4]
  wire [9:0] _T_8767; // @[Cat.scala 30:58:@51952.4]
  wire [9:0] _T_8769; // @[Cat.scala 30:58:@51954.4]
  wire [9:0] _T_8771; // @[Cat.scala 30:58:@51956.4]
  wire [9:0] _T_8773; // @[Cat.scala 30:58:@51958.4]
  wire [9:0] _T_8775; // @[Cat.scala 30:58:@51960.4]
  wire [9:0] _T_8777; // @[Cat.scala 30:58:@51962.4]
  wire [9:0] _T_8779; // @[Cat.scala 30:58:@51964.4]
  wire [9:0] _T_8781; // @[Cat.scala 30:58:@51966.4]
  wire [9:0] _T_8783; // @[Cat.scala 30:58:@51968.4]
  wire [9:0] _T_8785; // @[Cat.scala 30:58:@51970.4]
  wire [9:0] _T_8787; // @[Cat.scala 30:58:@51972.4]
  wire [9:0] _T_8789; // @[Cat.scala 30:58:@51974.4]
  wire [9:0] _T_8791; // @[Cat.scala 30:58:@51976.4]
  wire [9:0] _T_8793; // @[Cat.scala 30:58:@51978.4]
  wire [9:0] _T_8794; // @[Mux.scala 31:69:@51979.4]
  wire [9:0] _T_8795; // @[Mux.scala 31:69:@51980.4]
  wire [9:0] _T_8796; // @[Mux.scala 31:69:@51981.4]
  wire [9:0] _T_8797; // @[Mux.scala 31:69:@51982.4]
  wire [9:0] _T_8798; // @[Mux.scala 31:69:@51983.4]
  wire [9:0] _T_8799; // @[Mux.scala 31:69:@51984.4]
  wire [9:0] _T_8800; // @[Mux.scala 31:69:@51985.4]
  wire [9:0] _T_8801; // @[Mux.scala 31:69:@51986.4]
  wire [9:0] _T_8802; // @[Mux.scala 31:69:@51987.4]
  wire [9:0] _T_8803; // @[Mux.scala 31:69:@51988.4]
  wire [9:0] _T_8804; // @[Mux.scala 31:69:@51989.4]
  wire [9:0] _T_8805; // @[Mux.scala 31:69:@51990.4]
  wire [9:0] _T_8806; // @[Mux.scala 31:69:@51991.4]
  wire [9:0] _T_8807; // @[Mux.scala 31:69:@51992.4]
  wire  _T_8967; // @[package.scala 96:25:@52209.4 package.scala 96:25:@52210.4]
  wire [7:0] _T_8971; // @[Mux.scala 31:69:@52219.4]
  wire  _T_8964; // @[package.scala 96:25:@52201.4 package.scala 96:25:@52202.4]
  wire [7:0] _T_8972; // @[Mux.scala 31:69:@52220.4]
  wire  _T_8961; // @[package.scala 96:25:@52193.4 package.scala 96:25:@52194.4]
  wire [7:0] _T_8973; // @[Mux.scala 31:69:@52221.4]
  wire  _T_8958; // @[package.scala 96:25:@52185.4 package.scala 96:25:@52186.4]
  wire [7:0] _T_8974; // @[Mux.scala 31:69:@52222.4]
  wire  _T_8955; // @[package.scala 96:25:@52177.4 package.scala 96:25:@52178.4]
  wire [7:0] _T_8975; // @[Mux.scala 31:69:@52223.4]
  wire  _T_8952; // @[package.scala 96:25:@52169.4 package.scala 96:25:@52170.4]
  wire [7:0] _T_8976; // @[Mux.scala 31:69:@52224.4]
  wire  _T_8949; // @[package.scala 96:25:@52161.4 package.scala 96:25:@52162.4]
  wire [7:0] _T_8977; // @[Mux.scala 31:69:@52225.4]
  wire  _T_8946; // @[package.scala 96:25:@52153.4 package.scala 96:25:@52154.4]
  wire [7:0] _T_8978; // @[Mux.scala 31:69:@52226.4]
  wire  _T_8943; // @[package.scala 96:25:@52145.4 package.scala 96:25:@52146.4]
  wire [7:0] _T_8979; // @[Mux.scala 31:69:@52227.4]
  wire  _T_8940; // @[package.scala 96:25:@52137.4 package.scala 96:25:@52138.4]
  wire [7:0] _T_8980; // @[Mux.scala 31:69:@52228.4]
  wire  _T_8937; // @[package.scala 96:25:@52129.4 package.scala 96:25:@52130.4]
  wire [7:0] _T_8981; // @[Mux.scala 31:69:@52229.4]
  wire  _T_8934; // @[package.scala 96:25:@52121.4 package.scala 96:25:@52122.4]
  wire [7:0] _T_8982; // @[Mux.scala 31:69:@52230.4]
  wire  _T_8931; // @[package.scala 96:25:@52113.4 package.scala 96:25:@52114.4]
  wire [7:0] _T_8983; // @[Mux.scala 31:69:@52231.4]
  wire  _T_8928; // @[package.scala 96:25:@52105.4 package.scala 96:25:@52106.4]
  wire [7:0] _T_8984; // @[Mux.scala 31:69:@52232.4]
  wire  _T_8925; // @[package.scala 96:25:@52097.4 package.scala 96:25:@52098.4]
  wire [7:0] _T_8985; // @[Mux.scala 31:69:@52233.4]
  wire  _T_8922; // @[package.scala 96:25:@52089.4 package.scala 96:25:@52090.4]
  wire [7:0] _T_8986; // @[Mux.scala 31:69:@52234.4]
  wire  _T_8919; // @[package.scala 96:25:@52081.4 package.scala 96:25:@52082.4]
  wire [7:0] _T_8987; // @[Mux.scala 31:69:@52235.4]
  wire  _T_8916; // @[package.scala 96:25:@52073.4 package.scala 96:25:@52074.4]
  wire [7:0] _T_8988; // @[Mux.scala 31:69:@52236.4]
  wire  _T_8913; // @[package.scala 96:25:@52065.4 package.scala 96:25:@52066.4]
  wire  _T_9146; // @[package.scala 96:25:@52449.4 package.scala 96:25:@52450.4]
  wire [7:0] _T_9150; // @[Mux.scala 31:69:@52459.4]
  wire  _T_9143; // @[package.scala 96:25:@52441.4 package.scala 96:25:@52442.4]
  wire [7:0] _T_9151; // @[Mux.scala 31:69:@52460.4]
  wire  _T_9140; // @[package.scala 96:25:@52433.4 package.scala 96:25:@52434.4]
  wire [7:0] _T_9152; // @[Mux.scala 31:69:@52461.4]
  wire  _T_9137; // @[package.scala 96:25:@52425.4 package.scala 96:25:@52426.4]
  wire [7:0] _T_9153; // @[Mux.scala 31:69:@52462.4]
  wire  _T_9134; // @[package.scala 96:25:@52417.4 package.scala 96:25:@52418.4]
  wire [7:0] _T_9154; // @[Mux.scala 31:69:@52463.4]
  wire  _T_9131; // @[package.scala 96:25:@52409.4 package.scala 96:25:@52410.4]
  wire [7:0] _T_9155; // @[Mux.scala 31:69:@52464.4]
  wire  _T_9128; // @[package.scala 96:25:@52401.4 package.scala 96:25:@52402.4]
  wire [7:0] _T_9156; // @[Mux.scala 31:69:@52465.4]
  wire  _T_9125; // @[package.scala 96:25:@52393.4 package.scala 96:25:@52394.4]
  wire [7:0] _T_9157; // @[Mux.scala 31:69:@52466.4]
  wire  _T_9122; // @[package.scala 96:25:@52385.4 package.scala 96:25:@52386.4]
  wire [7:0] _T_9158; // @[Mux.scala 31:69:@52467.4]
  wire  _T_9119; // @[package.scala 96:25:@52377.4 package.scala 96:25:@52378.4]
  wire [7:0] _T_9159; // @[Mux.scala 31:69:@52468.4]
  wire  _T_9116; // @[package.scala 96:25:@52369.4 package.scala 96:25:@52370.4]
  wire [7:0] _T_9160; // @[Mux.scala 31:69:@52469.4]
  wire  _T_9113; // @[package.scala 96:25:@52361.4 package.scala 96:25:@52362.4]
  wire [7:0] _T_9161; // @[Mux.scala 31:69:@52470.4]
  wire  _T_9110; // @[package.scala 96:25:@52353.4 package.scala 96:25:@52354.4]
  wire [7:0] _T_9162; // @[Mux.scala 31:69:@52471.4]
  wire  _T_9107; // @[package.scala 96:25:@52345.4 package.scala 96:25:@52346.4]
  wire [7:0] _T_9163; // @[Mux.scala 31:69:@52472.4]
  wire  _T_9104; // @[package.scala 96:25:@52337.4 package.scala 96:25:@52338.4]
  wire [7:0] _T_9164; // @[Mux.scala 31:69:@52473.4]
  wire  _T_9101; // @[package.scala 96:25:@52329.4 package.scala 96:25:@52330.4]
  wire [7:0] _T_9165; // @[Mux.scala 31:69:@52474.4]
  wire  _T_9098; // @[package.scala 96:25:@52321.4 package.scala 96:25:@52322.4]
  wire [7:0] _T_9166; // @[Mux.scala 31:69:@52475.4]
  wire  _T_9095; // @[package.scala 96:25:@52313.4 package.scala 96:25:@52314.4]
  wire [7:0] _T_9167; // @[Mux.scala 31:69:@52476.4]
  wire  _T_9092; // @[package.scala 96:25:@52305.4 package.scala 96:25:@52306.4]
  wire  _T_9325; // @[package.scala 96:25:@52689.4 package.scala 96:25:@52690.4]
  wire [7:0] _T_9329; // @[Mux.scala 31:69:@52699.4]
  wire  _T_9322; // @[package.scala 96:25:@52681.4 package.scala 96:25:@52682.4]
  wire [7:0] _T_9330; // @[Mux.scala 31:69:@52700.4]
  wire  _T_9319; // @[package.scala 96:25:@52673.4 package.scala 96:25:@52674.4]
  wire [7:0] _T_9331; // @[Mux.scala 31:69:@52701.4]
  wire  _T_9316; // @[package.scala 96:25:@52665.4 package.scala 96:25:@52666.4]
  wire [7:0] _T_9332; // @[Mux.scala 31:69:@52702.4]
  wire  _T_9313; // @[package.scala 96:25:@52657.4 package.scala 96:25:@52658.4]
  wire [7:0] _T_9333; // @[Mux.scala 31:69:@52703.4]
  wire  _T_9310; // @[package.scala 96:25:@52649.4 package.scala 96:25:@52650.4]
  wire [7:0] _T_9334; // @[Mux.scala 31:69:@52704.4]
  wire  _T_9307; // @[package.scala 96:25:@52641.4 package.scala 96:25:@52642.4]
  wire [7:0] _T_9335; // @[Mux.scala 31:69:@52705.4]
  wire  _T_9304; // @[package.scala 96:25:@52633.4 package.scala 96:25:@52634.4]
  wire [7:0] _T_9336; // @[Mux.scala 31:69:@52706.4]
  wire  _T_9301; // @[package.scala 96:25:@52625.4 package.scala 96:25:@52626.4]
  wire [7:0] _T_9337; // @[Mux.scala 31:69:@52707.4]
  wire  _T_9298; // @[package.scala 96:25:@52617.4 package.scala 96:25:@52618.4]
  wire [7:0] _T_9338; // @[Mux.scala 31:69:@52708.4]
  wire  _T_9295; // @[package.scala 96:25:@52609.4 package.scala 96:25:@52610.4]
  wire [7:0] _T_9339; // @[Mux.scala 31:69:@52709.4]
  wire  _T_9292; // @[package.scala 96:25:@52601.4 package.scala 96:25:@52602.4]
  wire [7:0] _T_9340; // @[Mux.scala 31:69:@52710.4]
  wire  _T_9289; // @[package.scala 96:25:@52593.4 package.scala 96:25:@52594.4]
  wire [7:0] _T_9341; // @[Mux.scala 31:69:@52711.4]
  wire  _T_9286; // @[package.scala 96:25:@52585.4 package.scala 96:25:@52586.4]
  wire [7:0] _T_9342; // @[Mux.scala 31:69:@52712.4]
  wire  _T_9283; // @[package.scala 96:25:@52577.4 package.scala 96:25:@52578.4]
  wire [7:0] _T_9343; // @[Mux.scala 31:69:@52713.4]
  wire  _T_9280; // @[package.scala 96:25:@52569.4 package.scala 96:25:@52570.4]
  wire [7:0] _T_9344; // @[Mux.scala 31:69:@52714.4]
  wire  _T_9277; // @[package.scala 96:25:@52561.4 package.scala 96:25:@52562.4]
  wire [7:0] _T_9345; // @[Mux.scala 31:69:@52715.4]
  wire  _T_9274; // @[package.scala 96:25:@52553.4 package.scala 96:25:@52554.4]
  wire [7:0] _T_9346; // @[Mux.scala 31:69:@52716.4]
  wire  _T_9271; // @[package.scala 96:25:@52545.4 package.scala 96:25:@52546.4]
  wire  _T_9504; // @[package.scala 96:25:@52929.4 package.scala 96:25:@52930.4]
  wire [7:0] _T_9508; // @[Mux.scala 31:69:@52939.4]
  wire  _T_9501; // @[package.scala 96:25:@52921.4 package.scala 96:25:@52922.4]
  wire [7:0] _T_9509; // @[Mux.scala 31:69:@52940.4]
  wire  _T_9498; // @[package.scala 96:25:@52913.4 package.scala 96:25:@52914.4]
  wire [7:0] _T_9510; // @[Mux.scala 31:69:@52941.4]
  wire  _T_9495; // @[package.scala 96:25:@52905.4 package.scala 96:25:@52906.4]
  wire [7:0] _T_9511; // @[Mux.scala 31:69:@52942.4]
  wire  _T_9492; // @[package.scala 96:25:@52897.4 package.scala 96:25:@52898.4]
  wire [7:0] _T_9512; // @[Mux.scala 31:69:@52943.4]
  wire  _T_9489; // @[package.scala 96:25:@52889.4 package.scala 96:25:@52890.4]
  wire [7:0] _T_9513; // @[Mux.scala 31:69:@52944.4]
  wire  _T_9486; // @[package.scala 96:25:@52881.4 package.scala 96:25:@52882.4]
  wire [7:0] _T_9514; // @[Mux.scala 31:69:@52945.4]
  wire  _T_9483; // @[package.scala 96:25:@52873.4 package.scala 96:25:@52874.4]
  wire [7:0] _T_9515; // @[Mux.scala 31:69:@52946.4]
  wire  _T_9480; // @[package.scala 96:25:@52865.4 package.scala 96:25:@52866.4]
  wire [7:0] _T_9516; // @[Mux.scala 31:69:@52947.4]
  wire  _T_9477; // @[package.scala 96:25:@52857.4 package.scala 96:25:@52858.4]
  wire [7:0] _T_9517; // @[Mux.scala 31:69:@52948.4]
  wire  _T_9474; // @[package.scala 96:25:@52849.4 package.scala 96:25:@52850.4]
  wire [7:0] _T_9518; // @[Mux.scala 31:69:@52949.4]
  wire  _T_9471; // @[package.scala 96:25:@52841.4 package.scala 96:25:@52842.4]
  wire [7:0] _T_9519; // @[Mux.scala 31:69:@52950.4]
  wire  _T_9468; // @[package.scala 96:25:@52833.4 package.scala 96:25:@52834.4]
  wire [7:0] _T_9520; // @[Mux.scala 31:69:@52951.4]
  wire  _T_9465; // @[package.scala 96:25:@52825.4 package.scala 96:25:@52826.4]
  wire [7:0] _T_9521; // @[Mux.scala 31:69:@52952.4]
  wire  _T_9462; // @[package.scala 96:25:@52817.4 package.scala 96:25:@52818.4]
  wire [7:0] _T_9522; // @[Mux.scala 31:69:@52953.4]
  wire  _T_9459; // @[package.scala 96:25:@52809.4 package.scala 96:25:@52810.4]
  wire [7:0] _T_9523; // @[Mux.scala 31:69:@52954.4]
  wire  _T_9456; // @[package.scala 96:25:@52801.4 package.scala 96:25:@52802.4]
  wire [7:0] _T_9524; // @[Mux.scala 31:69:@52955.4]
  wire  _T_9453; // @[package.scala 96:25:@52793.4 package.scala 96:25:@52794.4]
  wire [7:0] _T_9525; // @[Mux.scala 31:69:@52956.4]
  wire  _T_9450; // @[package.scala 96:25:@52785.4 package.scala 96:25:@52786.4]
  wire  _T_9683; // @[package.scala 96:25:@53169.4 package.scala 96:25:@53170.4]
  wire [7:0] _T_9687; // @[Mux.scala 31:69:@53179.4]
  wire  _T_9680; // @[package.scala 96:25:@53161.4 package.scala 96:25:@53162.4]
  wire [7:0] _T_9688; // @[Mux.scala 31:69:@53180.4]
  wire  _T_9677; // @[package.scala 96:25:@53153.4 package.scala 96:25:@53154.4]
  wire [7:0] _T_9689; // @[Mux.scala 31:69:@53181.4]
  wire  _T_9674; // @[package.scala 96:25:@53145.4 package.scala 96:25:@53146.4]
  wire [7:0] _T_9690; // @[Mux.scala 31:69:@53182.4]
  wire  _T_9671; // @[package.scala 96:25:@53137.4 package.scala 96:25:@53138.4]
  wire [7:0] _T_9691; // @[Mux.scala 31:69:@53183.4]
  wire  _T_9668; // @[package.scala 96:25:@53129.4 package.scala 96:25:@53130.4]
  wire [7:0] _T_9692; // @[Mux.scala 31:69:@53184.4]
  wire  _T_9665; // @[package.scala 96:25:@53121.4 package.scala 96:25:@53122.4]
  wire [7:0] _T_9693; // @[Mux.scala 31:69:@53185.4]
  wire  _T_9662; // @[package.scala 96:25:@53113.4 package.scala 96:25:@53114.4]
  wire [7:0] _T_9694; // @[Mux.scala 31:69:@53186.4]
  wire  _T_9659; // @[package.scala 96:25:@53105.4 package.scala 96:25:@53106.4]
  wire [7:0] _T_9695; // @[Mux.scala 31:69:@53187.4]
  wire  _T_9656; // @[package.scala 96:25:@53097.4 package.scala 96:25:@53098.4]
  wire [7:0] _T_9696; // @[Mux.scala 31:69:@53188.4]
  wire  _T_9653; // @[package.scala 96:25:@53089.4 package.scala 96:25:@53090.4]
  wire [7:0] _T_9697; // @[Mux.scala 31:69:@53189.4]
  wire  _T_9650; // @[package.scala 96:25:@53081.4 package.scala 96:25:@53082.4]
  wire [7:0] _T_9698; // @[Mux.scala 31:69:@53190.4]
  wire  _T_9647; // @[package.scala 96:25:@53073.4 package.scala 96:25:@53074.4]
  wire [7:0] _T_9699; // @[Mux.scala 31:69:@53191.4]
  wire  _T_9644; // @[package.scala 96:25:@53065.4 package.scala 96:25:@53066.4]
  wire [7:0] _T_9700; // @[Mux.scala 31:69:@53192.4]
  wire  _T_9641; // @[package.scala 96:25:@53057.4 package.scala 96:25:@53058.4]
  wire [7:0] _T_9701; // @[Mux.scala 31:69:@53193.4]
  wire  _T_9638; // @[package.scala 96:25:@53049.4 package.scala 96:25:@53050.4]
  wire [7:0] _T_9702; // @[Mux.scala 31:69:@53194.4]
  wire  _T_9635; // @[package.scala 96:25:@53041.4 package.scala 96:25:@53042.4]
  wire [7:0] _T_9703; // @[Mux.scala 31:69:@53195.4]
  wire  _T_9632; // @[package.scala 96:25:@53033.4 package.scala 96:25:@53034.4]
  wire [7:0] _T_9704; // @[Mux.scala 31:69:@53196.4]
  wire  _T_9629; // @[package.scala 96:25:@53025.4 package.scala 96:25:@53026.4]
  wire  _T_9862; // @[package.scala 96:25:@53409.4 package.scala 96:25:@53410.4]
  wire [7:0] _T_9866; // @[Mux.scala 31:69:@53419.4]
  wire  _T_9859; // @[package.scala 96:25:@53401.4 package.scala 96:25:@53402.4]
  wire [7:0] _T_9867; // @[Mux.scala 31:69:@53420.4]
  wire  _T_9856; // @[package.scala 96:25:@53393.4 package.scala 96:25:@53394.4]
  wire [7:0] _T_9868; // @[Mux.scala 31:69:@53421.4]
  wire  _T_9853; // @[package.scala 96:25:@53385.4 package.scala 96:25:@53386.4]
  wire [7:0] _T_9869; // @[Mux.scala 31:69:@53422.4]
  wire  _T_9850; // @[package.scala 96:25:@53377.4 package.scala 96:25:@53378.4]
  wire [7:0] _T_9870; // @[Mux.scala 31:69:@53423.4]
  wire  _T_9847; // @[package.scala 96:25:@53369.4 package.scala 96:25:@53370.4]
  wire [7:0] _T_9871; // @[Mux.scala 31:69:@53424.4]
  wire  _T_9844; // @[package.scala 96:25:@53361.4 package.scala 96:25:@53362.4]
  wire [7:0] _T_9872; // @[Mux.scala 31:69:@53425.4]
  wire  _T_9841; // @[package.scala 96:25:@53353.4 package.scala 96:25:@53354.4]
  wire [7:0] _T_9873; // @[Mux.scala 31:69:@53426.4]
  wire  _T_9838; // @[package.scala 96:25:@53345.4 package.scala 96:25:@53346.4]
  wire [7:0] _T_9874; // @[Mux.scala 31:69:@53427.4]
  wire  _T_9835; // @[package.scala 96:25:@53337.4 package.scala 96:25:@53338.4]
  wire [7:0] _T_9875; // @[Mux.scala 31:69:@53428.4]
  wire  _T_9832; // @[package.scala 96:25:@53329.4 package.scala 96:25:@53330.4]
  wire [7:0] _T_9876; // @[Mux.scala 31:69:@53429.4]
  wire  _T_9829; // @[package.scala 96:25:@53321.4 package.scala 96:25:@53322.4]
  wire [7:0] _T_9877; // @[Mux.scala 31:69:@53430.4]
  wire  _T_9826; // @[package.scala 96:25:@53313.4 package.scala 96:25:@53314.4]
  wire [7:0] _T_9878; // @[Mux.scala 31:69:@53431.4]
  wire  _T_9823; // @[package.scala 96:25:@53305.4 package.scala 96:25:@53306.4]
  wire [7:0] _T_9879; // @[Mux.scala 31:69:@53432.4]
  wire  _T_9820; // @[package.scala 96:25:@53297.4 package.scala 96:25:@53298.4]
  wire [7:0] _T_9880; // @[Mux.scala 31:69:@53433.4]
  wire  _T_9817; // @[package.scala 96:25:@53289.4 package.scala 96:25:@53290.4]
  wire [7:0] _T_9881; // @[Mux.scala 31:69:@53434.4]
  wire  _T_9814; // @[package.scala 96:25:@53281.4 package.scala 96:25:@53282.4]
  wire [7:0] _T_9882; // @[Mux.scala 31:69:@53435.4]
  wire  _T_9811; // @[package.scala 96:25:@53273.4 package.scala 96:25:@53274.4]
  wire [7:0] _T_9883; // @[Mux.scala 31:69:@53436.4]
  wire  _T_9808; // @[package.scala 96:25:@53265.4 package.scala 96:25:@53266.4]
  wire  _T_10041; // @[package.scala 96:25:@53649.4 package.scala 96:25:@53650.4]
  wire [7:0] _T_10045; // @[Mux.scala 31:69:@53659.4]
  wire  _T_10038; // @[package.scala 96:25:@53641.4 package.scala 96:25:@53642.4]
  wire [7:0] _T_10046; // @[Mux.scala 31:69:@53660.4]
  wire  _T_10035; // @[package.scala 96:25:@53633.4 package.scala 96:25:@53634.4]
  wire [7:0] _T_10047; // @[Mux.scala 31:69:@53661.4]
  wire  _T_10032; // @[package.scala 96:25:@53625.4 package.scala 96:25:@53626.4]
  wire [7:0] _T_10048; // @[Mux.scala 31:69:@53662.4]
  wire  _T_10029; // @[package.scala 96:25:@53617.4 package.scala 96:25:@53618.4]
  wire [7:0] _T_10049; // @[Mux.scala 31:69:@53663.4]
  wire  _T_10026; // @[package.scala 96:25:@53609.4 package.scala 96:25:@53610.4]
  wire [7:0] _T_10050; // @[Mux.scala 31:69:@53664.4]
  wire  _T_10023; // @[package.scala 96:25:@53601.4 package.scala 96:25:@53602.4]
  wire [7:0] _T_10051; // @[Mux.scala 31:69:@53665.4]
  wire  _T_10020; // @[package.scala 96:25:@53593.4 package.scala 96:25:@53594.4]
  wire [7:0] _T_10052; // @[Mux.scala 31:69:@53666.4]
  wire  _T_10017; // @[package.scala 96:25:@53585.4 package.scala 96:25:@53586.4]
  wire [7:0] _T_10053; // @[Mux.scala 31:69:@53667.4]
  wire  _T_10014; // @[package.scala 96:25:@53577.4 package.scala 96:25:@53578.4]
  wire [7:0] _T_10054; // @[Mux.scala 31:69:@53668.4]
  wire  _T_10011; // @[package.scala 96:25:@53569.4 package.scala 96:25:@53570.4]
  wire [7:0] _T_10055; // @[Mux.scala 31:69:@53669.4]
  wire  _T_10008; // @[package.scala 96:25:@53561.4 package.scala 96:25:@53562.4]
  wire [7:0] _T_10056; // @[Mux.scala 31:69:@53670.4]
  wire  _T_10005; // @[package.scala 96:25:@53553.4 package.scala 96:25:@53554.4]
  wire [7:0] _T_10057; // @[Mux.scala 31:69:@53671.4]
  wire  _T_10002; // @[package.scala 96:25:@53545.4 package.scala 96:25:@53546.4]
  wire [7:0] _T_10058; // @[Mux.scala 31:69:@53672.4]
  wire  _T_9999; // @[package.scala 96:25:@53537.4 package.scala 96:25:@53538.4]
  wire [7:0] _T_10059; // @[Mux.scala 31:69:@53673.4]
  wire  _T_9996; // @[package.scala 96:25:@53529.4 package.scala 96:25:@53530.4]
  wire [7:0] _T_10060; // @[Mux.scala 31:69:@53674.4]
  wire  _T_9993; // @[package.scala 96:25:@53521.4 package.scala 96:25:@53522.4]
  wire [7:0] _T_10061; // @[Mux.scala 31:69:@53675.4]
  wire  _T_9990; // @[package.scala 96:25:@53513.4 package.scala 96:25:@53514.4]
  wire [7:0] _T_10062; // @[Mux.scala 31:69:@53676.4]
  wire  _T_9987; // @[package.scala 96:25:@53505.4 package.scala 96:25:@53506.4]
  wire  _T_10220; // @[package.scala 96:25:@53889.4 package.scala 96:25:@53890.4]
  wire [7:0] _T_10224; // @[Mux.scala 31:69:@53899.4]
  wire  _T_10217; // @[package.scala 96:25:@53881.4 package.scala 96:25:@53882.4]
  wire [7:0] _T_10225; // @[Mux.scala 31:69:@53900.4]
  wire  _T_10214; // @[package.scala 96:25:@53873.4 package.scala 96:25:@53874.4]
  wire [7:0] _T_10226; // @[Mux.scala 31:69:@53901.4]
  wire  _T_10211; // @[package.scala 96:25:@53865.4 package.scala 96:25:@53866.4]
  wire [7:0] _T_10227; // @[Mux.scala 31:69:@53902.4]
  wire  _T_10208; // @[package.scala 96:25:@53857.4 package.scala 96:25:@53858.4]
  wire [7:0] _T_10228; // @[Mux.scala 31:69:@53903.4]
  wire  _T_10205; // @[package.scala 96:25:@53849.4 package.scala 96:25:@53850.4]
  wire [7:0] _T_10229; // @[Mux.scala 31:69:@53904.4]
  wire  _T_10202; // @[package.scala 96:25:@53841.4 package.scala 96:25:@53842.4]
  wire [7:0] _T_10230; // @[Mux.scala 31:69:@53905.4]
  wire  _T_10199; // @[package.scala 96:25:@53833.4 package.scala 96:25:@53834.4]
  wire [7:0] _T_10231; // @[Mux.scala 31:69:@53906.4]
  wire  _T_10196; // @[package.scala 96:25:@53825.4 package.scala 96:25:@53826.4]
  wire [7:0] _T_10232; // @[Mux.scala 31:69:@53907.4]
  wire  _T_10193; // @[package.scala 96:25:@53817.4 package.scala 96:25:@53818.4]
  wire [7:0] _T_10233; // @[Mux.scala 31:69:@53908.4]
  wire  _T_10190; // @[package.scala 96:25:@53809.4 package.scala 96:25:@53810.4]
  wire [7:0] _T_10234; // @[Mux.scala 31:69:@53909.4]
  wire  _T_10187; // @[package.scala 96:25:@53801.4 package.scala 96:25:@53802.4]
  wire [7:0] _T_10235; // @[Mux.scala 31:69:@53910.4]
  wire  _T_10184; // @[package.scala 96:25:@53793.4 package.scala 96:25:@53794.4]
  wire [7:0] _T_10236; // @[Mux.scala 31:69:@53911.4]
  wire  _T_10181; // @[package.scala 96:25:@53785.4 package.scala 96:25:@53786.4]
  wire [7:0] _T_10237; // @[Mux.scala 31:69:@53912.4]
  wire  _T_10178; // @[package.scala 96:25:@53777.4 package.scala 96:25:@53778.4]
  wire [7:0] _T_10238; // @[Mux.scala 31:69:@53913.4]
  wire  _T_10175; // @[package.scala 96:25:@53769.4 package.scala 96:25:@53770.4]
  wire [7:0] _T_10239; // @[Mux.scala 31:69:@53914.4]
  wire  _T_10172; // @[package.scala 96:25:@53761.4 package.scala 96:25:@53762.4]
  wire [7:0] _T_10240; // @[Mux.scala 31:69:@53915.4]
  wire  _T_10169; // @[package.scala 96:25:@53753.4 package.scala 96:25:@53754.4]
  wire [7:0] _T_10241; // @[Mux.scala 31:69:@53916.4]
  wire  _T_10166; // @[package.scala 96:25:@53745.4 package.scala 96:25:@53746.4]
  wire  _T_10399; // @[package.scala 96:25:@54129.4 package.scala 96:25:@54130.4]
  wire [7:0] _T_10403; // @[Mux.scala 31:69:@54139.4]
  wire  _T_10396; // @[package.scala 96:25:@54121.4 package.scala 96:25:@54122.4]
  wire [7:0] _T_10404; // @[Mux.scala 31:69:@54140.4]
  wire  _T_10393; // @[package.scala 96:25:@54113.4 package.scala 96:25:@54114.4]
  wire [7:0] _T_10405; // @[Mux.scala 31:69:@54141.4]
  wire  _T_10390; // @[package.scala 96:25:@54105.4 package.scala 96:25:@54106.4]
  wire [7:0] _T_10406; // @[Mux.scala 31:69:@54142.4]
  wire  _T_10387; // @[package.scala 96:25:@54097.4 package.scala 96:25:@54098.4]
  wire [7:0] _T_10407; // @[Mux.scala 31:69:@54143.4]
  wire  _T_10384; // @[package.scala 96:25:@54089.4 package.scala 96:25:@54090.4]
  wire [7:0] _T_10408; // @[Mux.scala 31:69:@54144.4]
  wire  _T_10381; // @[package.scala 96:25:@54081.4 package.scala 96:25:@54082.4]
  wire [7:0] _T_10409; // @[Mux.scala 31:69:@54145.4]
  wire  _T_10378; // @[package.scala 96:25:@54073.4 package.scala 96:25:@54074.4]
  wire [7:0] _T_10410; // @[Mux.scala 31:69:@54146.4]
  wire  _T_10375; // @[package.scala 96:25:@54065.4 package.scala 96:25:@54066.4]
  wire [7:0] _T_10411; // @[Mux.scala 31:69:@54147.4]
  wire  _T_10372; // @[package.scala 96:25:@54057.4 package.scala 96:25:@54058.4]
  wire [7:0] _T_10412; // @[Mux.scala 31:69:@54148.4]
  wire  _T_10369; // @[package.scala 96:25:@54049.4 package.scala 96:25:@54050.4]
  wire [7:0] _T_10413; // @[Mux.scala 31:69:@54149.4]
  wire  _T_10366; // @[package.scala 96:25:@54041.4 package.scala 96:25:@54042.4]
  wire [7:0] _T_10414; // @[Mux.scala 31:69:@54150.4]
  wire  _T_10363; // @[package.scala 96:25:@54033.4 package.scala 96:25:@54034.4]
  wire [7:0] _T_10415; // @[Mux.scala 31:69:@54151.4]
  wire  _T_10360; // @[package.scala 96:25:@54025.4 package.scala 96:25:@54026.4]
  wire [7:0] _T_10416; // @[Mux.scala 31:69:@54152.4]
  wire  _T_10357; // @[package.scala 96:25:@54017.4 package.scala 96:25:@54018.4]
  wire [7:0] _T_10417; // @[Mux.scala 31:69:@54153.4]
  wire  _T_10354; // @[package.scala 96:25:@54009.4 package.scala 96:25:@54010.4]
  wire [7:0] _T_10418; // @[Mux.scala 31:69:@54154.4]
  wire  _T_10351; // @[package.scala 96:25:@54001.4 package.scala 96:25:@54002.4]
  wire [7:0] _T_10419; // @[Mux.scala 31:69:@54155.4]
  wire  _T_10348; // @[package.scala 96:25:@53993.4 package.scala 96:25:@53994.4]
  wire [7:0] _T_10420; // @[Mux.scala 31:69:@54156.4]
  wire  _T_10345; // @[package.scala 96:25:@53985.4 package.scala 96:25:@53986.4]
  wire  _T_10578; // @[package.scala 96:25:@54369.4 package.scala 96:25:@54370.4]
  wire [7:0] _T_10582; // @[Mux.scala 31:69:@54379.4]
  wire  _T_10575; // @[package.scala 96:25:@54361.4 package.scala 96:25:@54362.4]
  wire [7:0] _T_10583; // @[Mux.scala 31:69:@54380.4]
  wire  _T_10572; // @[package.scala 96:25:@54353.4 package.scala 96:25:@54354.4]
  wire [7:0] _T_10584; // @[Mux.scala 31:69:@54381.4]
  wire  _T_10569; // @[package.scala 96:25:@54345.4 package.scala 96:25:@54346.4]
  wire [7:0] _T_10585; // @[Mux.scala 31:69:@54382.4]
  wire  _T_10566; // @[package.scala 96:25:@54337.4 package.scala 96:25:@54338.4]
  wire [7:0] _T_10586; // @[Mux.scala 31:69:@54383.4]
  wire  _T_10563; // @[package.scala 96:25:@54329.4 package.scala 96:25:@54330.4]
  wire [7:0] _T_10587; // @[Mux.scala 31:69:@54384.4]
  wire  _T_10560; // @[package.scala 96:25:@54321.4 package.scala 96:25:@54322.4]
  wire [7:0] _T_10588; // @[Mux.scala 31:69:@54385.4]
  wire  _T_10557; // @[package.scala 96:25:@54313.4 package.scala 96:25:@54314.4]
  wire [7:0] _T_10589; // @[Mux.scala 31:69:@54386.4]
  wire  _T_10554; // @[package.scala 96:25:@54305.4 package.scala 96:25:@54306.4]
  wire [7:0] _T_10590; // @[Mux.scala 31:69:@54387.4]
  wire  _T_10551; // @[package.scala 96:25:@54297.4 package.scala 96:25:@54298.4]
  wire [7:0] _T_10591; // @[Mux.scala 31:69:@54388.4]
  wire  _T_10548; // @[package.scala 96:25:@54289.4 package.scala 96:25:@54290.4]
  wire [7:0] _T_10592; // @[Mux.scala 31:69:@54389.4]
  wire  _T_10545; // @[package.scala 96:25:@54281.4 package.scala 96:25:@54282.4]
  wire [7:0] _T_10593; // @[Mux.scala 31:69:@54390.4]
  wire  _T_10542; // @[package.scala 96:25:@54273.4 package.scala 96:25:@54274.4]
  wire [7:0] _T_10594; // @[Mux.scala 31:69:@54391.4]
  wire  _T_10539; // @[package.scala 96:25:@54265.4 package.scala 96:25:@54266.4]
  wire [7:0] _T_10595; // @[Mux.scala 31:69:@54392.4]
  wire  _T_10536; // @[package.scala 96:25:@54257.4 package.scala 96:25:@54258.4]
  wire [7:0] _T_10596; // @[Mux.scala 31:69:@54393.4]
  wire  _T_10533; // @[package.scala 96:25:@54249.4 package.scala 96:25:@54250.4]
  wire [7:0] _T_10597; // @[Mux.scala 31:69:@54394.4]
  wire  _T_10530; // @[package.scala 96:25:@54241.4 package.scala 96:25:@54242.4]
  wire [7:0] _T_10598; // @[Mux.scala 31:69:@54395.4]
  wire  _T_10527; // @[package.scala 96:25:@54233.4 package.scala 96:25:@54234.4]
  wire [7:0] _T_10599; // @[Mux.scala 31:69:@54396.4]
  wire  _T_10524; // @[package.scala 96:25:@54225.4 package.scala 96:25:@54226.4]
  wire  _T_10757; // @[package.scala 96:25:@54609.4 package.scala 96:25:@54610.4]
  wire [7:0] _T_10761; // @[Mux.scala 31:69:@54619.4]
  wire  _T_10754; // @[package.scala 96:25:@54601.4 package.scala 96:25:@54602.4]
  wire [7:0] _T_10762; // @[Mux.scala 31:69:@54620.4]
  wire  _T_10751; // @[package.scala 96:25:@54593.4 package.scala 96:25:@54594.4]
  wire [7:0] _T_10763; // @[Mux.scala 31:69:@54621.4]
  wire  _T_10748; // @[package.scala 96:25:@54585.4 package.scala 96:25:@54586.4]
  wire [7:0] _T_10764; // @[Mux.scala 31:69:@54622.4]
  wire  _T_10745; // @[package.scala 96:25:@54577.4 package.scala 96:25:@54578.4]
  wire [7:0] _T_10765; // @[Mux.scala 31:69:@54623.4]
  wire  _T_10742; // @[package.scala 96:25:@54569.4 package.scala 96:25:@54570.4]
  wire [7:0] _T_10766; // @[Mux.scala 31:69:@54624.4]
  wire  _T_10739; // @[package.scala 96:25:@54561.4 package.scala 96:25:@54562.4]
  wire [7:0] _T_10767; // @[Mux.scala 31:69:@54625.4]
  wire  _T_10736; // @[package.scala 96:25:@54553.4 package.scala 96:25:@54554.4]
  wire [7:0] _T_10768; // @[Mux.scala 31:69:@54626.4]
  wire  _T_10733; // @[package.scala 96:25:@54545.4 package.scala 96:25:@54546.4]
  wire [7:0] _T_10769; // @[Mux.scala 31:69:@54627.4]
  wire  _T_10730; // @[package.scala 96:25:@54537.4 package.scala 96:25:@54538.4]
  wire [7:0] _T_10770; // @[Mux.scala 31:69:@54628.4]
  wire  _T_10727; // @[package.scala 96:25:@54529.4 package.scala 96:25:@54530.4]
  wire [7:0] _T_10771; // @[Mux.scala 31:69:@54629.4]
  wire  _T_10724; // @[package.scala 96:25:@54521.4 package.scala 96:25:@54522.4]
  wire [7:0] _T_10772; // @[Mux.scala 31:69:@54630.4]
  wire  _T_10721; // @[package.scala 96:25:@54513.4 package.scala 96:25:@54514.4]
  wire [7:0] _T_10773; // @[Mux.scala 31:69:@54631.4]
  wire  _T_10718; // @[package.scala 96:25:@54505.4 package.scala 96:25:@54506.4]
  wire [7:0] _T_10774; // @[Mux.scala 31:69:@54632.4]
  wire  _T_10715; // @[package.scala 96:25:@54497.4 package.scala 96:25:@54498.4]
  wire [7:0] _T_10775; // @[Mux.scala 31:69:@54633.4]
  wire  _T_10712; // @[package.scala 96:25:@54489.4 package.scala 96:25:@54490.4]
  wire [7:0] _T_10776; // @[Mux.scala 31:69:@54634.4]
  wire  _T_10709; // @[package.scala 96:25:@54481.4 package.scala 96:25:@54482.4]
  wire [7:0] _T_10777; // @[Mux.scala 31:69:@54635.4]
  wire  _T_10706; // @[package.scala 96:25:@54473.4 package.scala 96:25:@54474.4]
  wire [7:0] _T_10778; // @[Mux.scala 31:69:@54636.4]
  wire  _T_10703; // @[package.scala 96:25:@54465.4 package.scala 96:25:@54466.4]
  wire  _T_10936; // @[package.scala 96:25:@54849.4 package.scala 96:25:@54850.4]
  wire [7:0] _T_10940; // @[Mux.scala 31:69:@54859.4]
  wire  _T_10933; // @[package.scala 96:25:@54841.4 package.scala 96:25:@54842.4]
  wire [7:0] _T_10941; // @[Mux.scala 31:69:@54860.4]
  wire  _T_10930; // @[package.scala 96:25:@54833.4 package.scala 96:25:@54834.4]
  wire [7:0] _T_10942; // @[Mux.scala 31:69:@54861.4]
  wire  _T_10927; // @[package.scala 96:25:@54825.4 package.scala 96:25:@54826.4]
  wire [7:0] _T_10943; // @[Mux.scala 31:69:@54862.4]
  wire  _T_10924; // @[package.scala 96:25:@54817.4 package.scala 96:25:@54818.4]
  wire [7:0] _T_10944; // @[Mux.scala 31:69:@54863.4]
  wire  _T_10921; // @[package.scala 96:25:@54809.4 package.scala 96:25:@54810.4]
  wire [7:0] _T_10945; // @[Mux.scala 31:69:@54864.4]
  wire  _T_10918; // @[package.scala 96:25:@54801.4 package.scala 96:25:@54802.4]
  wire [7:0] _T_10946; // @[Mux.scala 31:69:@54865.4]
  wire  _T_10915; // @[package.scala 96:25:@54793.4 package.scala 96:25:@54794.4]
  wire [7:0] _T_10947; // @[Mux.scala 31:69:@54866.4]
  wire  _T_10912; // @[package.scala 96:25:@54785.4 package.scala 96:25:@54786.4]
  wire [7:0] _T_10948; // @[Mux.scala 31:69:@54867.4]
  wire  _T_10909; // @[package.scala 96:25:@54777.4 package.scala 96:25:@54778.4]
  wire [7:0] _T_10949; // @[Mux.scala 31:69:@54868.4]
  wire  _T_10906; // @[package.scala 96:25:@54769.4 package.scala 96:25:@54770.4]
  wire [7:0] _T_10950; // @[Mux.scala 31:69:@54869.4]
  wire  _T_10903; // @[package.scala 96:25:@54761.4 package.scala 96:25:@54762.4]
  wire [7:0] _T_10951; // @[Mux.scala 31:69:@54870.4]
  wire  _T_10900; // @[package.scala 96:25:@54753.4 package.scala 96:25:@54754.4]
  wire [7:0] _T_10952; // @[Mux.scala 31:69:@54871.4]
  wire  _T_10897; // @[package.scala 96:25:@54745.4 package.scala 96:25:@54746.4]
  wire [7:0] _T_10953; // @[Mux.scala 31:69:@54872.4]
  wire  _T_10894; // @[package.scala 96:25:@54737.4 package.scala 96:25:@54738.4]
  wire [7:0] _T_10954; // @[Mux.scala 31:69:@54873.4]
  wire  _T_10891; // @[package.scala 96:25:@54729.4 package.scala 96:25:@54730.4]
  wire [7:0] _T_10955; // @[Mux.scala 31:69:@54874.4]
  wire  _T_10888; // @[package.scala 96:25:@54721.4 package.scala 96:25:@54722.4]
  wire [7:0] _T_10956; // @[Mux.scala 31:69:@54875.4]
  wire  _T_10885; // @[package.scala 96:25:@54713.4 package.scala 96:25:@54714.4]
  wire [7:0] _T_10957; // @[Mux.scala 31:69:@54876.4]
  wire  _T_10882; // @[package.scala 96:25:@54705.4 package.scala 96:25:@54706.4]
  wire  _T_11115; // @[package.scala 96:25:@55089.4 package.scala 96:25:@55090.4]
  wire [7:0] _T_11119; // @[Mux.scala 31:69:@55099.4]
  wire  _T_11112; // @[package.scala 96:25:@55081.4 package.scala 96:25:@55082.4]
  wire [7:0] _T_11120; // @[Mux.scala 31:69:@55100.4]
  wire  _T_11109; // @[package.scala 96:25:@55073.4 package.scala 96:25:@55074.4]
  wire [7:0] _T_11121; // @[Mux.scala 31:69:@55101.4]
  wire  _T_11106; // @[package.scala 96:25:@55065.4 package.scala 96:25:@55066.4]
  wire [7:0] _T_11122; // @[Mux.scala 31:69:@55102.4]
  wire  _T_11103; // @[package.scala 96:25:@55057.4 package.scala 96:25:@55058.4]
  wire [7:0] _T_11123; // @[Mux.scala 31:69:@55103.4]
  wire  _T_11100; // @[package.scala 96:25:@55049.4 package.scala 96:25:@55050.4]
  wire [7:0] _T_11124; // @[Mux.scala 31:69:@55104.4]
  wire  _T_11097; // @[package.scala 96:25:@55041.4 package.scala 96:25:@55042.4]
  wire [7:0] _T_11125; // @[Mux.scala 31:69:@55105.4]
  wire  _T_11094; // @[package.scala 96:25:@55033.4 package.scala 96:25:@55034.4]
  wire [7:0] _T_11126; // @[Mux.scala 31:69:@55106.4]
  wire  _T_11091; // @[package.scala 96:25:@55025.4 package.scala 96:25:@55026.4]
  wire [7:0] _T_11127; // @[Mux.scala 31:69:@55107.4]
  wire  _T_11088; // @[package.scala 96:25:@55017.4 package.scala 96:25:@55018.4]
  wire [7:0] _T_11128; // @[Mux.scala 31:69:@55108.4]
  wire  _T_11085; // @[package.scala 96:25:@55009.4 package.scala 96:25:@55010.4]
  wire [7:0] _T_11129; // @[Mux.scala 31:69:@55109.4]
  wire  _T_11082; // @[package.scala 96:25:@55001.4 package.scala 96:25:@55002.4]
  wire [7:0] _T_11130; // @[Mux.scala 31:69:@55110.4]
  wire  _T_11079; // @[package.scala 96:25:@54993.4 package.scala 96:25:@54994.4]
  wire [7:0] _T_11131; // @[Mux.scala 31:69:@55111.4]
  wire  _T_11076; // @[package.scala 96:25:@54985.4 package.scala 96:25:@54986.4]
  wire [7:0] _T_11132; // @[Mux.scala 31:69:@55112.4]
  wire  _T_11073; // @[package.scala 96:25:@54977.4 package.scala 96:25:@54978.4]
  wire [7:0] _T_11133; // @[Mux.scala 31:69:@55113.4]
  wire  _T_11070; // @[package.scala 96:25:@54969.4 package.scala 96:25:@54970.4]
  wire [7:0] _T_11134; // @[Mux.scala 31:69:@55114.4]
  wire  _T_11067; // @[package.scala 96:25:@54961.4 package.scala 96:25:@54962.4]
  wire [7:0] _T_11135; // @[Mux.scala 31:69:@55115.4]
  wire  _T_11064; // @[package.scala 96:25:@54953.4 package.scala 96:25:@54954.4]
  wire [7:0] _T_11136; // @[Mux.scala 31:69:@55116.4]
  wire  _T_11061; // @[package.scala 96:25:@54945.4 package.scala 96:25:@54946.4]
  wire  _T_11294; // @[package.scala 96:25:@55329.4 package.scala 96:25:@55330.4]
  wire [7:0] _T_11298; // @[Mux.scala 31:69:@55339.4]
  wire  _T_11291; // @[package.scala 96:25:@55321.4 package.scala 96:25:@55322.4]
  wire [7:0] _T_11299; // @[Mux.scala 31:69:@55340.4]
  wire  _T_11288; // @[package.scala 96:25:@55313.4 package.scala 96:25:@55314.4]
  wire [7:0] _T_11300; // @[Mux.scala 31:69:@55341.4]
  wire  _T_11285; // @[package.scala 96:25:@55305.4 package.scala 96:25:@55306.4]
  wire [7:0] _T_11301; // @[Mux.scala 31:69:@55342.4]
  wire  _T_11282; // @[package.scala 96:25:@55297.4 package.scala 96:25:@55298.4]
  wire [7:0] _T_11302; // @[Mux.scala 31:69:@55343.4]
  wire  _T_11279; // @[package.scala 96:25:@55289.4 package.scala 96:25:@55290.4]
  wire [7:0] _T_11303; // @[Mux.scala 31:69:@55344.4]
  wire  _T_11276; // @[package.scala 96:25:@55281.4 package.scala 96:25:@55282.4]
  wire [7:0] _T_11304; // @[Mux.scala 31:69:@55345.4]
  wire  _T_11273; // @[package.scala 96:25:@55273.4 package.scala 96:25:@55274.4]
  wire [7:0] _T_11305; // @[Mux.scala 31:69:@55346.4]
  wire  _T_11270; // @[package.scala 96:25:@55265.4 package.scala 96:25:@55266.4]
  wire [7:0] _T_11306; // @[Mux.scala 31:69:@55347.4]
  wire  _T_11267; // @[package.scala 96:25:@55257.4 package.scala 96:25:@55258.4]
  wire [7:0] _T_11307; // @[Mux.scala 31:69:@55348.4]
  wire  _T_11264; // @[package.scala 96:25:@55249.4 package.scala 96:25:@55250.4]
  wire [7:0] _T_11308; // @[Mux.scala 31:69:@55349.4]
  wire  _T_11261; // @[package.scala 96:25:@55241.4 package.scala 96:25:@55242.4]
  wire [7:0] _T_11309; // @[Mux.scala 31:69:@55350.4]
  wire  _T_11258; // @[package.scala 96:25:@55233.4 package.scala 96:25:@55234.4]
  wire [7:0] _T_11310; // @[Mux.scala 31:69:@55351.4]
  wire  _T_11255; // @[package.scala 96:25:@55225.4 package.scala 96:25:@55226.4]
  wire [7:0] _T_11311; // @[Mux.scala 31:69:@55352.4]
  wire  _T_11252; // @[package.scala 96:25:@55217.4 package.scala 96:25:@55218.4]
  wire [7:0] _T_11312; // @[Mux.scala 31:69:@55353.4]
  wire  _T_11249; // @[package.scala 96:25:@55209.4 package.scala 96:25:@55210.4]
  wire [7:0] _T_11313; // @[Mux.scala 31:69:@55354.4]
  wire  _T_11246; // @[package.scala 96:25:@55201.4 package.scala 96:25:@55202.4]
  wire [7:0] _T_11314; // @[Mux.scala 31:69:@55355.4]
  wire  _T_11243; // @[package.scala 96:25:@55193.4 package.scala 96:25:@55194.4]
  wire [7:0] _T_11315; // @[Mux.scala 31:69:@55356.4]
  wire  _T_11240; // @[package.scala 96:25:@55185.4 package.scala 96:25:@55186.4]
  wire  _T_11473; // @[package.scala 96:25:@55569.4 package.scala 96:25:@55570.4]
  wire [7:0] _T_11477; // @[Mux.scala 31:69:@55579.4]
  wire  _T_11470; // @[package.scala 96:25:@55561.4 package.scala 96:25:@55562.4]
  wire [7:0] _T_11478; // @[Mux.scala 31:69:@55580.4]
  wire  _T_11467; // @[package.scala 96:25:@55553.4 package.scala 96:25:@55554.4]
  wire [7:0] _T_11479; // @[Mux.scala 31:69:@55581.4]
  wire  _T_11464; // @[package.scala 96:25:@55545.4 package.scala 96:25:@55546.4]
  wire [7:0] _T_11480; // @[Mux.scala 31:69:@55582.4]
  wire  _T_11461; // @[package.scala 96:25:@55537.4 package.scala 96:25:@55538.4]
  wire [7:0] _T_11481; // @[Mux.scala 31:69:@55583.4]
  wire  _T_11458; // @[package.scala 96:25:@55529.4 package.scala 96:25:@55530.4]
  wire [7:0] _T_11482; // @[Mux.scala 31:69:@55584.4]
  wire  _T_11455; // @[package.scala 96:25:@55521.4 package.scala 96:25:@55522.4]
  wire [7:0] _T_11483; // @[Mux.scala 31:69:@55585.4]
  wire  _T_11452; // @[package.scala 96:25:@55513.4 package.scala 96:25:@55514.4]
  wire [7:0] _T_11484; // @[Mux.scala 31:69:@55586.4]
  wire  _T_11449; // @[package.scala 96:25:@55505.4 package.scala 96:25:@55506.4]
  wire [7:0] _T_11485; // @[Mux.scala 31:69:@55587.4]
  wire  _T_11446; // @[package.scala 96:25:@55497.4 package.scala 96:25:@55498.4]
  wire [7:0] _T_11486; // @[Mux.scala 31:69:@55588.4]
  wire  _T_11443; // @[package.scala 96:25:@55489.4 package.scala 96:25:@55490.4]
  wire [7:0] _T_11487; // @[Mux.scala 31:69:@55589.4]
  wire  _T_11440; // @[package.scala 96:25:@55481.4 package.scala 96:25:@55482.4]
  wire [7:0] _T_11488; // @[Mux.scala 31:69:@55590.4]
  wire  _T_11437; // @[package.scala 96:25:@55473.4 package.scala 96:25:@55474.4]
  wire [7:0] _T_11489; // @[Mux.scala 31:69:@55591.4]
  wire  _T_11434; // @[package.scala 96:25:@55465.4 package.scala 96:25:@55466.4]
  wire [7:0] _T_11490; // @[Mux.scala 31:69:@55592.4]
  wire  _T_11431; // @[package.scala 96:25:@55457.4 package.scala 96:25:@55458.4]
  wire [7:0] _T_11491; // @[Mux.scala 31:69:@55593.4]
  wire  _T_11428; // @[package.scala 96:25:@55449.4 package.scala 96:25:@55450.4]
  wire [7:0] _T_11492; // @[Mux.scala 31:69:@55594.4]
  wire  _T_11425; // @[package.scala 96:25:@55441.4 package.scala 96:25:@55442.4]
  wire [7:0] _T_11493; // @[Mux.scala 31:69:@55595.4]
  wire  _T_11422; // @[package.scala 96:25:@55433.4 package.scala 96:25:@55434.4]
  wire [7:0] _T_11494; // @[Mux.scala 31:69:@55596.4]
  wire  _T_11419; // @[package.scala 96:25:@55425.4 package.scala 96:25:@55426.4]
  wire  _T_11652; // @[package.scala 96:25:@55809.4 package.scala 96:25:@55810.4]
  wire [7:0] _T_11656; // @[Mux.scala 31:69:@55819.4]
  wire  _T_11649; // @[package.scala 96:25:@55801.4 package.scala 96:25:@55802.4]
  wire [7:0] _T_11657; // @[Mux.scala 31:69:@55820.4]
  wire  _T_11646; // @[package.scala 96:25:@55793.4 package.scala 96:25:@55794.4]
  wire [7:0] _T_11658; // @[Mux.scala 31:69:@55821.4]
  wire  _T_11643; // @[package.scala 96:25:@55785.4 package.scala 96:25:@55786.4]
  wire [7:0] _T_11659; // @[Mux.scala 31:69:@55822.4]
  wire  _T_11640; // @[package.scala 96:25:@55777.4 package.scala 96:25:@55778.4]
  wire [7:0] _T_11660; // @[Mux.scala 31:69:@55823.4]
  wire  _T_11637; // @[package.scala 96:25:@55769.4 package.scala 96:25:@55770.4]
  wire [7:0] _T_11661; // @[Mux.scala 31:69:@55824.4]
  wire  _T_11634; // @[package.scala 96:25:@55761.4 package.scala 96:25:@55762.4]
  wire [7:0] _T_11662; // @[Mux.scala 31:69:@55825.4]
  wire  _T_11631; // @[package.scala 96:25:@55753.4 package.scala 96:25:@55754.4]
  wire [7:0] _T_11663; // @[Mux.scala 31:69:@55826.4]
  wire  _T_11628; // @[package.scala 96:25:@55745.4 package.scala 96:25:@55746.4]
  wire [7:0] _T_11664; // @[Mux.scala 31:69:@55827.4]
  wire  _T_11625; // @[package.scala 96:25:@55737.4 package.scala 96:25:@55738.4]
  wire [7:0] _T_11665; // @[Mux.scala 31:69:@55828.4]
  wire  _T_11622; // @[package.scala 96:25:@55729.4 package.scala 96:25:@55730.4]
  wire [7:0] _T_11666; // @[Mux.scala 31:69:@55829.4]
  wire  _T_11619; // @[package.scala 96:25:@55721.4 package.scala 96:25:@55722.4]
  wire [7:0] _T_11667; // @[Mux.scala 31:69:@55830.4]
  wire  _T_11616; // @[package.scala 96:25:@55713.4 package.scala 96:25:@55714.4]
  wire [7:0] _T_11668; // @[Mux.scala 31:69:@55831.4]
  wire  _T_11613; // @[package.scala 96:25:@55705.4 package.scala 96:25:@55706.4]
  wire [7:0] _T_11669; // @[Mux.scala 31:69:@55832.4]
  wire  _T_11610; // @[package.scala 96:25:@55697.4 package.scala 96:25:@55698.4]
  wire [7:0] _T_11670; // @[Mux.scala 31:69:@55833.4]
  wire  _T_11607; // @[package.scala 96:25:@55689.4 package.scala 96:25:@55690.4]
  wire [7:0] _T_11671; // @[Mux.scala 31:69:@55834.4]
  wire  _T_11604; // @[package.scala 96:25:@55681.4 package.scala 96:25:@55682.4]
  wire [7:0] _T_11672; // @[Mux.scala 31:69:@55835.4]
  wire  _T_11601; // @[package.scala 96:25:@55673.4 package.scala 96:25:@55674.4]
  wire [7:0] _T_11673; // @[Mux.scala 31:69:@55836.4]
  wire  _T_11598; // @[package.scala 96:25:@55665.4 package.scala 96:25:@55666.4]
  wire  _T_11831; // @[package.scala 96:25:@56049.4 package.scala 96:25:@56050.4]
  wire [7:0] _T_11835; // @[Mux.scala 31:69:@56059.4]
  wire  _T_11828; // @[package.scala 96:25:@56041.4 package.scala 96:25:@56042.4]
  wire [7:0] _T_11836; // @[Mux.scala 31:69:@56060.4]
  wire  _T_11825; // @[package.scala 96:25:@56033.4 package.scala 96:25:@56034.4]
  wire [7:0] _T_11837; // @[Mux.scala 31:69:@56061.4]
  wire  _T_11822; // @[package.scala 96:25:@56025.4 package.scala 96:25:@56026.4]
  wire [7:0] _T_11838; // @[Mux.scala 31:69:@56062.4]
  wire  _T_11819; // @[package.scala 96:25:@56017.4 package.scala 96:25:@56018.4]
  wire [7:0] _T_11839; // @[Mux.scala 31:69:@56063.4]
  wire  _T_11816; // @[package.scala 96:25:@56009.4 package.scala 96:25:@56010.4]
  wire [7:0] _T_11840; // @[Mux.scala 31:69:@56064.4]
  wire  _T_11813; // @[package.scala 96:25:@56001.4 package.scala 96:25:@56002.4]
  wire [7:0] _T_11841; // @[Mux.scala 31:69:@56065.4]
  wire  _T_11810; // @[package.scala 96:25:@55993.4 package.scala 96:25:@55994.4]
  wire [7:0] _T_11842; // @[Mux.scala 31:69:@56066.4]
  wire  _T_11807; // @[package.scala 96:25:@55985.4 package.scala 96:25:@55986.4]
  wire [7:0] _T_11843; // @[Mux.scala 31:69:@56067.4]
  wire  _T_11804; // @[package.scala 96:25:@55977.4 package.scala 96:25:@55978.4]
  wire [7:0] _T_11844; // @[Mux.scala 31:69:@56068.4]
  wire  _T_11801; // @[package.scala 96:25:@55969.4 package.scala 96:25:@55970.4]
  wire [7:0] _T_11845; // @[Mux.scala 31:69:@56069.4]
  wire  _T_11798; // @[package.scala 96:25:@55961.4 package.scala 96:25:@55962.4]
  wire [7:0] _T_11846; // @[Mux.scala 31:69:@56070.4]
  wire  _T_11795; // @[package.scala 96:25:@55953.4 package.scala 96:25:@55954.4]
  wire [7:0] _T_11847; // @[Mux.scala 31:69:@56071.4]
  wire  _T_11792; // @[package.scala 96:25:@55945.4 package.scala 96:25:@55946.4]
  wire [7:0] _T_11848; // @[Mux.scala 31:69:@56072.4]
  wire  _T_11789; // @[package.scala 96:25:@55937.4 package.scala 96:25:@55938.4]
  wire [7:0] _T_11849; // @[Mux.scala 31:69:@56073.4]
  wire  _T_11786; // @[package.scala 96:25:@55929.4 package.scala 96:25:@55930.4]
  wire [7:0] _T_11850; // @[Mux.scala 31:69:@56074.4]
  wire  _T_11783; // @[package.scala 96:25:@55921.4 package.scala 96:25:@55922.4]
  wire [7:0] _T_11851; // @[Mux.scala 31:69:@56075.4]
  wire  _T_11780; // @[package.scala 96:25:@55913.4 package.scala 96:25:@55914.4]
  wire [7:0] _T_11852; // @[Mux.scala 31:69:@56076.4]
  wire  _T_11777; // @[package.scala 96:25:@55905.4 package.scala 96:25:@55906.4]
  wire  _T_12010; // @[package.scala 96:25:@56289.4 package.scala 96:25:@56290.4]
  wire [7:0] _T_12014; // @[Mux.scala 31:69:@56299.4]
  wire  _T_12007; // @[package.scala 96:25:@56281.4 package.scala 96:25:@56282.4]
  wire [7:0] _T_12015; // @[Mux.scala 31:69:@56300.4]
  wire  _T_12004; // @[package.scala 96:25:@56273.4 package.scala 96:25:@56274.4]
  wire [7:0] _T_12016; // @[Mux.scala 31:69:@56301.4]
  wire  _T_12001; // @[package.scala 96:25:@56265.4 package.scala 96:25:@56266.4]
  wire [7:0] _T_12017; // @[Mux.scala 31:69:@56302.4]
  wire  _T_11998; // @[package.scala 96:25:@56257.4 package.scala 96:25:@56258.4]
  wire [7:0] _T_12018; // @[Mux.scala 31:69:@56303.4]
  wire  _T_11995; // @[package.scala 96:25:@56249.4 package.scala 96:25:@56250.4]
  wire [7:0] _T_12019; // @[Mux.scala 31:69:@56304.4]
  wire  _T_11992; // @[package.scala 96:25:@56241.4 package.scala 96:25:@56242.4]
  wire [7:0] _T_12020; // @[Mux.scala 31:69:@56305.4]
  wire  _T_11989; // @[package.scala 96:25:@56233.4 package.scala 96:25:@56234.4]
  wire [7:0] _T_12021; // @[Mux.scala 31:69:@56306.4]
  wire  _T_11986; // @[package.scala 96:25:@56225.4 package.scala 96:25:@56226.4]
  wire [7:0] _T_12022; // @[Mux.scala 31:69:@56307.4]
  wire  _T_11983; // @[package.scala 96:25:@56217.4 package.scala 96:25:@56218.4]
  wire [7:0] _T_12023; // @[Mux.scala 31:69:@56308.4]
  wire  _T_11980; // @[package.scala 96:25:@56209.4 package.scala 96:25:@56210.4]
  wire [7:0] _T_12024; // @[Mux.scala 31:69:@56309.4]
  wire  _T_11977; // @[package.scala 96:25:@56201.4 package.scala 96:25:@56202.4]
  wire [7:0] _T_12025; // @[Mux.scala 31:69:@56310.4]
  wire  _T_11974; // @[package.scala 96:25:@56193.4 package.scala 96:25:@56194.4]
  wire [7:0] _T_12026; // @[Mux.scala 31:69:@56311.4]
  wire  _T_11971; // @[package.scala 96:25:@56185.4 package.scala 96:25:@56186.4]
  wire [7:0] _T_12027; // @[Mux.scala 31:69:@56312.4]
  wire  _T_11968; // @[package.scala 96:25:@56177.4 package.scala 96:25:@56178.4]
  wire [7:0] _T_12028; // @[Mux.scala 31:69:@56313.4]
  wire  _T_11965; // @[package.scala 96:25:@56169.4 package.scala 96:25:@56170.4]
  wire [7:0] _T_12029; // @[Mux.scala 31:69:@56314.4]
  wire  _T_11962; // @[package.scala 96:25:@56161.4 package.scala 96:25:@56162.4]
  wire [7:0] _T_12030; // @[Mux.scala 31:69:@56315.4]
  wire  _T_11959; // @[package.scala 96:25:@56153.4 package.scala 96:25:@56154.4]
  wire [7:0] _T_12031; // @[Mux.scala 31:69:@56316.4]
  wire  _T_11956; // @[package.scala 96:25:@56145.4 package.scala 96:25:@56146.4]
  wire  _T_12189; // @[package.scala 96:25:@56529.4 package.scala 96:25:@56530.4]
  wire [7:0] _T_12193; // @[Mux.scala 31:69:@56539.4]
  wire  _T_12186; // @[package.scala 96:25:@56521.4 package.scala 96:25:@56522.4]
  wire [7:0] _T_12194; // @[Mux.scala 31:69:@56540.4]
  wire  _T_12183; // @[package.scala 96:25:@56513.4 package.scala 96:25:@56514.4]
  wire [7:0] _T_12195; // @[Mux.scala 31:69:@56541.4]
  wire  _T_12180; // @[package.scala 96:25:@56505.4 package.scala 96:25:@56506.4]
  wire [7:0] _T_12196; // @[Mux.scala 31:69:@56542.4]
  wire  _T_12177; // @[package.scala 96:25:@56497.4 package.scala 96:25:@56498.4]
  wire [7:0] _T_12197; // @[Mux.scala 31:69:@56543.4]
  wire  _T_12174; // @[package.scala 96:25:@56489.4 package.scala 96:25:@56490.4]
  wire [7:0] _T_12198; // @[Mux.scala 31:69:@56544.4]
  wire  _T_12171; // @[package.scala 96:25:@56481.4 package.scala 96:25:@56482.4]
  wire [7:0] _T_12199; // @[Mux.scala 31:69:@56545.4]
  wire  _T_12168; // @[package.scala 96:25:@56473.4 package.scala 96:25:@56474.4]
  wire [7:0] _T_12200; // @[Mux.scala 31:69:@56546.4]
  wire  _T_12165; // @[package.scala 96:25:@56465.4 package.scala 96:25:@56466.4]
  wire [7:0] _T_12201; // @[Mux.scala 31:69:@56547.4]
  wire  _T_12162; // @[package.scala 96:25:@56457.4 package.scala 96:25:@56458.4]
  wire [7:0] _T_12202; // @[Mux.scala 31:69:@56548.4]
  wire  _T_12159; // @[package.scala 96:25:@56449.4 package.scala 96:25:@56450.4]
  wire [7:0] _T_12203; // @[Mux.scala 31:69:@56549.4]
  wire  _T_12156; // @[package.scala 96:25:@56441.4 package.scala 96:25:@56442.4]
  wire [7:0] _T_12204; // @[Mux.scala 31:69:@56550.4]
  wire  _T_12153; // @[package.scala 96:25:@56433.4 package.scala 96:25:@56434.4]
  wire [7:0] _T_12205; // @[Mux.scala 31:69:@56551.4]
  wire  _T_12150; // @[package.scala 96:25:@56425.4 package.scala 96:25:@56426.4]
  wire [7:0] _T_12206; // @[Mux.scala 31:69:@56552.4]
  wire  _T_12147; // @[package.scala 96:25:@56417.4 package.scala 96:25:@56418.4]
  wire [7:0] _T_12207; // @[Mux.scala 31:69:@56553.4]
  wire  _T_12144; // @[package.scala 96:25:@56409.4 package.scala 96:25:@56410.4]
  wire [7:0] _T_12208; // @[Mux.scala 31:69:@56554.4]
  wire  _T_12141; // @[package.scala 96:25:@56401.4 package.scala 96:25:@56402.4]
  wire [7:0] _T_12209; // @[Mux.scala 31:69:@56555.4]
  wire  _T_12138; // @[package.scala 96:25:@56393.4 package.scala 96:25:@56394.4]
  wire [7:0] _T_12210; // @[Mux.scala 31:69:@56556.4]
  wire  _T_12135; // @[package.scala 96:25:@56385.4 package.scala 96:25:@56386.4]
  wire  _T_12368; // @[package.scala 96:25:@56769.4 package.scala 96:25:@56770.4]
  wire [7:0] _T_12372; // @[Mux.scala 31:69:@56779.4]
  wire  _T_12365; // @[package.scala 96:25:@56761.4 package.scala 96:25:@56762.4]
  wire [7:0] _T_12373; // @[Mux.scala 31:69:@56780.4]
  wire  _T_12362; // @[package.scala 96:25:@56753.4 package.scala 96:25:@56754.4]
  wire [7:0] _T_12374; // @[Mux.scala 31:69:@56781.4]
  wire  _T_12359; // @[package.scala 96:25:@56745.4 package.scala 96:25:@56746.4]
  wire [7:0] _T_12375; // @[Mux.scala 31:69:@56782.4]
  wire  _T_12356; // @[package.scala 96:25:@56737.4 package.scala 96:25:@56738.4]
  wire [7:0] _T_12376; // @[Mux.scala 31:69:@56783.4]
  wire  _T_12353; // @[package.scala 96:25:@56729.4 package.scala 96:25:@56730.4]
  wire [7:0] _T_12377; // @[Mux.scala 31:69:@56784.4]
  wire  _T_12350; // @[package.scala 96:25:@56721.4 package.scala 96:25:@56722.4]
  wire [7:0] _T_12378; // @[Mux.scala 31:69:@56785.4]
  wire  _T_12347; // @[package.scala 96:25:@56713.4 package.scala 96:25:@56714.4]
  wire [7:0] _T_12379; // @[Mux.scala 31:69:@56786.4]
  wire  _T_12344; // @[package.scala 96:25:@56705.4 package.scala 96:25:@56706.4]
  wire [7:0] _T_12380; // @[Mux.scala 31:69:@56787.4]
  wire  _T_12341; // @[package.scala 96:25:@56697.4 package.scala 96:25:@56698.4]
  wire [7:0] _T_12381; // @[Mux.scala 31:69:@56788.4]
  wire  _T_12338; // @[package.scala 96:25:@56689.4 package.scala 96:25:@56690.4]
  wire [7:0] _T_12382; // @[Mux.scala 31:69:@56789.4]
  wire  _T_12335; // @[package.scala 96:25:@56681.4 package.scala 96:25:@56682.4]
  wire [7:0] _T_12383; // @[Mux.scala 31:69:@56790.4]
  wire  _T_12332; // @[package.scala 96:25:@56673.4 package.scala 96:25:@56674.4]
  wire [7:0] _T_12384; // @[Mux.scala 31:69:@56791.4]
  wire  _T_12329; // @[package.scala 96:25:@56665.4 package.scala 96:25:@56666.4]
  wire [7:0] _T_12385; // @[Mux.scala 31:69:@56792.4]
  wire  _T_12326; // @[package.scala 96:25:@56657.4 package.scala 96:25:@56658.4]
  wire [7:0] _T_12386; // @[Mux.scala 31:69:@56793.4]
  wire  _T_12323; // @[package.scala 96:25:@56649.4 package.scala 96:25:@56650.4]
  wire [7:0] _T_12387; // @[Mux.scala 31:69:@56794.4]
  wire  _T_12320; // @[package.scala 96:25:@56641.4 package.scala 96:25:@56642.4]
  wire [7:0] _T_12388; // @[Mux.scala 31:69:@56795.4]
  wire  _T_12317; // @[package.scala 96:25:@56633.4 package.scala 96:25:@56634.4]
  wire [7:0] _T_12389; // @[Mux.scala 31:69:@56796.4]
  wire  _T_12314; // @[package.scala 96:25:@56625.4 package.scala 96:25:@56626.4]
  wire  _T_12547; // @[package.scala 96:25:@57009.4 package.scala 96:25:@57010.4]
  wire [7:0] _T_12551; // @[Mux.scala 31:69:@57019.4]
  wire  _T_12544; // @[package.scala 96:25:@57001.4 package.scala 96:25:@57002.4]
  wire [7:0] _T_12552; // @[Mux.scala 31:69:@57020.4]
  wire  _T_12541; // @[package.scala 96:25:@56993.4 package.scala 96:25:@56994.4]
  wire [7:0] _T_12553; // @[Mux.scala 31:69:@57021.4]
  wire  _T_12538; // @[package.scala 96:25:@56985.4 package.scala 96:25:@56986.4]
  wire [7:0] _T_12554; // @[Mux.scala 31:69:@57022.4]
  wire  _T_12535; // @[package.scala 96:25:@56977.4 package.scala 96:25:@56978.4]
  wire [7:0] _T_12555; // @[Mux.scala 31:69:@57023.4]
  wire  _T_12532; // @[package.scala 96:25:@56969.4 package.scala 96:25:@56970.4]
  wire [7:0] _T_12556; // @[Mux.scala 31:69:@57024.4]
  wire  _T_12529; // @[package.scala 96:25:@56961.4 package.scala 96:25:@56962.4]
  wire [7:0] _T_12557; // @[Mux.scala 31:69:@57025.4]
  wire  _T_12526; // @[package.scala 96:25:@56953.4 package.scala 96:25:@56954.4]
  wire [7:0] _T_12558; // @[Mux.scala 31:69:@57026.4]
  wire  _T_12523; // @[package.scala 96:25:@56945.4 package.scala 96:25:@56946.4]
  wire [7:0] _T_12559; // @[Mux.scala 31:69:@57027.4]
  wire  _T_12520; // @[package.scala 96:25:@56937.4 package.scala 96:25:@56938.4]
  wire [7:0] _T_12560; // @[Mux.scala 31:69:@57028.4]
  wire  _T_12517; // @[package.scala 96:25:@56929.4 package.scala 96:25:@56930.4]
  wire [7:0] _T_12561; // @[Mux.scala 31:69:@57029.4]
  wire  _T_12514; // @[package.scala 96:25:@56921.4 package.scala 96:25:@56922.4]
  wire [7:0] _T_12562; // @[Mux.scala 31:69:@57030.4]
  wire  _T_12511; // @[package.scala 96:25:@56913.4 package.scala 96:25:@56914.4]
  wire [7:0] _T_12563; // @[Mux.scala 31:69:@57031.4]
  wire  _T_12508; // @[package.scala 96:25:@56905.4 package.scala 96:25:@56906.4]
  wire [7:0] _T_12564; // @[Mux.scala 31:69:@57032.4]
  wire  _T_12505; // @[package.scala 96:25:@56897.4 package.scala 96:25:@56898.4]
  wire [7:0] _T_12565; // @[Mux.scala 31:69:@57033.4]
  wire  _T_12502; // @[package.scala 96:25:@56889.4 package.scala 96:25:@56890.4]
  wire [7:0] _T_12566; // @[Mux.scala 31:69:@57034.4]
  wire  _T_12499; // @[package.scala 96:25:@56881.4 package.scala 96:25:@56882.4]
  wire [7:0] _T_12567; // @[Mux.scala 31:69:@57035.4]
  wire  _T_12496; // @[package.scala 96:25:@56873.4 package.scala 96:25:@56874.4]
  wire [7:0] _T_12568; // @[Mux.scala 31:69:@57036.4]
  wire  _T_12493; // @[package.scala 96:25:@56865.4 package.scala 96:25:@56866.4]
  wire  _T_12726; // @[package.scala 96:25:@57249.4 package.scala 96:25:@57250.4]
  wire [7:0] _T_12730; // @[Mux.scala 31:69:@57259.4]
  wire  _T_12723; // @[package.scala 96:25:@57241.4 package.scala 96:25:@57242.4]
  wire [7:0] _T_12731; // @[Mux.scala 31:69:@57260.4]
  wire  _T_12720; // @[package.scala 96:25:@57233.4 package.scala 96:25:@57234.4]
  wire [7:0] _T_12732; // @[Mux.scala 31:69:@57261.4]
  wire  _T_12717; // @[package.scala 96:25:@57225.4 package.scala 96:25:@57226.4]
  wire [7:0] _T_12733; // @[Mux.scala 31:69:@57262.4]
  wire  _T_12714; // @[package.scala 96:25:@57217.4 package.scala 96:25:@57218.4]
  wire [7:0] _T_12734; // @[Mux.scala 31:69:@57263.4]
  wire  _T_12711; // @[package.scala 96:25:@57209.4 package.scala 96:25:@57210.4]
  wire [7:0] _T_12735; // @[Mux.scala 31:69:@57264.4]
  wire  _T_12708; // @[package.scala 96:25:@57201.4 package.scala 96:25:@57202.4]
  wire [7:0] _T_12736; // @[Mux.scala 31:69:@57265.4]
  wire  _T_12705; // @[package.scala 96:25:@57193.4 package.scala 96:25:@57194.4]
  wire [7:0] _T_12737; // @[Mux.scala 31:69:@57266.4]
  wire  _T_12702; // @[package.scala 96:25:@57185.4 package.scala 96:25:@57186.4]
  wire [7:0] _T_12738; // @[Mux.scala 31:69:@57267.4]
  wire  _T_12699; // @[package.scala 96:25:@57177.4 package.scala 96:25:@57178.4]
  wire [7:0] _T_12739; // @[Mux.scala 31:69:@57268.4]
  wire  _T_12696; // @[package.scala 96:25:@57169.4 package.scala 96:25:@57170.4]
  wire [7:0] _T_12740; // @[Mux.scala 31:69:@57269.4]
  wire  _T_12693; // @[package.scala 96:25:@57161.4 package.scala 96:25:@57162.4]
  wire [7:0] _T_12741; // @[Mux.scala 31:69:@57270.4]
  wire  _T_12690; // @[package.scala 96:25:@57153.4 package.scala 96:25:@57154.4]
  wire [7:0] _T_12742; // @[Mux.scala 31:69:@57271.4]
  wire  _T_12687; // @[package.scala 96:25:@57145.4 package.scala 96:25:@57146.4]
  wire [7:0] _T_12743; // @[Mux.scala 31:69:@57272.4]
  wire  _T_12684; // @[package.scala 96:25:@57137.4 package.scala 96:25:@57138.4]
  wire [7:0] _T_12744; // @[Mux.scala 31:69:@57273.4]
  wire  _T_12681; // @[package.scala 96:25:@57129.4 package.scala 96:25:@57130.4]
  wire [7:0] _T_12745; // @[Mux.scala 31:69:@57274.4]
  wire  _T_12678; // @[package.scala 96:25:@57121.4 package.scala 96:25:@57122.4]
  wire [7:0] _T_12746; // @[Mux.scala 31:69:@57275.4]
  wire  _T_12675; // @[package.scala 96:25:@57113.4 package.scala 96:25:@57114.4]
  wire [7:0] _T_12747; // @[Mux.scala 31:69:@57276.4]
  wire  _T_12672; // @[package.scala 96:25:@57105.4 package.scala 96:25:@57106.4]
  wire  _T_12905; // @[package.scala 96:25:@57489.4 package.scala 96:25:@57490.4]
  wire [7:0] _T_12909; // @[Mux.scala 31:69:@57499.4]
  wire  _T_12902; // @[package.scala 96:25:@57481.4 package.scala 96:25:@57482.4]
  wire [7:0] _T_12910; // @[Mux.scala 31:69:@57500.4]
  wire  _T_12899; // @[package.scala 96:25:@57473.4 package.scala 96:25:@57474.4]
  wire [7:0] _T_12911; // @[Mux.scala 31:69:@57501.4]
  wire  _T_12896; // @[package.scala 96:25:@57465.4 package.scala 96:25:@57466.4]
  wire [7:0] _T_12912; // @[Mux.scala 31:69:@57502.4]
  wire  _T_12893; // @[package.scala 96:25:@57457.4 package.scala 96:25:@57458.4]
  wire [7:0] _T_12913; // @[Mux.scala 31:69:@57503.4]
  wire  _T_12890; // @[package.scala 96:25:@57449.4 package.scala 96:25:@57450.4]
  wire [7:0] _T_12914; // @[Mux.scala 31:69:@57504.4]
  wire  _T_12887; // @[package.scala 96:25:@57441.4 package.scala 96:25:@57442.4]
  wire [7:0] _T_12915; // @[Mux.scala 31:69:@57505.4]
  wire  _T_12884; // @[package.scala 96:25:@57433.4 package.scala 96:25:@57434.4]
  wire [7:0] _T_12916; // @[Mux.scala 31:69:@57506.4]
  wire  _T_12881; // @[package.scala 96:25:@57425.4 package.scala 96:25:@57426.4]
  wire [7:0] _T_12917; // @[Mux.scala 31:69:@57507.4]
  wire  _T_12878; // @[package.scala 96:25:@57417.4 package.scala 96:25:@57418.4]
  wire [7:0] _T_12918; // @[Mux.scala 31:69:@57508.4]
  wire  _T_12875; // @[package.scala 96:25:@57409.4 package.scala 96:25:@57410.4]
  wire [7:0] _T_12919; // @[Mux.scala 31:69:@57509.4]
  wire  _T_12872; // @[package.scala 96:25:@57401.4 package.scala 96:25:@57402.4]
  wire [7:0] _T_12920; // @[Mux.scala 31:69:@57510.4]
  wire  _T_12869; // @[package.scala 96:25:@57393.4 package.scala 96:25:@57394.4]
  wire [7:0] _T_12921; // @[Mux.scala 31:69:@57511.4]
  wire  _T_12866; // @[package.scala 96:25:@57385.4 package.scala 96:25:@57386.4]
  wire [7:0] _T_12922; // @[Mux.scala 31:69:@57512.4]
  wire  _T_12863; // @[package.scala 96:25:@57377.4 package.scala 96:25:@57378.4]
  wire [7:0] _T_12923; // @[Mux.scala 31:69:@57513.4]
  wire  _T_12860; // @[package.scala 96:25:@57369.4 package.scala 96:25:@57370.4]
  wire [7:0] _T_12924; // @[Mux.scala 31:69:@57514.4]
  wire  _T_12857; // @[package.scala 96:25:@57361.4 package.scala 96:25:@57362.4]
  wire [7:0] _T_12925; // @[Mux.scala 31:69:@57515.4]
  wire  _T_12854; // @[package.scala 96:25:@57353.4 package.scala 96:25:@57354.4]
  wire [7:0] _T_12926; // @[Mux.scala 31:69:@57516.4]
  wire  _T_12851; // @[package.scala 96:25:@57345.4 package.scala 96:25:@57346.4]
  wire  _T_13084; // @[package.scala 96:25:@57729.4 package.scala 96:25:@57730.4]
  wire [7:0] _T_13088; // @[Mux.scala 31:69:@57739.4]
  wire  _T_13081; // @[package.scala 96:25:@57721.4 package.scala 96:25:@57722.4]
  wire [7:0] _T_13089; // @[Mux.scala 31:69:@57740.4]
  wire  _T_13078; // @[package.scala 96:25:@57713.4 package.scala 96:25:@57714.4]
  wire [7:0] _T_13090; // @[Mux.scala 31:69:@57741.4]
  wire  _T_13075; // @[package.scala 96:25:@57705.4 package.scala 96:25:@57706.4]
  wire [7:0] _T_13091; // @[Mux.scala 31:69:@57742.4]
  wire  _T_13072; // @[package.scala 96:25:@57697.4 package.scala 96:25:@57698.4]
  wire [7:0] _T_13092; // @[Mux.scala 31:69:@57743.4]
  wire  _T_13069; // @[package.scala 96:25:@57689.4 package.scala 96:25:@57690.4]
  wire [7:0] _T_13093; // @[Mux.scala 31:69:@57744.4]
  wire  _T_13066; // @[package.scala 96:25:@57681.4 package.scala 96:25:@57682.4]
  wire [7:0] _T_13094; // @[Mux.scala 31:69:@57745.4]
  wire  _T_13063; // @[package.scala 96:25:@57673.4 package.scala 96:25:@57674.4]
  wire [7:0] _T_13095; // @[Mux.scala 31:69:@57746.4]
  wire  _T_13060; // @[package.scala 96:25:@57665.4 package.scala 96:25:@57666.4]
  wire [7:0] _T_13096; // @[Mux.scala 31:69:@57747.4]
  wire  _T_13057; // @[package.scala 96:25:@57657.4 package.scala 96:25:@57658.4]
  wire [7:0] _T_13097; // @[Mux.scala 31:69:@57748.4]
  wire  _T_13054; // @[package.scala 96:25:@57649.4 package.scala 96:25:@57650.4]
  wire [7:0] _T_13098; // @[Mux.scala 31:69:@57749.4]
  wire  _T_13051; // @[package.scala 96:25:@57641.4 package.scala 96:25:@57642.4]
  wire [7:0] _T_13099; // @[Mux.scala 31:69:@57750.4]
  wire  _T_13048; // @[package.scala 96:25:@57633.4 package.scala 96:25:@57634.4]
  wire [7:0] _T_13100; // @[Mux.scala 31:69:@57751.4]
  wire  _T_13045; // @[package.scala 96:25:@57625.4 package.scala 96:25:@57626.4]
  wire [7:0] _T_13101; // @[Mux.scala 31:69:@57752.4]
  wire  _T_13042; // @[package.scala 96:25:@57617.4 package.scala 96:25:@57618.4]
  wire [7:0] _T_13102; // @[Mux.scala 31:69:@57753.4]
  wire  _T_13039; // @[package.scala 96:25:@57609.4 package.scala 96:25:@57610.4]
  wire [7:0] _T_13103; // @[Mux.scala 31:69:@57754.4]
  wire  _T_13036; // @[package.scala 96:25:@57601.4 package.scala 96:25:@57602.4]
  wire [7:0] _T_13104; // @[Mux.scala 31:69:@57755.4]
  wire  _T_13033; // @[package.scala 96:25:@57593.4 package.scala 96:25:@57594.4]
  wire [7:0] _T_13105; // @[Mux.scala 31:69:@57756.4]
  wire  _T_13030; // @[package.scala 96:25:@57585.4 package.scala 96:25:@57586.4]
  wire  _T_13263; // @[package.scala 96:25:@57969.4 package.scala 96:25:@57970.4]
  wire [7:0] _T_13267; // @[Mux.scala 31:69:@57979.4]
  wire  _T_13260; // @[package.scala 96:25:@57961.4 package.scala 96:25:@57962.4]
  wire [7:0] _T_13268; // @[Mux.scala 31:69:@57980.4]
  wire  _T_13257; // @[package.scala 96:25:@57953.4 package.scala 96:25:@57954.4]
  wire [7:0] _T_13269; // @[Mux.scala 31:69:@57981.4]
  wire  _T_13254; // @[package.scala 96:25:@57945.4 package.scala 96:25:@57946.4]
  wire [7:0] _T_13270; // @[Mux.scala 31:69:@57982.4]
  wire  _T_13251; // @[package.scala 96:25:@57937.4 package.scala 96:25:@57938.4]
  wire [7:0] _T_13271; // @[Mux.scala 31:69:@57983.4]
  wire  _T_13248; // @[package.scala 96:25:@57929.4 package.scala 96:25:@57930.4]
  wire [7:0] _T_13272; // @[Mux.scala 31:69:@57984.4]
  wire  _T_13245; // @[package.scala 96:25:@57921.4 package.scala 96:25:@57922.4]
  wire [7:0] _T_13273; // @[Mux.scala 31:69:@57985.4]
  wire  _T_13242; // @[package.scala 96:25:@57913.4 package.scala 96:25:@57914.4]
  wire [7:0] _T_13274; // @[Mux.scala 31:69:@57986.4]
  wire  _T_13239; // @[package.scala 96:25:@57905.4 package.scala 96:25:@57906.4]
  wire [7:0] _T_13275; // @[Mux.scala 31:69:@57987.4]
  wire  _T_13236; // @[package.scala 96:25:@57897.4 package.scala 96:25:@57898.4]
  wire [7:0] _T_13276; // @[Mux.scala 31:69:@57988.4]
  wire  _T_13233; // @[package.scala 96:25:@57889.4 package.scala 96:25:@57890.4]
  wire [7:0] _T_13277; // @[Mux.scala 31:69:@57989.4]
  wire  _T_13230; // @[package.scala 96:25:@57881.4 package.scala 96:25:@57882.4]
  wire [7:0] _T_13278; // @[Mux.scala 31:69:@57990.4]
  wire  _T_13227; // @[package.scala 96:25:@57873.4 package.scala 96:25:@57874.4]
  wire [7:0] _T_13279; // @[Mux.scala 31:69:@57991.4]
  wire  _T_13224; // @[package.scala 96:25:@57865.4 package.scala 96:25:@57866.4]
  wire [7:0] _T_13280; // @[Mux.scala 31:69:@57992.4]
  wire  _T_13221; // @[package.scala 96:25:@57857.4 package.scala 96:25:@57858.4]
  wire [7:0] _T_13281; // @[Mux.scala 31:69:@57993.4]
  wire  _T_13218; // @[package.scala 96:25:@57849.4 package.scala 96:25:@57850.4]
  wire [7:0] _T_13282; // @[Mux.scala 31:69:@57994.4]
  wire  _T_13215; // @[package.scala 96:25:@57841.4 package.scala 96:25:@57842.4]
  wire [7:0] _T_13283; // @[Mux.scala 31:69:@57995.4]
  wire  _T_13212; // @[package.scala 96:25:@57833.4 package.scala 96:25:@57834.4]
  wire [7:0] _T_13284; // @[Mux.scala 31:69:@57996.4]
  wire  _T_13209; // @[package.scala 96:25:@57825.4 package.scala 96:25:@57826.4]
  wire  _T_13442; // @[package.scala 96:25:@58209.4 package.scala 96:25:@58210.4]
  wire [7:0] _T_13446; // @[Mux.scala 31:69:@58219.4]
  wire  _T_13439; // @[package.scala 96:25:@58201.4 package.scala 96:25:@58202.4]
  wire [7:0] _T_13447; // @[Mux.scala 31:69:@58220.4]
  wire  _T_13436; // @[package.scala 96:25:@58193.4 package.scala 96:25:@58194.4]
  wire [7:0] _T_13448; // @[Mux.scala 31:69:@58221.4]
  wire  _T_13433; // @[package.scala 96:25:@58185.4 package.scala 96:25:@58186.4]
  wire [7:0] _T_13449; // @[Mux.scala 31:69:@58222.4]
  wire  _T_13430; // @[package.scala 96:25:@58177.4 package.scala 96:25:@58178.4]
  wire [7:0] _T_13450; // @[Mux.scala 31:69:@58223.4]
  wire  _T_13427; // @[package.scala 96:25:@58169.4 package.scala 96:25:@58170.4]
  wire [7:0] _T_13451; // @[Mux.scala 31:69:@58224.4]
  wire  _T_13424; // @[package.scala 96:25:@58161.4 package.scala 96:25:@58162.4]
  wire [7:0] _T_13452; // @[Mux.scala 31:69:@58225.4]
  wire  _T_13421; // @[package.scala 96:25:@58153.4 package.scala 96:25:@58154.4]
  wire [7:0] _T_13453; // @[Mux.scala 31:69:@58226.4]
  wire  _T_13418; // @[package.scala 96:25:@58145.4 package.scala 96:25:@58146.4]
  wire [7:0] _T_13454; // @[Mux.scala 31:69:@58227.4]
  wire  _T_13415; // @[package.scala 96:25:@58137.4 package.scala 96:25:@58138.4]
  wire [7:0] _T_13455; // @[Mux.scala 31:69:@58228.4]
  wire  _T_13412; // @[package.scala 96:25:@58129.4 package.scala 96:25:@58130.4]
  wire [7:0] _T_13456; // @[Mux.scala 31:69:@58229.4]
  wire  _T_13409; // @[package.scala 96:25:@58121.4 package.scala 96:25:@58122.4]
  wire [7:0] _T_13457; // @[Mux.scala 31:69:@58230.4]
  wire  _T_13406; // @[package.scala 96:25:@58113.4 package.scala 96:25:@58114.4]
  wire [7:0] _T_13458; // @[Mux.scala 31:69:@58231.4]
  wire  _T_13403; // @[package.scala 96:25:@58105.4 package.scala 96:25:@58106.4]
  wire [7:0] _T_13459; // @[Mux.scala 31:69:@58232.4]
  wire  _T_13400; // @[package.scala 96:25:@58097.4 package.scala 96:25:@58098.4]
  wire [7:0] _T_13460; // @[Mux.scala 31:69:@58233.4]
  wire  _T_13397; // @[package.scala 96:25:@58089.4 package.scala 96:25:@58090.4]
  wire [7:0] _T_13461; // @[Mux.scala 31:69:@58234.4]
  wire  _T_13394; // @[package.scala 96:25:@58081.4 package.scala 96:25:@58082.4]
  wire [7:0] _T_13462; // @[Mux.scala 31:69:@58235.4]
  wire  _T_13391; // @[package.scala 96:25:@58073.4 package.scala 96:25:@58074.4]
  wire [7:0] _T_13463; // @[Mux.scala 31:69:@58236.4]
  wire  _T_13388; // @[package.scala 96:25:@58065.4 package.scala 96:25:@58066.4]
  wire  _T_13621; // @[package.scala 96:25:@58449.4 package.scala 96:25:@58450.4]
  wire [7:0] _T_13625; // @[Mux.scala 31:69:@58459.4]
  wire  _T_13618; // @[package.scala 96:25:@58441.4 package.scala 96:25:@58442.4]
  wire [7:0] _T_13626; // @[Mux.scala 31:69:@58460.4]
  wire  _T_13615; // @[package.scala 96:25:@58433.4 package.scala 96:25:@58434.4]
  wire [7:0] _T_13627; // @[Mux.scala 31:69:@58461.4]
  wire  _T_13612; // @[package.scala 96:25:@58425.4 package.scala 96:25:@58426.4]
  wire [7:0] _T_13628; // @[Mux.scala 31:69:@58462.4]
  wire  _T_13609; // @[package.scala 96:25:@58417.4 package.scala 96:25:@58418.4]
  wire [7:0] _T_13629; // @[Mux.scala 31:69:@58463.4]
  wire  _T_13606; // @[package.scala 96:25:@58409.4 package.scala 96:25:@58410.4]
  wire [7:0] _T_13630; // @[Mux.scala 31:69:@58464.4]
  wire  _T_13603; // @[package.scala 96:25:@58401.4 package.scala 96:25:@58402.4]
  wire [7:0] _T_13631; // @[Mux.scala 31:69:@58465.4]
  wire  _T_13600; // @[package.scala 96:25:@58393.4 package.scala 96:25:@58394.4]
  wire [7:0] _T_13632; // @[Mux.scala 31:69:@58466.4]
  wire  _T_13597; // @[package.scala 96:25:@58385.4 package.scala 96:25:@58386.4]
  wire [7:0] _T_13633; // @[Mux.scala 31:69:@58467.4]
  wire  _T_13594; // @[package.scala 96:25:@58377.4 package.scala 96:25:@58378.4]
  wire [7:0] _T_13634; // @[Mux.scala 31:69:@58468.4]
  wire  _T_13591; // @[package.scala 96:25:@58369.4 package.scala 96:25:@58370.4]
  wire [7:0] _T_13635; // @[Mux.scala 31:69:@58469.4]
  wire  _T_13588; // @[package.scala 96:25:@58361.4 package.scala 96:25:@58362.4]
  wire [7:0] _T_13636; // @[Mux.scala 31:69:@58470.4]
  wire  _T_13585; // @[package.scala 96:25:@58353.4 package.scala 96:25:@58354.4]
  wire [7:0] _T_13637; // @[Mux.scala 31:69:@58471.4]
  wire  _T_13582; // @[package.scala 96:25:@58345.4 package.scala 96:25:@58346.4]
  wire [7:0] _T_13638; // @[Mux.scala 31:69:@58472.4]
  wire  _T_13579; // @[package.scala 96:25:@58337.4 package.scala 96:25:@58338.4]
  wire [7:0] _T_13639; // @[Mux.scala 31:69:@58473.4]
  wire  _T_13576; // @[package.scala 96:25:@58329.4 package.scala 96:25:@58330.4]
  wire [7:0] _T_13640; // @[Mux.scala 31:69:@58474.4]
  wire  _T_13573; // @[package.scala 96:25:@58321.4 package.scala 96:25:@58322.4]
  wire [7:0] _T_13641; // @[Mux.scala 31:69:@58475.4]
  wire  _T_13570; // @[package.scala 96:25:@58313.4 package.scala 96:25:@58314.4]
  wire [7:0] _T_13642; // @[Mux.scala 31:69:@58476.4]
  wire  _T_13567; // @[package.scala 96:25:@58305.4 package.scala 96:25:@58306.4]
  wire  _T_13800; // @[package.scala 96:25:@58689.4 package.scala 96:25:@58690.4]
  wire [7:0] _T_13804; // @[Mux.scala 31:69:@58699.4]
  wire  _T_13797; // @[package.scala 96:25:@58681.4 package.scala 96:25:@58682.4]
  wire [7:0] _T_13805; // @[Mux.scala 31:69:@58700.4]
  wire  _T_13794; // @[package.scala 96:25:@58673.4 package.scala 96:25:@58674.4]
  wire [7:0] _T_13806; // @[Mux.scala 31:69:@58701.4]
  wire  _T_13791; // @[package.scala 96:25:@58665.4 package.scala 96:25:@58666.4]
  wire [7:0] _T_13807; // @[Mux.scala 31:69:@58702.4]
  wire  _T_13788; // @[package.scala 96:25:@58657.4 package.scala 96:25:@58658.4]
  wire [7:0] _T_13808; // @[Mux.scala 31:69:@58703.4]
  wire  _T_13785; // @[package.scala 96:25:@58649.4 package.scala 96:25:@58650.4]
  wire [7:0] _T_13809; // @[Mux.scala 31:69:@58704.4]
  wire  _T_13782; // @[package.scala 96:25:@58641.4 package.scala 96:25:@58642.4]
  wire [7:0] _T_13810; // @[Mux.scala 31:69:@58705.4]
  wire  _T_13779; // @[package.scala 96:25:@58633.4 package.scala 96:25:@58634.4]
  wire [7:0] _T_13811; // @[Mux.scala 31:69:@58706.4]
  wire  _T_13776; // @[package.scala 96:25:@58625.4 package.scala 96:25:@58626.4]
  wire [7:0] _T_13812; // @[Mux.scala 31:69:@58707.4]
  wire  _T_13773; // @[package.scala 96:25:@58617.4 package.scala 96:25:@58618.4]
  wire [7:0] _T_13813; // @[Mux.scala 31:69:@58708.4]
  wire  _T_13770; // @[package.scala 96:25:@58609.4 package.scala 96:25:@58610.4]
  wire [7:0] _T_13814; // @[Mux.scala 31:69:@58709.4]
  wire  _T_13767; // @[package.scala 96:25:@58601.4 package.scala 96:25:@58602.4]
  wire [7:0] _T_13815; // @[Mux.scala 31:69:@58710.4]
  wire  _T_13764; // @[package.scala 96:25:@58593.4 package.scala 96:25:@58594.4]
  wire [7:0] _T_13816; // @[Mux.scala 31:69:@58711.4]
  wire  _T_13761; // @[package.scala 96:25:@58585.4 package.scala 96:25:@58586.4]
  wire [7:0] _T_13817; // @[Mux.scala 31:69:@58712.4]
  wire  _T_13758; // @[package.scala 96:25:@58577.4 package.scala 96:25:@58578.4]
  wire [7:0] _T_13818; // @[Mux.scala 31:69:@58713.4]
  wire  _T_13755; // @[package.scala 96:25:@58569.4 package.scala 96:25:@58570.4]
  wire [7:0] _T_13819; // @[Mux.scala 31:69:@58714.4]
  wire  _T_13752; // @[package.scala 96:25:@58561.4 package.scala 96:25:@58562.4]
  wire [7:0] _T_13820; // @[Mux.scala 31:69:@58715.4]
  wire  _T_13749; // @[package.scala 96:25:@58553.4 package.scala 96:25:@58554.4]
  wire [7:0] _T_13821; // @[Mux.scala 31:69:@58716.4]
  wire  _T_13746; // @[package.scala 96:25:@58545.4 package.scala 96:25:@58546.4]
  wire  _T_13979; // @[package.scala 96:25:@58929.4 package.scala 96:25:@58930.4]
  wire [7:0] _T_13983; // @[Mux.scala 31:69:@58939.4]
  wire  _T_13976; // @[package.scala 96:25:@58921.4 package.scala 96:25:@58922.4]
  wire [7:0] _T_13984; // @[Mux.scala 31:69:@58940.4]
  wire  _T_13973; // @[package.scala 96:25:@58913.4 package.scala 96:25:@58914.4]
  wire [7:0] _T_13985; // @[Mux.scala 31:69:@58941.4]
  wire  _T_13970; // @[package.scala 96:25:@58905.4 package.scala 96:25:@58906.4]
  wire [7:0] _T_13986; // @[Mux.scala 31:69:@58942.4]
  wire  _T_13967; // @[package.scala 96:25:@58897.4 package.scala 96:25:@58898.4]
  wire [7:0] _T_13987; // @[Mux.scala 31:69:@58943.4]
  wire  _T_13964; // @[package.scala 96:25:@58889.4 package.scala 96:25:@58890.4]
  wire [7:0] _T_13988; // @[Mux.scala 31:69:@58944.4]
  wire  _T_13961; // @[package.scala 96:25:@58881.4 package.scala 96:25:@58882.4]
  wire [7:0] _T_13989; // @[Mux.scala 31:69:@58945.4]
  wire  _T_13958; // @[package.scala 96:25:@58873.4 package.scala 96:25:@58874.4]
  wire [7:0] _T_13990; // @[Mux.scala 31:69:@58946.4]
  wire  _T_13955; // @[package.scala 96:25:@58865.4 package.scala 96:25:@58866.4]
  wire [7:0] _T_13991; // @[Mux.scala 31:69:@58947.4]
  wire  _T_13952; // @[package.scala 96:25:@58857.4 package.scala 96:25:@58858.4]
  wire [7:0] _T_13992; // @[Mux.scala 31:69:@58948.4]
  wire  _T_13949; // @[package.scala 96:25:@58849.4 package.scala 96:25:@58850.4]
  wire [7:0] _T_13993; // @[Mux.scala 31:69:@58949.4]
  wire  _T_13946; // @[package.scala 96:25:@58841.4 package.scala 96:25:@58842.4]
  wire [7:0] _T_13994; // @[Mux.scala 31:69:@58950.4]
  wire  _T_13943; // @[package.scala 96:25:@58833.4 package.scala 96:25:@58834.4]
  wire [7:0] _T_13995; // @[Mux.scala 31:69:@58951.4]
  wire  _T_13940; // @[package.scala 96:25:@58825.4 package.scala 96:25:@58826.4]
  wire [7:0] _T_13996; // @[Mux.scala 31:69:@58952.4]
  wire  _T_13937; // @[package.scala 96:25:@58817.4 package.scala 96:25:@58818.4]
  wire [7:0] _T_13997; // @[Mux.scala 31:69:@58953.4]
  wire  _T_13934; // @[package.scala 96:25:@58809.4 package.scala 96:25:@58810.4]
  wire [7:0] _T_13998; // @[Mux.scala 31:69:@58954.4]
  wire  _T_13931; // @[package.scala 96:25:@58801.4 package.scala 96:25:@58802.4]
  wire [7:0] _T_13999; // @[Mux.scala 31:69:@58955.4]
  wire  _T_13928; // @[package.scala 96:25:@58793.4 package.scala 96:25:@58794.4]
  wire [7:0] _T_14000; // @[Mux.scala 31:69:@58956.4]
  wire  _T_13925; // @[package.scala 96:25:@58785.4 package.scala 96:25:@58786.4]
  wire  _T_14158; // @[package.scala 96:25:@59169.4 package.scala 96:25:@59170.4]
  wire [7:0] _T_14162; // @[Mux.scala 31:69:@59179.4]
  wire  _T_14155; // @[package.scala 96:25:@59161.4 package.scala 96:25:@59162.4]
  wire [7:0] _T_14163; // @[Mux.scala 31:69:@59180.4]
  wire  _T_14152; // @[package.scala 96:25:@59153.4 package.scala 96:25:@59154.4]
  wire [7:0] _T_14164; // @[Mux.scala 31:69:@59181.4]
  wire  _T_14149; // @[package.scala 96:25:@59145.4 package.scala 96:25:@59146.4]
  wire [7:0] _T_14165; // @[Mux.scala 31:69:@59182.4]
  wire  _T_14146; // @[package.scala 96:25:@59137.4 package.scala 96:25:@59138.4]
  wire [7:0] _T_14166; // @[Mux.scala 31:69:@59183.4]
  wire  _T_14143; // @[package.scala 96:25:@59129.4 package.scala 96:25:@59130.4]
  wire [7:0] _T_14167; // @[Mux.scala 31:69:@59184.4]
  wire  _T_14140; // @[package.scala 96:25:@59121.4 package.scala 96:25:@59122.4]
  wire [7:0] _T_14168; // @[Mux.scala 31:69:@59185.4]
  wire  _T_14137; // @[package.scala 96:25:@59113.4 package.scala 96:25:@59114.4]
  wire [7:0] _T_14169; // @[Mux.scala 31:69:@59186.4]
  wire  _T_14134; // @[package.scala 96:25:@59105.4 package.scala 96:25:@59106.4]
  wire [7:0] _T_14170; // @[Mux.scala 31:69:@59187.4]
  wire  _T_14131; // @[package.scala 96:25:@59097.4 package.scala 96:25:@59098.4]
  wire [7:0] _T_14171; // @[Mux.scala 31:69:@59188.4]
  wire  _T_14128; // @[package.scala 96:25:@59089.4 package.scala 96:25:@59090.4]
  wire [7:0] _T_14172; // @[Mux.scala 31:69:@59189.4]
  wire  _T_14125; // @[package.scala 96:25:@59081.4 package.scala 96:25:@59082.4]
  wire [7:0] _T_14173; // @[Mux.scala 31:69:@59190.4]
  wire  _T_14122; // @[package.scala 96:25:@59073.4 package.scala 96:25:@59074.4]
  wire [7:0] _T_14174; // @[Mux.scala 31:69:@59191.4]
  wire  _T_14119; // @[package.scala 96:25:@59065.4 package.scala 96:25:@59066.4]
  wire [7:0] _T_14175; // @[Mux.scala 31:69:@59192.4]
  wire  _T_14116; // @[package.scala 96:25:@59057.4 package.scala 96:25:@59058.4]
  wire [7:0] _T_14176; // @[Mux.scala 31:69:@59193.4]
  wire  _T_14113; // @[package.scala 96:25:@59049.4 package.scala 96:25:@59050.4]
  wire [7:0] _T_14177; // @[Mux.scala 31:69:@59194.4]
  wire  _T_14110; // @[package.scala 96:25:@59041.4 package.scala 96:25:@59042.4]
  wire [7:0] _T_14178; // @[Mux.scala 31:69:@59195.4]
  wire  _T_14107; // @[package.scala 96:25:@59033.4 package.scala 96:25:@59034.4]
  wire [7:0] _T_14179; // @[Mux.scala 31:69:@59196.4]
  wire  _T_14104; // @[package.scala 96:25:@59025.4 package.scala 96:25:@59026.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@44319.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@44335.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@44351.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@44367.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@44383.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@44399.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@44415.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@44431.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@44447.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@44463.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@44479.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@44495.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@44511.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@44527.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@44543.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@44559.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  Mem1D_5 Mem1D_16 ( // @[MemPrimitives.scala 64:21:@44575.4]
    .clock(Mem1D_16_clock),
    .reset(Mem1D_16_reset),
    .io_r_ofs_0(Mem1D_16_io_r_ofs_0),
    .io_r_backpressure(Mem1D_16_io_r_backpressure),
    .io_w_ofs_0(Mem1D_16_io_w_ofs_0),
    .io_w_data_0(Mem1D_16_io_w_data_0),
    .io_w_en_0(Mem1D_16_io_w_en_0),
    .io_output(Mem1D_16_io_output)
  );
  Mem1D_5 Mem1D_17 ( // @[MemPrimitives.scala 64:21:@44591.4]
    .clock(Mem1D_17_clock),
    .reset(Mem1D_17_reset),
    .io_r_ofs_0(Mem1D_17_io_r_ofs_0),
    .io_r_backpressure(Mem1D_17_io_r_backpressure),
    .io_w_ofs_0(Mem1D_17_io_w_ofs_0),
    .io_w_data_0(Mem1D_17_io_w_data_0),
    .io_w_en_0(Mem1D_17_io_w_en_0),
    .io_output(Mem1D_17_io_output)
  );
  Mem1D_5 Mem1D_18 ( // @[MemPrimitives.scala 64:21:@44607.4]
    .clock(Mem1D_18_clock),
    .reset(Mem1D_18_reset),
    .io_r_ofs_0(Mem1D_18_io_r_ofs_0),
    .io_r_backpressure(Mem1D_18_io_r_backpressure),
    .io_w_ofs_0(Mem1D_18_io_w_ofs_0),
    .io_w_data_0(Mem1D_18_io_w_data_0),
    .io_w_en_0(Mem1D_18_io_w_en_0),
    .io_output(Mem1D_18_io_output)
  );
  Mem1D_5 Mem1D_19 ( // @[MemPrimitives.scala 64:21:@44623.4]
    .clock(Mem1D_19_clock),
    .reset(Mem1D_19_reset),
    .io_r_ofs_0(Mem1D_19_io_r_ofs_0),
    .io_r_backpressure(Mem1D_19_io_r_backpressure),
    .io_w_ofs_0(Mem1D_19_io_w_ofs_0),
    .io_w_data_0(Mem1D_19_io_w_data_0),
    .io_w_en_0(Mem1D_19_io_w_en_0),
    .io_output(Mem1D_19_io_output)
  );
  Mem1D_5 Mem1D_20 ( // @[MemPrimitives.scala 64:21:@44639.4]
    .clock(Mem1D_20_clock),
    .reset(Mem1D_20_reset),
    .io_r_ofs_0(Mem1D_20_io_r_ofs_0),
    .io_r_backpressure(Mem1D_20_io_r_backpressure),
    .io_w_ofs_0(Mem1D_20_io_w_ofs_0),
    .io_w_data_0(Mem1D_20_io_w_data_0),
    .io_w_en_0(Mem1D_20_io_w_en_0),
    .io_output(Mem1D_20_io_output)
  );
  Mem1D_5 Mem1D_21 ( // @[MemPrimitives.scala 64:21:@44655.4]
    .clock(Mem1D_21_clock),
    .reset(Mem1D_21_reset),
    .io_r_ofs_0(Mem1D_21_io_r_ofs_0),
    .io_r_backpressure(Mem1D_21_io_r_backpressure),
    .io_w_ofs_0(Mem1D_21_io_w_ofs_0),
    .io_w_data_0(Mem1D_21_io_w_data_0),
    .io_w_en_0(Mem1D_21_io_w_en_0),
    .io_output(Mem1D_21_io_output)
  );
  Mem1D_5 Mem1D_22 ( // @[MemPrimitives.scala 64:21:@44671.4]
    .clock(Mem1D_22_clock),
    .reset(Mem1D_22_reset),
    .io_r_ofs_0(Mem1D_22_io_r_ofs_0),
    .io_r_backpressure(Mem1D_22_io_r_backpressure),
    .io_w_ofs_0(Mem1D_22_io_w_ofs_0),
    .io_w_data_0(Mem1D_22_io_w_data_0),
    .io_w_en_0(Mem1D_22_io_w_en_0),
    .io_output(Mem1D_22_io_output)
  );
  Mem1D_5 Mem1D_23 ( // @[MemPrimitives.scala 64:21:@44687.4]
    .clock(Mem1D_23_clock),
    .reset(Mem1D_23_reset),
    .io_r_ofs_0(Mem1D_23_io_r_ofs_0),
    .io_r_backpressure(Mem1D_23_io_r_backpressure),
    .io_w_ofs_0(Mem1D_23_io_w_ofs_0),
    .io_w_data_0(Mem1D_23_io_w_data_0),
    .io_w_en_0(Mem1D_23_io_w_en_0),
    .io_output(Mem1D_23_io_output)
  );
  Mem1D_5 Mem1D_24 ( // @[MemPrimitives.scala 64:21:@44703.4]
    .clock(Mem1D_24_clock),
    .reset(Mem1D_24_reset),
    .io_r_ofs_0(Mem1D_24_io_r_ofs_0),
    .io_r_backpressure(Mem1D_24_io_r_backpressure),
    .io_w_ofs_0(Mem1D_24_io_w_ofs_0),
    .io_w_data_0(Mem1D_24_io_w_data_0),
    .io_w_en_0(Mem1D_24_io_w_en_0),
    .io_output(Mem1D_24_io_output)
  );
  Mem1D_5 Mem1D_25 ( // @[MemPrimitives.scala 64:21:@44719.4]
    .clock(Mem1D_25_clock),
    .reset(Mem1D_25_reset),
    .io_r_ofs_0(Mem1D_25_io_r_ofs_0),
    .io_r_backpressure(Mem1D_25_io_r_backpressure),
    .io_w_ofs_0(Mem1D_25_io_w_ofs_0),
    .io_w_data_0(Mem1D_25_io_w_data_0),
    .io_w_en_0(Mem1D_25_io_w_en_0),
    .io_output(Mem1D_25_io_output)
  );
  Mem1D_5 Mem1D_26 ( // @[MemPrimitives.scala 64:21:@44735.4]
    .clock(Mem1D_26_clock),
    .reset(Mem1D_26_reset),
    .io_r_ofs_0(Mem1D_26_io_r_ofs_0),
    .io_r_backpressure(Mem1D_26_io_r_backpressure),
    .io_w_ofs_0(Mem1D_26_io_w_ofs_0),
    .io_w_data_0(Mem1D_26_io_w_data_0),
    .io_w_en_0(Mem1D_26_io_w_en_0),
    .io_output(Mem1D_26_io_output)
  );
  Mem1D_5 Mem1D_27 ( // @[MemPrimitives.scala 64:21:@44751.4]
    .clock(Mem1D_27_clock),
    .reset(Mem1D_27_reset),
    .io_r_ofs_0(Mem1D_27_io_r_ofs_0),
    .io_r_backpressure(Mem1D_27_io_r_backpressure),
    .io_w_ofs_0(Mem1D_27_io_w_ofs_0),
    .io_w_data_0(Mem1D_27_io_w_data_0),
    .io_w_en_0(Mem1D_27_io_w_en_0),
    .io_output(Mem1D_27_io_output)
  );
  Mem1D_5 Mem1D_28 ( // @[MemPrimitives.scala 64:21:@44767.4]
    .clock(Mem1D_28_clock),
    .reset(Mem1D_28_reset),
    .io_r_ofs_0(Mem1D_28_io_r_ofs_0),
    .io_r_backpressure(Mem1D_28_io_r_backpressure),
    .io_w_ofs_0(Mem1D_28_io_w_ofs_0),
    .io_w_data_0(Mem1D_28_io_w_data_0),
    .io_w_en_0(Mem1D_28_io_w_en_0),
    .io_output(Mem1D_28_io_output)
  );
  Mem1D_5 Mem1D_29 ( // @[MemPrimitives.scala 64:21:@44783.4]
    .clock(Mem1D_29_clock),
    .reset(Mem1D_29_reset),
    .io_r_ofs_0(Mem1D_29_io_r_ofs_0),
    .io_r_backpressure(Mem1D_29_io_r_backpressure),
    .io_w_ofs_0(Mem1D_29_io_w_ofs_0),
    .io_w_data_0(Mem1D_29_io_w_data_0),
    .io_w_en_0(Mem1D_29_io_w_en_0),
    .io_output(Mem1D_29_io_output)
  );
  Mem1D_5 Mem1D_30 ( // @[MemPrimitives.scala 64:21:@44799.4]
    .clock(Mem1D_30_clock),
    .reset(Mem1D_30_reset),
    .io_r_ofs_0(Mem1D_30_io_r_ofs_0),
    .io_r_backpressure(Mem1D_30_io_r_backpressure),
    .io_w_ofs_0(Mem1D_30_io_w_ofs_0),
    .io_w_data_0(Mem1D_30_io_w_data_0),
    .io_w_en_0(Mem1D_30_io_w_en_0),
    .io_output(Mem1D_30_io_output)
  );
  Mem1D_5 Mem1D_31 ( // @[MemPrimitives.scala 64:21:@44815.4]
    .clock(Mem1D_31_clock),
    .reset(Mem1D_31_reset),
    .io_r_ofs_0(Mem1D_31_io_r_ofs_0),
    .io_r_backpressure(Mem1D_31_io_r_backpressure),
    .io_w_ofs_0(Mem1D_31_io_w_ofs_0),
    .io_w_data_0(Mem1D_31_io_w_data_0),
    .io_w_en_0(Mem1D_31_io_w_en_0),
    .io_output(Mem1D_31_io_output)
  );
  Mem1D_5 Mem1D_32 ( // @[MemPrimitives.scala 64:21:@44831.4]
    .clock(Mem1D_32_clock),
    .reset(Mem1D_32_reset),
    .io_r_ofs_0(Mem1D_32_io_r_ofs_0),
    .io_r_backpressure(Mem1D_32_io_r_backpressure),
    .io_w_ofs_0(Mem1D_32_io_w_ofs_0),
    .io_w_data_0(Mem1D_32_io_w_data_0),
    .io_w_en_0(Mem1D_32_io_w_en_0),
    .io_output(Mem1D_32_io_output)
  );
  Mem1D_5 Mem1D_33 ( // @[MemPrimitives.scala 64:21:@44847.4]
    .clock(Mem1D_33_clock),
    .reset(Mem1D_33_reset),
    .io_r_ofs_0(Mem1D_33_io_r_ofs_0),
    .io_r_backpressure(Mem1D_33_io_r_backpressure),
    .io_w_ofs_0(Mem1D_33_io_w_ofs_0),
    .io_w_data_0(Mem1D_33_io_w_data_0),
    .io_w_en_0(Mem1D_33_io_w_en_0),
    .io_output(Mem1D_33_io_output)
  );
  Mem1D_5 Mem1D_34 ( // @[MemPrimitives.scala 64:21:@44863.4]
    .clock(Mem1D_34_clock),
    .reset(Mem1D_34_reset),
    .io_r_ofs_0(Mem1D_34_io_r_ofs_0),
    .io_r_backpressure(Mem1D_34_io_r_backpressure),
    .io_w_ofs_0(Mem1D_34_io_w_ofs_0),
    .io_w_data_0(Mem1D_34_io_w_data_0),
    .io_w_en_0(Mem1D_34_io_w_en_0),
    .io_output(Mem1D_34_io_output)
  );
  Mem1D_5 Mem1D_35 ( // @[MemPrimitives.scala 64:21:@44879.4]
    .clock(Mem1D_35_clock),
    .reset(Mem1D_35_reset),
    .io_r_ofs_0(Mem1D_35_io_r_ofs_0),
    .io_r_backpressure(Mem1D_35_io_r_backpressure),
    .io_w_ofs_0(Mem1D_35_io_w_ofs_0),
    .io_w_data_0(Mem1D_35_io_w_data_0),
    .io_w_en_0(Mem1D_35_io_w_en_0),
    .io_output(Mem1D_35_io_output)
  );
  Mem1D_5 Mem1D_36 ( // @[MemPrimitives.scala 64:21:@44895.4]
    .clock(Mem1D_36_clock),
    .reset(Mem1D_36_reset),
    .io_r_ofs_0(Mem1D_36_io_r_ofs_0),
    .io_r_backpressure(Mem1D_36_io_r_backpressure),
    .io_w_ofs_0(Mem1D_36_io_w_ofs_0),
    .io_w_data_0(Mem1D_36_io_w_data_0),
    .io_w_en_0(Mem1D_36_io_w_en_0),
    .io_output(Mem1D_36_io_output)
  );
  Mem1D_5 Mem1D_37 ( // @[MemPrimitives.scala 64:21:@44911.4]
    .clock(Mem1D_37_clock),
    .reset(Mem1D_37_reset),
    .io_r_ofs_0(Mem1D_37_io_r_ofs_0),
    .io_r_backpressure(Mem1D_37_io_r_backpressure),
    .io_w_ofs_0(Mem1D_37_io_w_ofs_0),
    .io_w_data_0(Mem1D_37_io_w_data_0),
    .io_w_en_0(Mem1D_37_io_w_en_0),
    .io_output(Mem1D_37_io_output)
  );
  Mem1D_5 Mem1D_38 ( // @[MemPrimitives.scala 64:21:@44927.4]
    .clock(Mem1D_38_clock),
    .reset(Mem1D_38_reset),
    .io_r_ofs_0(Mem1D_38_io_r_ofs_0),
    .io_r_backpressure(Mem1D_38_io_r_backpressure),
    .io_w_ofs_0(Mem1D_38_io_w_ofs_0),
    .io_w_data_0(Mem1D_38_io_w_data_0),
    .io_w_en_0(Mem1D_38_io_w_en_0),
    .io_output(Mem1D_38_io_output)
  );
  Mem1D_5 Mem1D_39 ( // @[MemPrimitives.scala 64:21:@44943.4]
    .clock(Mem1D_39_clock),
    .reset(Mem1D_39_reset),
    .io_r_ofs_0(Mem1D_39_io_r_ofs_0),
    .io_r_backpressure(Mem1D_39_io_r_backpressure),
    .io_w_ofs_0(Mem1D_39_io_w_ofs_0),
    .io_w_data_0(Mem1D_39_io_w_data_0),
    .io_w_en_0(Mem1D_39_io_w_en_0),
    .io_output(Mem1D_39_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 121:29:@46339.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_ins_9(StickySelects_io_ins_9),
    .io_ins_10(StickySelects_io_ins_10),
    .io_ins_11(StickySelects_io_ins_11),
    .io_ins_12(StickySelects_io_ins_12),
    .io_ins_13(StickySelects_io_ins_13),
    .io_ins_14(StickySelects_io_ins_14),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8),
    .io_outs_9(StickySelects_io_outs_9),
    .io_outs_10(StickySelects_io_outs_10),
    .io_outs_11(StickySelects_io_outs_11),
    .io_outs_12(StickySelects_io_outs_12),
    .io_outs_13(StickySelects_io_outs_13),
    .io_outs_14(StickySelects_io_outs_14)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 121:29:@46482.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_ins_9(StickySelects_1_io_ins_9),
    .io_ins_10(StickySelects_1_io_ins_10),
    .io_ins_11(StickySelects_1_io_ins_11),
    .io_ins_12(StickySelects_1_io_ins_12),
    .io_ins_13(StickySelects_1_io_ins_13),
    .io_ins_14(StickySelects_1_io_ins_14),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8),
    .io_outs_9(StickySelects_1_io_outs_9),
    .io_outs_10(StickySelects_1_io_outs_10),
    .io_outs_11(StickySelects_1_io_outs_11),
    .io_outs_12(StickySelects_1_io_outs_12),
    .io_outs_13(StickySelects_1_io_outs_13),
    .io_outs_14(StickySelects_1_io_outs_14)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@46625.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_ins_9(StickySelects_2_io_ins_9),
    .io_ins_10(StickySelects_2_io_ins_10),
    .io_ins_11(StickySelects_2_io_ins_11),
    .io_ins_12(StickySelects_2_io_ins_12),
    .io_ins_13(StickySelects_2_io_ins_13),
    .io_ins_14(StickySelects_2_io_ins_14),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8),
    .io_outs_9(StickySelects_2_io_outs_9),
    .io_outs_10(StickySelects_2_io_outs_10),
    .io_outs_11(StickySelects_2_io_outs_11),
    .io_outs_12(StickySelects_2_io_outs_12),
    .io_outs_13(StickySelects_2_io_outs_13),
    .io_outs_14(StickySelects_2_io_outs_14)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@46768.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_ins_9(StickySelects_3_io_ins_9),
    .io_ins_10(StickySelects_3_io_ins_10),
    .io_ins_11(StickySelects_3_io_ins_11),
    .io_ins_12(StickySelects_3_io_ins_12),
    .io_ins_13(StickySelects_3_io_ins_13),
    .io_ins_14(StickySelects_3_io_ins_14),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8),
    .io_outs_9(StickySelects_3_io_outs_9),
    .io_outs_10(StickySelects_3_io_outs_10),
    .io_outs_11(StickySelects_3_io_outs_11),
    .io_outs_12(StickySelects_3_io_outs_12),
    .io_outs_13(StickySelects_3_io_outs_13),
    .io_outs_14(StickySelects_3_io_outs_14)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 121:29:@46911.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_ins_9(StickySelects_4_io_ins_9),
    .io_ins_10(StickySelects_4_io_ins_10),
    .io_ins_11(StickySelects_4_io_ins_11),
    .io_ins_12(StickySelects_4_io_ins_12),
    .io_ins_13(StickySelects_4_io_ins_13),
    .io_ins_14(StickySelects_4_io_ins_14),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8),
    .io_outs_9(StickySelects_4_io_outs_9),
    .io_outs_10(StickySelects_4_io_outs_10),
    .io_outs_11(StickySelects_4_io_outs_11),
    .io_outs_12(StickySelects_4_io_outs_12),
    .io_outs_13(StickySelects_4_io_outs_13),
    .io_outs_14(StickySelects_4_io_outs_14)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 121:29:@47054.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_ins_9(StickySelects_5_io_ins_9),
    .io_ins_10(StickySelects_5_io_ins_10),
    .io_ins_11(StickySelects_5_io_ins_11),
    .io_ins_12(StickySelects_5_io_ins_12),
    .io_ins_13(StickySelects_5_io_ins_13),
    .io_ins_14(StickySelects_5_io_ins_14),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8),
    .io_outs_9(StickySelects_5_io_outs_9),
    .io_outs_10(StickySelects_5_io_outs_10),
    .io_outs_11(StickySelects_5_io_outs_11),
    .io_outs_12(StickySelects_5_io_outs_12),
    .io_outs_13(StickySelects_5_io_outs_13),
    .io_outs_14(StickySelects_5_io_outs_14)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@47197.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_ins_9(StickySelects_6_io_ins_9),
    .io_ins_10(StickySelects_6_io_ins_10),
    .io_ins_11(StickySelects_6_io_ins_11),
    .io_ins_12(StickySelects_6_io_ins_12),
    .io_ins_13(StickySelects_6_io_ins_13),
    .io_ins_14(StickySelects_6_io_ins_14),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8),
    .io_outs_9(StickySelects_6_io_outs_9),
    .io_outs_10(StickySelects_6_io_outs_10),
    .io_outs_11(StickySelects_6_io_outs_11),
    .io_outs_12(StickySelects_6_io_outs_12),
    .io_outs_13(StickySelects_6_io_outs_13),
    .io_outs_14(StickySelects_6_io_outs_14)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@47340.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_ins_9(StickySelects_7_io_ins_9),
    .io_ins_10(StickySelects_7_io_ins_10),
    .io_ins_11(StickySelects_7_io_ins_11),
    .io_ins_12(StickySelects_7_io_ins_12),
    .io_ins_13(StickySelects_7_io_ins_13),
    .io_ins_14(StickySelects_7_io_ins_14),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8),
    .io_outs_9(StickySelects_7_io_outs_9),
    .io_outs_10(StickySelects_7_io_outs_10),
    .io_outs_11(StickySelects_7_io_outs_11),
    .io_outs_12(StickySelects_7_io_outs_12),
    .io_outs_13(StickySelects_7_io_outs_13),
    .io_outs_14(StickySelects_7_io_outs_14)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 121:29:@47483.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_ins_9(StickySelects_8_io_ins_9),
    .io_ins_10(StickySelects_8_io_ins_10),
    .io_ins_11(StickySelects_8_io_ins_11),
    .io_ins_12(StickySelects_8_io_ins_12),
    .io_ins_13(StickySelects_8_io_ins_13),
    .io_ins_14(StickySelects_8_io_ins_14),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8),
    .io_outs_9(StickySelects_8_io_outs_9),
    .io_outs_10(StickySelects_8_io_outs_10),
    .io_outs_11(StickySelects_8_io_outs_11),
    .io_outs_12(StickySelects_8_io_outs_12),
    .io_outs_13(StickySelects_8_io_outs_13),
    .io_outs_14(StickySelects_8_io_outs_14)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 121:29:@47626.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_ins_9(StickySelects_9_io_ins_9),
    .io_ins_10(StickySelects_9_io_ins_10),
    .io_ins_11(StickySelects_9_io_ins_11),
    .io_ins_12(StickySelects_9_io_ins_12),
    .io_ins_13(StickySelects_9_io_ins_13),
    .io_ins_14(StickySelects_9_io_ins_14),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8),
    .io_outs_9(StickySelects_9_io_outs_9),
    .io_outs_10(StickySelects_9_io_outs_10),
    .io_outs_11(StickySelects_9_io_outs_11),
    .io_outs_12(StickySelects_9_io_outs_12),
    .io_outs_13(StickySelects_9_io_outs_13),
    .io_outs_14(StickySelects_9_io_outs_14)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@47769.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_ins_9(StickySelects_10_io_ins_9),
    .io_ins_10(StickySelects_10_io_ins_10),
    .io_ins_11(StickySelects_10_io_ins_11),
    .io_ins_12(StickySelects_10_io_ins_12),
    .io_ins_13(StickySelects_10_io_ins_13),
    .io_ins_14(StickySelects_10_io_ins_14),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8),
    .io_outs_9(StickySelects_10_io_outs_9),
    .io_outs_10(StickySelects_10_io_outs_10),
    .io_outs_11(StickySelects_10_io_outs_11),
    .io_outs_12(StickySelects_10_io_outs_12),
    .io_outs_13(StickySelects_10_io_outs_13),
    .io_outs_14(StickySelects_10_io_outs_14)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@47912.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_ins_9(StickySelects_11_io_ins_9),
    .io_ins_10(StickySelects_11_io_ins_10),
    .io_ins_11(StickySelects_11_io_ins_11),
    .io_ins_12(StickySelects_11_io_ins_12),
    .io_ins_13(StickySelects_11_io_ins_13),
    .io_ins_14(StickySelects_11_io_ins_14),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8),
    .io_outs_9(StickySelects_11_io_outs_9),
    .io_outs_10(StickySelects_11_io_outs_10),
    .io_outs_11(StickySelects_11_io_outs_11),
    .io_outs_12(StickySelects_11_io_outs_12),
    .io_outs_13(StickySelects_11_io_outs_13),
    .io_outs_14(StickySelects_11_io_outs_14)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 121:29:@48055.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_ins_6(StickySelects_12_io_ins_6),
    .io_ins_7(StickySelects_12_io_ins_7),
    .io_ins_8(StickySelects_12_io_ins_8),
    .io_ins_9(StickySelects_12_io_ins_9),
    .io_ins_10(StickySelects_12_io_ins_10),
    .io_ins_11(StickySelects_12_io_ins_11),
    .io_ins_12(StickySelects_12_io_ins_12),
    .io_ins_13(StickySelects_12_io_ins_13),
    .io_ins_14(StickySelects_12_io_ins_14),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5),
    .io_outs_6(StickySelects_12_io_outs_6),
    .io_outs_7(StickySelects_12_io_outs_7),
    .io_outs_8(StickySelects_12_io_outs_8),
    .io_outs_9(StickySelects_12_io_outs_9),
    .io_outs_10(StickySelects_12_io_outs_10),
    .io_outs_11(StickySelects_12_io_outs_11),
    .io_outs_12(StickySelects_12_io_outs_12),
    .io_outs_13(StickySelects_12_io_outs_13),
    .io_outs_14(StickySelects_12_io_outs_14)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 121:29:@48198.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_ins_6(StickySelects_13_io_ins_6),
    .io_ins_7(StickySelects_13_io_ins_7),
    .io_ins_8(StickySelects_13_io_ins_8),
    .io_ins_9(StickySelects_13_io_ins_9),
    .io_ins_10(StickySelects_13_io_ins_10),
    .io_ins_11(StickySelects_13_io_ins_11),
    .io_ins_12(StickySelects_13_io_ins_12),
    .io_ins_13(StickySelects_13_io_ins_13),
    .io_ins_14(StickySelects_13_io_ins_14),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5),
    .io_outs_6(StickySelects_13_io_outs_6),
    .io_outs_7(StickySelects_13_io_outs_7),
    .io_outs_8(StickySelects_13_io_outs_8),
    .io_outs_9(StickySelects_13_io_outs_9),
    .io_outs_10(StickySelects_13_io_outs_10),
    .io_outs_11(StickySelects_13_io_outs_11),
    .io_outs_12(StickySelects_13_io_outs_12),
    .io_outs_13(StickySelects_13_io_outs_13),
    .io_outs_14(StickySelects_13_io_outs_14)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@48341.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_ins_8(StickySelects_14_io_ins_8),
    .io_ins_9(StickySelects_14_io_ins_9),
    .io_ins_10(StickySelects_14_io_ins_10),
    .io_ins_11(StickySelects_14_io_ins_11),
    .io_ins_12(StickySelects_14_io_ins_12),
    .io_ins_13(StickySelects_14_io_ins_13),
    .io_ins_14(StickySelects_14_io_ins_14),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7),
    .io_outs_8(StickySelects_14_io_outs_8),
    .io_outs_9(StickySelects_14_io_outs_9),
    .io_outs_10(StickySelects_14_io_outs_10),
    .io_outs_11(StickySelects_14_io_outs_11),
    .io_outs_12(StickySelects_14_io_outs_12),
    .io_outs_13(StickySelects_14_io_outs_13),
    .io_outs_14(StickySelects_14_io_outs_14)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@48484.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_ins_8(StickySelects_15_io_ins_8),
    .io_ins_9(StickySelects_15_io_ins_9),
    .io_ins_10(StickySelects_15_io_ins_10),
    .io_ins_11(StickySelects_15_io_ins_11),
    .io_ins_12(StickySelects_15_io_ins_12),
    .io_ins_13(StickySelects_15_io_ins_13),
    .io_ins_14(StickySelects_15_io_ins_14),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7),
    .io_outs_8(StickySelects_15_io_outs_8),
    .io_outs_9(StickySelects_15_io_outs_9),
    .io_outs_10(StickySelects_15_io_outs_10),
    .io_outs_11(StickySelects_15_io_outs_11),
    .io_outs_12(StickySelects_15_io_outs_12),
    .io_outs_13(StickySelects_15_io_outs_13),
    .io_outs_14(StickySelects_15_io_outs_14)
  );
  StickySelects_1 StickySelects_16 ( // @[MemPrimitives.scala 121:29:@48627.4]
    .clock(StickySelects_16_clock),
    .reset(StickySelects_16_reset),
    .io_ins_0(StickySelects_16_io_ins_0),
    .io_ins_1(StickySelects_16_io_ins_1),
    .io_ins_2(StickySelects_16_io_ins_2),
    .io_ins_3(StickySelects_16_io_ins_3),
    .io_ins_4(StickySelects_16_io_ins_4),
    .io_ins_5(StickySelects_16_io_ins_5),
    .io_ins_6(StickySelects_16_io_ins_6),
    .io_ins_7(StickySelects_16_io_ins_7),
    .io_ins_8(StickySelects_16_io_ins_8),
    .io_ins_9(StickySelects_16_io_ins_9),
    .io_ins_10(StickySelects_16_io_ins_10),
    .io_ins_11(StickySelects_16_io_ins_11),
    .io_ins_12(StickySelects_16_io_ins_12),
    .io_ins_13(StickySelects_16_io_ins_13),
    .io_ins_14(StickySelects_16_io_ins_14),
    .io_outs_0(StickySelects_16_io_outs_0),
    .io_outs_1(StickySelects_16_io_outs_1),
    .io_outs_2(StickySelects_16_io_outs_2),
    .io_outs_3(StickySelects_16_io_outs_3),
    .io_outs_4(StickySelects_16_io_outs_4),
    .io_outs_5(StickySelects_16_io_outs_5),
    .io_outs_6(StickySelects_16_io_outs_6),
    .io_outs_7(StickySelects_16_io_outs_7),
    .io_outs_8(StickySelects_16_io_outs_8),
    .io_outs_9(StickySelects_16_io_outs_9),
    .io_outs_10(StickySelects_16_io_outs_10),
    .io_outs_11(StickySelects_16_io_outs_11),
    .io_outs_12(StickySelects_16_io_outs_12),
    .io_outs_13(StickySelects_16_io_outs_13),
    .io_outs_14(StickySelects_16_io_outs_14)
  );
  StickySelects_1 StickySelects_17 ( // @[MemPrimitives.scala 121:29:@48770.4]
    .clock(StickySelects_17_clock),
    .reset(StickySelects_17_reset),
    .io_ins_0(StickySelects_17_io_ins_0),
    .io_ins_1(StickySelects_17_io_ins_1),
    .io_ins_2(StickySelects_17_io_ins_2),
    .io_ins_3(StickySelects_17_io_ins_3),
    .io_ins_4(StickySelects_17_io_ins_4),
    .io_ins_5(StickySelects_17_io_ins_5),
    .io_ins_6(StickySelects_17_io_ins_6),
    .io_ins_7(StickySelects_17_io_ins_7),
    .io_ins_8(StickySelects_17_io_ins_8),
    .io_ins_9(StickySelects_17_io_ins_9),
    .io_ins_10(StickySelects_17_io_ins_10),
    .io_ins_11(StickySelects_17_io_ins_11),
    .io_ins_12(StickySelects_17_io_ins_12),
    .io_ins_13(StickySelects_17_io_ins_13),
    .io_ins_14(StickySelects_17_io_ins_14),
    .io_outs_0(StickySelects_17_io_outs_0),
    .io_outs_1(StickySelects_17_io_outs_1),
    .io_outs_2(StickySelects_17_io_outs_2),
    .io_outs_3(StickySelects_17_io_outs_3),
    .io_outs_4(StickySelects_17_io_outs_4),
    .io_outs_5(StickySelects_17_io_outs_5),
    .io_outs_6(StickySelects_17_io_outs_6),
    .io_outs_7(StickySelects_17_io_outs_7),
    .io_outs_8(StickySelects_17_io_outs_8),
    .io_outs_9(StickySelects_17_io_outs_9),
    .io_outs_10(StickySelects_17_io_outs_10),
    .io_outs_11(StickySelects_17_io_outs_11),
    .io_outs_12(StickySelects_17_io_outs_12),
    .io_outs_13(StickySelects_17_io_outs_13),
    .io_outs_14(StickySelects_17_io_outs_14)
  );
  StickySelects_1 StickySelects_18 ( // @[MemPrimitives.scala 121:29:@48913.4]
    .clock(StickySelects_18_clock),
    .reset(StickySelects_18_reset),
    .io_ins_0(StickySelects_18_io_ins_0),
    .io_ins_1(StickySelects_18_io_ins_1),
    .io_ins_2(StickySelects_18_io_ins_2),
    .io_ins_3(StickySelects_18_io_ins_3),
    .io_ins_4(StickySelects_18_io_ins_4),
    .io_ins_5(StickySelects_18_io_ins_5),
    .io_ins_6(StickySelects_18_io_ins_6),
    .io_ins_7(StickySelects_18_io_ins_7),
    .io_ins_8(StickySelects_18_io_ins_8),
    .io_ins_9(StickySelects_18_io_ins_9),
    .io_ins_10(StickySelects_18_io_ins_10),
    .io_ins_11(StickySelects_18_io_ins_11),
    .io_ins_12(StickySelects_18_io_ins_12),
    .io_ins_13(StickySelects_18_io_ins_13),
    .io_ins_14(StickySelects_18_io_ins_14),
    .io_outs_0(StickySelects_18_io_outs_0),
    .io_outs_1(StickySelects_18_io_outs_1),
    .io_outs_2(StickySelects_18_io_outs_2),
    .io_outs_3(StickySelects_18_io_outs_3),
    .io_outs_4(StickySelects_18_io_outs_4),
    .io_outs_5(StickySelects_18_io_outs_5),
    .io_outs_6(StickySelects_18_io_outs_6),
    .io_outs_7(StickySelects_18_io_outs_7),
    .io_outs_8(StickySelects_18_io_outs_8),
    .io_outs_9(StickySelects_18_io_outs_9),
    .io_outs_10(StickySelects_18_io_outs_10),
    .io_outs_11(StickySelects_18_io_outs_11),
    .io_outs_12(StickySelects_18_io_outs_12),
    .io_outs_13(StickySelects_18_io_outs_13),
    .io_outs_14(StickySelects_18_io_outs_14)
  );
  StickySelects_1 StickySelects_19 ( // @[MemPrimitives.scala 121:29:@49056.4]
    .clock(StickySelects_19_clock),
    .reset(StickySelects_19_reset),
    .io_ins_0(StickySelects_19_io_ins_0),
    .io_ins_1(StickySelects_19_io_ins_1),
    .io_ins_2(StickySelects_19_io_ins_2),
    .io_ins_3(StickySelects_19_io_ins_3),
    .io_ins_4(StickySelects_19_io_ins_4),
    .io_ins_5(StickySelects_19_io_ins_5),
    .io_ins_6(StickySelects_19_io_ins_6),
    .io_ins_7(StickySelects_19_io_ins_7),
    .io_ins_8(StickySelects_19_io_ins_8),
    .io_ins_9(StickySelects_19_io_ins_9),
    .io_ins_10(StickySelects_19_io_ins_10),
    .io_ins_11(StickySelects_19_io_ins_11),
    .io_ins_12(StickySelects_19_io_ins_12),
    .io_ins_13(StickySelects_19_io_ins_13),
    .io_ins_14(StickySelects_19_io_ins_14),
    .io_outs_0(StickySelects_19_io_outs_0),
    .io_outs_1(StickySelects_19_io_outs_1),
    .io_outs_2(StickySelects_19_io_outs_2),
    .io_outs_3(StickySelects_19_io_outs_3),
    .io_outs_4(StickySelects_19_io_outs_4),
    .io_outs_5(StickySelects_19_io_outs_5),
    .io_outs_6(StickySelects_19_io_outs_6),
    .io_outs_7(StickySelects_19_io_outs_7),
    .io_outs_8(StickySelects_19_io_outs_8),
    .io_outs_9(StickySelects_19_io_outs_9),
    .io_outs_10(StickySelects_19_io_outs_10),
    .io_outs_11(StickySelects_19_io_outs_11),
    .io_outs_12(StickySelects_19_io_outs_12),
    .io_outs_13(StickySelects_19_io_outs_13),
    .io_outs_14(StickySelects_19_io_outs_14)
  );
  StickySelects_1 StickySelects_20 ( // @[MemPrimitives.scala 121:29:@49199.4]
    .clock(StickySelects_20_clock),
    .reset(StickySelects_20_reset),
    .io_ins_0(StickySelects_20_io_ins_0),
    .io_ins_1(StickySelects_20_io_ins_1),
    .io_ins_2(StickySelects_20_io_ins_2),
    .io_ins_3(StickySelects_20_io_ins_3),
    .io_ins_4(StickySelects_20_io_ins_4),
    .io_ins_5(StickySelects_20_io_ins_5),
    .io_ins_6(StickySelects_20_io_ins_6),
    .io_ins_7(StickySelects_20_io_ins_7),
    .io_ins_8(StickySelects_20_io_ins_8),
    .io_ins_9(StickySelects_20_io_ins_9),
    .io_ins_10(StickySelects_20_io_ins_10),
    .io_ins_11(StickySelects_20_io_ins_11),
    .io_ins_12(StickySelects_20_io_ins_12),
    .io_ins_13(StickySelects_20_io_ins_13),
    .io_ins_14(StickySelects_20_io_ins_14),
    .io_outs_0(StickySelects_20_io_outs_0),
    .io_outs_1(StickySelects_20_io_outs_1),
    .io_outs_2(StickySelects_20_io_outs_2),
    .io_outs_3(StickySelects_20_io_outs_3),
    .io_outs_4(StickySelects_20_io_outs_4),
    .io_outs_5(StickySelects_20_io_outs_5),
    .io_outs_6(StickySelects_20_io_outs_6),
    .io_outs_7(StickySelects_20_io_outs_7),
    .io_outs_8(StickySelects_20_io_outs_8),
    .io_outs_9(StickySelects_20_io_outs_9),
    .io_outs_10(StickySelects_20_io_outs_10),
    .io_outs_11(StickySelects_20_io_outs_11),
    .io_outs_12(StickySelects_20_io_outs_12),
    .io_outs_13(StickySelects_20_io_outs_13),
    .io_outs_14(StickySelects_20_io_outs_14)
  );
  StickySelects_1 StickySelects_21 ( // @[MemPrimitives.scala 121:29:@49342.4]
    .clock(StickySelects_21_clock),
    .reset(StickySelects_21_reset),
    .io_ins_0(StickySelects_21_io_ins_0),
    .io_ins_1(StickySelects_21_io_ins_1),
    .io_ins_2(StickySelects_21_io_ins_2),
    .io_ins_3(StickySelects_21_io_ins_3),
    .io_ins_4(StickySelects_21_io_ins_4),
    .io_ins_5(StickySelects_21_io_ins_5),
    .io_ins_6(StickySelects_21_io_ins_6),
    .io_ins_7(StickySelects_21_io_ins_7),
    .io_ins_8(StickySelects_21_io_ins_8),
    .io_ins_9(StickySelects_21_io_ins_9),
    .io_ins_10(StickySelects_21_io_ins_10),
    .io_ins_11(StickySelects_21_io_ins_11),
    .io_ins_12(StickySelects_21_io_ins_12),
    .io_ins_13(StickySelects_21_io_ins_13),
    .io_ins_14(StickySelects_21_io_ins_14),
    .io_outs_0(StickySelects_21_io_outs_0),
    .io_outs_1(StickySelects_21_io_outs_1),
    .io_outs_2(StickySelects_21_io_outs_2),
    .io_outs_3(StickySelects_21_io_outs_3),
    .io_outs_4(StickySelects_21_io_outs_4),
    .io_outs_5(StickySelects_21_io_outs_5),
    .io_outs_6(StickySelects_21_io_outs_6),
    .io_outs_7(StickySelects_21_io_outs_7),
    .io_outs_8(StickySelects_21_io_outs_8),
    .io_outs_9(StickySelects_21_io_outs_9),
    .io_outs_10(StickySelects_21_io_outs_10),
    .io_outs_11(StickySelects_21_io_outs_11),
    .io_outs_12(StickySelects_21_io_outs_12),
    .io_outs_13(StickySelects_21_io_outs_13),
    .io_outs_14(StickySelects_21_io_outs_14)
  );
  StickySelects_1 StickySelects_22 ( // @[MemPrimitives.scala 121:29:@49485.4]
    .clock(StickySelects_22_clock),
    .reset(StickySelects_22_reset),
    .io_ins_0(StickySelects_22_io_ins_0),
    .io_ins_1(StickySelects_22_io_ins_1),
    .io_ins_2(StickySelects_22_io_ins_2),
    .io_ins_3(StickySelects_22_io_ins_3),
    .io_ins_4(StickySelects_22_io_ins_4),
    .io_ins_5(StickySelects_22_io_ins_5),
    .io_ins_6(StickySelects_22_io_ins_6),
    .io_ins_7(StickySelects_22_io_ins_7),
    .io_ins_8(StickySelects_22_io_ins_8),
    .io_ins_9(StickySelects_22_io_ins_9),
    .io_ins_10(StickySelects_22_io_ins_10),
    .io_ins_11(StickySelects_22_io_ins_11),
    .io_ins_12(StickySelects_22_io_ins_12),
    .io_ins_13(StickySelects_22_io_ins_13),
    .io_ins_14(StickySelects_22_io_ins_14),
    .io_outs_0(StickySelects_22_io_outs_0),
    .io_outs_1(StickySelects_22_io_outs_1),
    .io_outs_2(StickySelects_22_io_outs_2),
    .io_outs_3(StickySelects_22_io_outs_3),
    .io_outs_4(StickySelects_22_io_outs_4),
    .io_outs_5(StickySelects_22_io_outs_5),
    .io_outs_6(StickySelects_22_io_outs_6),
    .io_outs_7(StickySelects_22_io_outs_7),
    .io_outs_8(StickySelects_22_io_outs_8),
    .io_outs_9(StickySelects_22_io_outs_9),
    .io_outs_10(StickySelects_22_io_outs_10),
    .io_outs_11(StickySelects_22_io_outs_11),
    .io_outs_12(StickySelects_22_io_outs_12),
    .io_outs_13(StickySelects_22_io_outs_13),
    .io_outs_14(StickySelects_22_io_outs_14)
  );
  StickySelects_1 StickySelects_23 ( // @[MemPrimitives.scala 121:29:@49628.4]
    .clock(StickySelects_23_clock),
    .reset(StickySelects_23_reset),
    .io_ins_0(StickySelects_23_io_ins_0),
    .io_ins_1(StickySelects_23_io_ins_1),
    .io_ins_2(StickySelects_23_io_ins_2),
    .io_ins_3(StickySelects_23_io_ins_3),
    .io_ins_4(StickySelects_23_io_ins_4),
    .io_ins_5(StickySelects_23_io_ins_5),
    .io_ins_6(StickySelects_23_io_ins_6),
    .io_ins_7(StickySelects_23_io_ins_7),
    .io_ins_8(StickySelects_23_io_ins_8),
    .io_ins_9(StickySelects_23_io_ins_9),
    .io_ins_10(StickySelects_23_io_ins_10),
    .io_ins_11(StickySelects_23_io_ins_11),
    .io_ins_12(StickySelects_23_io_ins_12),
    .io_ins_13(StickySelects_23_io_ins_13),
    .io_ins_14(StickySelects_23_io_ins_14),
    .io_outs_0(StickySelects_23_io_outs_0),
    .io_outs_1(StickySelects_23_io_outs_1),
    .io_outs_2(StickySelects_23_io_outs_2),
    .io_outs_3(StickySelects_23_io_outs_3),
    .io_outs_4(StickySelects_23_io_outs_4),
    .io_outs_5(StickySelects_23_io_outs_5),
    .io_outs_6(StickySelects_23_io_outs_6),
    .io_outs_7(StickySelects_23_io_outs_7),
    .io_outs_8(StickySelects_23_io_outs_8),
    .io_outs_9(StickySelects_23_io_outs_9),
    .io_outs_10(StickySelects_23_io_outs_10),
    .io_outs_11(StickySelects_23_io_outs_11),
    .io_outs_12(StickySelects_23_io_outs_12),
    .io_outs_13(StickySelects_23_io_outs_13),
    .io_outs_14(StickySelects_23_io_outs_14)
  );
  StickySelects_1 StickySelects_24 ( // @[MemPrimitives.scala 121:29:@49771.4]
    .clock(StickySelects_24_clock),
    .reset(StickySelects_24_reset),
    .io_ins_0(StickySelects_24_io_ins_0),
    .io_ins_1(StickySelects_24_io_ins_1),
    .io_ins_2(StickySelects_24_io_ins_2),
    .io_ins_3(StickySelects_24_io_ins_3),
    .io_ins_4(StickySelects_24_io_ins_4),
    .io_ins_5(StickySelects_24_io_ins_5),
    .io_ins_6(StickySelects_24_io_ins_6),
    .io_ins_7(StickySelects_24_io_ins_7),
    .io_ins_8(StickySelects_24_io_ins_8),
    .io_ins_9(StickySelects_24_io_ins_9),
    .io_ins_10(StickySelects_24_io_ins_10),
    .io_ins_11(StickySelects_24_io_ins_11),
    .io_ins_12(StickySelects_24_io_ins_12),
    .io_ins_13(StickySelects_24_io_ins_13),
    .io_ins_14(StickySelects_24_io_ins_14),
    .io_outs_0(StickySelects_24_io_outs_0),
    .io_outs_1(StickySelects_24_io_outs_1),
    .io_outs_2(StickySelects_24_io_outs_2),
    .io_outs_3(StickySelects_24_io_outs_3),
    .io_outs_4(StickySelects_24_io_outs_4),
    .io_outs_5(StickySelects_24_io_outs_5),
    .io_outs_6(StickySelects_24_io_outs_6),
    .io_outs_7(StickySelects_24_io_outs_7),
    .io_outs_8(StickySelects_24_io_outs_8),
    .io_outs_9(StickySelects_24_io_outs_9),
    .io_outs_10(StickySelects_24_io_outs_10),
    .io_outs_11(StickySelects_24_io_outs_11),
    .io_outs_12(StickySelects_24_io_outs_12),
    .io_outs_13(StickySelects_24_io_outs_13),
    .io_outs_14(StickySelects_24_io_outs_14)
  );
  StickySelects_1 StickySelects_25 ( // @[MemPrimitives.scala 121:29:@49914.4]
    .clock(StickySelects_25_clock),
    .reset(StickySelects_25_reset),
    .io_ins_0(StickySelects_25_io_ins_0),
    .io_ins_1(StickySelects_25_io_ins_1),
    .io_ins_2(StickySelects_25_io_ins_2),
    .io_ins_3(StickySelects_25_io_ins_3),
    .io_ins_4(StickySelects_25_io_ins_4),
    .io_ins_5(StickySelects_25_io_ins_5),
    .io_ins_6(StickySelects_25_io_ins_6),
    .io_ins_7(StickySelects_25_io_ins_7),
    .io_ins_8(StickySelects_25_io_ins_8),
    .io_ins_9(StickySelects_25_io_ins_9),
    .io_ins_10(StickySelects_25_io_ins_10),
    .io_ins_11(StickySelects_25_io_ins_11),
    .io_ins_12(StickySelects_25_io_ins_12),
    .io_ins_13(StickySelects_25_io_ins_13),
    .io_ins_14(StickySelects_25_io_ins_14),
    .io_outs_0(StickySelects_25_io_outs_0),
    .io_outs_1(StickySelects_25_io_outs_1),
    .io_outs_2(StickySelects_25_io_outs_2),
    .io_outs_3(StickySelects_25_io_outs_3),
    .io_outs_4(StickySelects_25_io_outs_4),
    .io_outs_5(StickySelects_25_io_outs_5),
    .io_outs_6(StickySelects_25_io_outs_6),
    .io_outs_7(StickySelects_25_io_outs_7),
    .io_outs_8(StickySelects_25_io_outs_8),
    .io_outs_9(StickySelects_25_io_outs_9),
    .io_outs_10(StickySelects_25_io_outs_10),
    .io_outs_11(StickySelects_25_io_outs_11),
    .io_outs_12(StickySelects_25_io_outs_12),
    .io_outs_13(StickySelects_25_io_outs_13),
    .io_outs_14(StickySelects_25_io_outs_14)
  );
  StickySelects_1 StickySelects_26 ( // @[MemPrimitives.scala 121:29:@50057.4]
    .clock(StickySelects_26_clock),
    .reset(StickySelects_26_reset),
    .io_ins_0(StickySelects_26_io_ins_0),
    .io_ins_1(StickySelects_26_io_ins_1),
    .io_ins_2(StickySelects_26_io_ins_2),
    .io_ins_3(StickySelects_26_io_ins_3),
    .io_ins_4(StickySelects_26_io_ins_4),
    .io_ins_5(StickySelects_26_io_ins_5),
    .io_ins_6(StickySelects_26_io_ins_6),
    .io_ins_7(StickySelects_26_io_ins_7),
    .io_ins_8(StickySelects_26_io_ins_8),
    .io_ins_9(StickySelects_26_io_ins_9),
    .io_ins_10(StickySelects_26_io_ins_10),
    .io_ins_11(StickySelects_26_io_ins_11),
    .io_ins_12(StickySelects_26_io_ins_12),
    .io_ins_13(StickySelects_26_io_ins_13),
    .io_ins_14(StickySelects_26_io_ins_14),
    .io_outs_0(StickySelects_26_io_outs_0),
    .io_outs_1(StickySelects_26_io_outs_1),
    .io_outs_2(StickySelects_26_io_outs_2),
    .io_outs_3(StickySelects_26_io_outs_3),
    .io_outs_4(StickySelects_26_io_outs_4),
    .io_outs_5(StickySelects_26_io_outs_5),
    .io_outs_6(StickySelects_26_io_outs_6),
    .io_outs_7(StickySelects_26_io_outs_7),
    .io_outs_8(StickySelects_26_io_outs_8),
    .io_outs_9(StickySelects_26_io_outs_9),
    .io_outs_10(StickySelects_26_io_outs_10),
    .io_outs_11(StickySelects_26_io_outs_11),
    .io_outs_12(StickySelects_26_io_outs_12),
    .io_outs_13(StickySelects_26_io_outs_13),
    .io_outs_14(StickySelects_26_io_outs_14)
  );
  StickySelects_1 StickySelects_27 ( // @[MemPrimitives.scala 121:29:@50200.4]
    .clock(StickySelects_27_clock),
    .reset(StickySelects_27_reset),
    .io_ins_0(StickySelects_27_io_ins_0),
    .io_ins_1(StickySelects_27_io_ins_1),
    .io_ins_2(StickySelects_27_io_ins_2),
    .io_ins_3(StickySelects_27_io_ins_3),
    .io_ins_4(StickySelects_27_io_ins_4),
    .io_ins_5(StickySelects_27_io_ins_5),
    .io_ins_6(StickySelects_27_io_ins_6),
    .io_ins_7(StickySelects_27_io_ins_7),
    .io_ins_8(StickySelects_27_io_ins_8),
    .io_ins_9(StickySelects_27_io_ins_9),
    .io_ins_10(StickySelects_27_io_ins_10),
    .io_ins_11(StickySelects_27_io_ins_11),
    .io_ins_12(StickySelects_27_io_ins_12),
    .io_ins_13(StickySelects_27_io_ins_13),
    .io_ins_14(StickySelects_27_io_ins_14),
    .io_outs_0(StickySelects_27_io_outs_0),
    .io_outs_1(StickySelects_27_io_outs_1),
    .io_outs_2(StickySelects_27_io_outs_2),
    .io_outs_3(StickySelects_27_io_outs_3),
    .io_outs_4(StickySelects_27_io_outs_4),
    .io_outs_5(StickySelects_27_io_outs_5),
    .io_outs_6(StickySelects_27_io_outs_6),
    .io_outs_7(StickySelects_27_io_outs_7),
    .io_outs_8(StickySelects_27_io_outs_8),
    .io_outs_9(StickySelects_27_io_outs_9),
    .io_outs_10(StickySelects_27_io_outs_10),
    .io_outs_11(StickySelects_27_io_outs_11),
    .io_outs_12(StickySelects_27_io_outs_12),
    .io_outs_13(StickySelects_27_io_outs_13),
    .io_outs_14(StickySelects_27_io_outs_14)
  );
  StickySelects_1 StickySelects_28 ( // @[MemPrimitives.scala 121:29:@50343.4]
    .clock(StickySelects_28_clock),
    .reset(StickySelects_28_reset),
    .io_ins_0(StickySelects_28_io_ins_0),
    .io_ins_1(StickySelects_28_io_ins_1),
    .io_ins_2(StickySelects_28_io_ins_2),
    .io_ins_3(StickySelects_28_io_ins_3),
    .io_ins_4(StickySelects_28_io_ins_4),
    .io_ins_5(StickySelects_28_io_ins_5),
    .io_ins_6(StickySelects_28_io_ins_6),
    .io_ins_7(StickySelects_28_io_ins_7),
    .io_ins_8(StickySelects_28_io_ins_8),
    .io_ins_9(StickySelects_28_io_ins_9),
    .io_ins_10(StickySelects_28_io_ins_10),
    .io_ins_11(StickySelects_28_io_ins_11),
    .io_ins_12(StickySelects_28_io_ins_12),
    .io_ins_13(StickySelects_28_io_ins_13),
    .io_ins_14(StickySelects_28_io_ins_14),
    .io_outs_0(StickySelects_28_io_outs_0),
    .io_outs_1(StickySelects_28_io_outs_1),
    .io_outs_2(StickySelects_28_io_outs_2),
    .io_outs_3(StickySelects_28_io_outs_3),
    .io_outs_4(StickySelects_28_io_outs_4),
    .io_outs_5(StickySelects_28_io_outs_5),
    .io_outs_6(StickySelects_28_io_outs_6),
    .io_outs_7(StickySelects_28_io_outs_7),
    .io_outs_8(StickySelects_28_io_outs_8),
    .io_outs_9(StickySelects_28_io_outs_9),
    .io_outs_10(StickySelects_28_io_outs_10),
    .io_outs_11(StickySelects_28_io_outs_11),
    .io_outs_12(StickySelects_28_io_outs_12),
    .io_outs_13(StickySelects_28_io_outs_13),
    .io_outs_14(StickySelects_28_io_outs_14)
  );
  StickySelects_1 StickySelects_29 ( // @[MemPrimitives.scala 121:29:@50486.4]
    .clock(StickySelects_29_clock),
    .reset(StickySelects_29_reset),
    .io_ins_0(StickySelects_29_io_ins_0),
    .io_ins_1(StickySelects_29_io_ins_1),
    .io_ins_2(StickySelects_29_io_ins_2),
    .io_ins_3(StickySelects_29_io_ins_3),
    .io_ins_4(StickySelects_29_io_ins_4),
    .io_ins_5(StickySelects_29_io_ins_5),
    .io_ins_6(StickySelects_29_io_ins_6),
    .io_ins_7(StickySelects_29_io_ins_7),
    .io_ins_8(StickySelects_29_io_ins_8),
    .io_ins_9(StickySelects_29_io_ins_9),
    .io_ins_10(StickySelects_29_io_ins_10),
    .io_ins_11(StickySelects_29_io_ins_11),
    .io_ins_12(StickySelects_29_io_ins_12),
    .io_ins_13(StickySelects_29_io_ins_13),
    .io_ins_14(StickySelects_29_io_ins_14),
    .io_outs_0(StickySelects_29_io_outs_0),
    .io_outs_1(StickySelects_29_io_outs_1),
    .io_outs_2(StickySelects_29_io_outs_2),
    .io_outs_3(StickySelects_29_io_outs_3),
    .io_outs_4(StickySelects_29_io_outs_4),
    .io_outs_5(StickySelects_29_io_outs_5),
    .io_outs_6(StickySelects_29_io_outs_6),
    .io_outs_7(StickySelects_29_io_outs_7),
    .io_outs_8(StickySelects_29_io_outs_8),
    .io_outs_9(StickySelects_29_io_outs_9),
    .io_outs_10(StickySelects_29_io_outs_10),
    .io_outs_11(StickySelects_29_io_outs_11),
    .io_outs_12(StickySelects_29_io_outs_12),
    .io_outs_13(StickySelects_29_io_outs_13),
    .io_outs_14(StickySelects_29_io_outs_14)
  );
  StickySelects_1 StickySelects_30 ( // @[MemPrimitives.scala 121:29:@50629.4]
    .clock(StickySelects_30_clock),
    .reset(StickySelects_30_reset),
    .io_ins_0(StickySelects_30_io_ins_0),
    .io_ins_1(StickySelects_30_io_ins_1),
    .io_ins_2(StickySelects_30_io_ins_2),
    .io_ins_3(StickySelects_30_io_ins_3),
    .io_ins_4(StickySelects_30_io_ins_4),
    .io_ins_5(StickySelects_30_io_ins_5),
    .io_ins_6(StickySelects_30_io_ins_6),
    .io_ins_7(StickySelects_30_io_ins_7),
    .io_ins_8(StickySelects_30_io_ins_8),
    .io_ins_9(StickySelects_30_io_ins_9),
    .io_ins_10(StickySelects_30_io_ins_10),
    .io_ins_11(StickySelects_30_io_ins_11),
    .io_ins_12(StickySelects_30_io_ins_12),
    .io_ins_13(StickySelects_30_io_ins_13),
    .io_ins_14(StickySelects_30_io_ins_14),
    .io_outs_0(StickySelects_30_io_outs_0),
    .io_outs_1(StickySelects_30_io_outs_1),
    .io_outs_2(StickySelects_30_io_outs_2),
    .io_outs_3(StickySelects_30_io_outs_3),
    .io_outs_4(StickySelects_30_io_outs_4),
    .io_outs_5(StickySelects_30_io_outs_5),
    .io_outs_6(StickySelects_30_io_outs_6),
    .io_outs_7(StickySelects_30_io_outs_7),
    .io_outs_8(StickySelects_30_io_outs_8),
    .io_outs_9(StickySelects_30_io_outs_9),
    .io_outs_10(StickySelects_30_io_outs_10),
    .io_outs_11(StickySelects_30_io_outs_11),
    .io_outs_12(StickySelects_30_io_outs_12),
    .io_outs_13(StickySelects_30_io_outs_13),
    .io_outs_14(StickySelects_30_io_outs_14)
  );
  StickySelects_1 StickySelects_31 ( // @[MemPrimitives.scala 121:29:@50772.4]
    .clock(StickySelects_31_clock),
    .reset(StickySelects_31_reset),
    .io_ins_0(StickySelects_31_io_ins_0),
    .io_ins_1(StickySelects_31_io_ins_1),
    .io_ins_2(StickySelects_31_io_ins_2),
    .io_ins_3(StickySelects_31_io_ins_3),
    .io_ins_4(StickySelects_31_io_ins_4),
    .io_ins_5(StickySelects_31_io_ins_5),
    .io_ins_6(StickySelects_31_io_ins_6),
    .io_ins_7(StickySelects_31_io_ins_7),
    .io_ins_8(StickySelects_31_io_ins_8),
    .io_ins_9(StickySelects_31_io_ins_9),
    .io_ins_10(StickySelects_31_io_ins_10),
    .io_ins_11(StickySelects_31_io_ins_11),
    .io_ins_12(StickySelects_31_io_ins_12),
    .io_ins_13(StickySelects_31_io_ins_13),
    .io_ins_14(StickySelects_31_io_ins_14),
    .io_outs_0(StickySelects_31_io_outs_0),
    .io_outs_1(StickySelects_31_io_outs_1),
    .io_outs_2(StickySelects_31_io_outs_2),
    .io_outs_3(StickySelects_31_io_outs_3),
    .io_outs_4(StickySelects_31_io_outs_4),
    .io_outs_5(StickySelects_31_io_outs_5),
    .io_outs_6(StickySelects_31_io_outs_6),
    .io_outs_7(StickySelects_31_io_outs_7),
    .io_outs_8(StickySelects_31_io_outs_8),
    .io_outs_9(StickySelects_31_io_outs_9),
    .io_outs_10(StickySelects_31_io_outs_10),
    .io_outs_11(StickySelects_31_io_outs_11),
    .io_outs_12(StickySelects_31_io_outs_12),
    .io_outs_13(StickySelects_31_io_outs_13),
    .io_outs_14(StickySelects_31_io_outs_14)
  );
  StickySelects_1 StickySelects_32 ( // @[MemPrimitives.scala 121:29:@50915.4]
    .clock(StickySelects_32_clock),
    .reset(StickySelects_32_reset),
    .io_ins_0(StickySelects_32_io_ins_0),
    .io_ins_1(StickySelects_32_io_ins_1),
    .io_ins_2(StickySelects_32_io_ins_2),
    .io_ins_3(StickySelects_32_io_ins_3),
    .io_ins_4(StickySelects_32_io_ins_4),
    .io_ins_5(StickySelects_32_io_ins_5),
    .io_ins_6(StickySelects_32_io_ins_6),
    .io_ins_7(StickySelects_32_io_ins_7),
    .io_ins_8(StickySelects_32_io_ins_8),
    .io_ins_9(StickySelects_32_io_ins_9),
    .io_ins_10(StickySelects_32_io_ins_10),
    .io_ins_11(StickySelects_32_io_ins_11),
    .io_ins_12(StickySelects_32_io_ins_12),
    .io_ins_13(StickySelects_32_io_ins_13),
    .io_ins_14(StickySelects_32_io_ins_14),
    .io_outs_0(StickySelects_32_io_outs_0),
    .io_outs_1(StickySelects_32_io_outs_1),
    .io_outs_2(StickySelects_32_io_outs_2),
    .io_outs_3(StickySelects_32_io_outs_3),
    .io_outs_4(StickySelects_32_io_outs_4),
    .io_outs_5(StickySelects_32_io_outs_5),
    .io_outs_6(StickySelects_32_io_outs_6),
    .io_outs_7(StickySelects_32_io_outs_7),
    .io_outs_8(StickySelects_32_io_outs_8),
    .io_outs_9(StickySelects_32_io_outs_9),
    .io_outs_10(StickySelects_32_io_outs_10),
    .io_outs_11(StickySelects_32_io_outs_11),
    .io_outs_12(StickySelects_32_io_outs_12),
    .io_outs_13(StickySelects_32_io_outs_13),
    .io_outs_14(StickySelects_32_io_outs_14)
  );
  StickySelects_1 StickySelects_33 ( // @[MemPrimitives.scala 121:29:@51058.4]
    .clock(StickySelects_33_clock),
    .reset(StickySelects_33_reset),
    .io_ins_0(StickySelects_33_io_ins_0),
    .io_ins_1(StickySelects_33_io_ins_1),
    .io_ins_2(StickySelects_33_io_ins_2),
    .io_ins_3(StickySelects_33_io_ins_3),
    .io_ins_4(StickySelects_33_io_ins_4),
    .io_ins_5(StickySelects_33_io_ins_5),
    .io_ins_6(StickySelects_33_io_ins_6),
    .io_ins_7(StickySelects_33_io_ins_7),
    .io_ins_8(StickySelects_33_io_ins_8),
    .io_ins_9(StickySelects_33_io_ins_9),
    .io_ins_10(StickySelects_33_io_ins_10),
    .io_ins_11(StickySelects_33_io_ins_11),
    .io_ins_12(StickySelects_33_io_ins_12),
    .io_ins_13(StickySelects_33_io_ins_13),
    .io_ins_14(StickySelects_33_io_ins_14),
    .io_outs_0(StickySelects_33_io_outs_0),
    .io_outs_1(StickySelects_33_io_outs_1),
    .io_outs_2(StickySelects_33_io_outs_2),
    .io_outs_3(StickySelects_33_io_outs_3),
    .io_outs_4(StickySelects_33_io_outs_4),
    .io_outs_5(StickySelects_33_io_outs_5),
    .io_outs_6(StickySelects_33_io_outs_6),
    .io_outs_7(StickySelects_33_io_outs_7),
    .io_outs_8(StickySelects_33_io_outs_8),
    .io_outs_9(StickySelects_33_io_outs_9),
    .io_outs_10(StickySelects_33_io_outs_10),
    .io_outs_11(StickySelects_33_io_outs_11),
    .io_outs_12(StickySelects_33_io_outs_12),
    .io_outs_13(StickySelects_33_io_outs_13),
    .io_outs_14(StickySelects_33_io_outs_14)
  );
  StickySelects_1 StickySelects_34 ( // @[MemPrimitives.scala 121:29:@51201.4]
    .clock(StickySelects_34_clock),
    .reset(StickySelects_34_reset),
    .io_ins_0(StickySelects_34_io_ins_0),
    .io_ins_1(StickySelects_34_io_ins_1),
    .io_ins_2(StickySelects_34_io_ins_2),
    .io_ins_3(StickySelects_34_io_ins_3),
    .io_ins_4(StickySelects_34_io_ins_4),
    .io_ins_5(StickySelects_34_io_ins_5),
    .io_ins_6(StickySelects_34_io_ins_6),
    .io_ins_7(StickySelects_34_io_ins_7),
    .io_ins_8(StickySelects_34_io_ins_8),
    .io_ins_9(StickySelects_34_io_ins_9),
    .io_ins_10(StickySelects_34_io_ins_10),
    .io_ins_11(StickySelects_34_io_ins_11),
    .io_ins_12(StickySelects_34_io_ins_12),
    .io_ins_13(StickySelects_34_io_ins_13),
    .io_ins_14(StickySelects_34_io_ins_14),
    .io_outs_0(StickySelects_34_io_outs_0),
    .io_outs_1(StickySelects_34_io_outs_1),
    .io_outs_2(StickySelects_34_io_outs_2),
    .io_outs_3(StickySelects_34_io_outs_3),
    .io_outs_4(StickySelects_34_io_outs_4),
    .io_outs_5(StickySelects_34_io_outs_5),
    .io_outs_6(StickySelects_34_io_outs_6),
    .io_outs_7(StickySelects_34_io_outs_7),
    .io_outs_8(StickySelects_34_io_outs_8),
    .io_outs_9(StickySelects_34_io_outs_9),
    .io_outs_10(StickySelects_34_io_outs_10),
    .io_outs_11(StickySelects_34_io_outs_11),
    .io_outs_12(StickySelects_34_io_outs_12),
    .io_outs_13(StickySelects_34_io_outs_13),
    .io_outs_14(StickySelects_34_io_outs_14)
  );
  StickySelects_1 StickySelects_35 ( // @[MemPrimitives.scala 121:29:@51344.4]
    .clock(StickySelects_35_clock),
    .reset(StickySelects_35_reset),
    .io_ins_0(StickySelects_35_io_ins_0),
    .io_ins_1(StickySelects_35_io_ins_1),
    .io_ins_2(StickySelects_35_io_ins_2),
    .io_ins_3(StickySelects_35_io_ins_3),
    .io_ins_4(StickySelects_35_io_ins_4),
    .io_ins_5(StickySelects_35_io_ins_5),
    .io_ins_6(StickySelects_35_io_ins_6),
    .io_ins_7(StickySelects_35_io_ins_7),
    .io_ins_8(StickySelects_35_io_ins_8),
    .io_ins_9(StickySelects_35_io_ins_9),
    .io_ins_10(StickySelects_35_io_ins_10),
    .io_ins_11(StickySelects_35_io_ins_11),
    .io_ins_12(StickySelects_35_io_ins_12),
    .io_ins_13(StickySelects_35_io_ins_13),
    .io_ins_14(StickySelects_35_io_ins_14),
    .io_outs_0(StickySelects_35_io_outs_0),
    .io_outs_1(StickySelects_35_io_outs_1),
    .io_outs_2(StickySelects_35_io_outs_2),
    .io_outs_3(StickySelects_35_io_outs_3),
    .io_outs_4(StickySelects_35_io_outs_4),
    .io_outs_5(StickySelects_35_io_outs_5),
    .io_outs_6(StickySelects_35_io_outs_6),
    .io_outs_7(StickySelects_35_io_outs_7),
    .io_outs_8(StickySelects_35_io_outs_8),
    .io_outs_9(StickySelects_35_io_outs_9),
    .io_outs_10(StickySelects_35_io_outs_10),
    .io_outs_11(StickySelects_35_io_outs_11),
    .io_outs_12(StickySelects_35_io_outs_12),
    .io_outs_13(StickySelects_35_io_outs_13),
    .io_outs_14(StickySelects_35_io_outs_14)
  );
  StickySelects_1 StickySelects_36 ( // @[MemPrimitives.scala 121:29:@51487.4]
    .clock(StickySelects_36_clock),
    .reset(StickySelects_36_reset),
    .io_ins_0(StickySelects_36_io_ins_0),
    .io_ins_1(StickySelects_36_io_ins_1),
    .io_ins_2(StickySelects_36_io_ins_2),
    .io_ins_3(StickySelects_36_io_ins_3),
    .io_ins_4(StickySelects_36_io_ins_4),
    .io_ins_5(StickySelects_36_io_ins_5),
    .io_ins_6(StickySelects_36_io_ins_6),
    .io_ins_7(StickySelects_36_io_ins_7),
    .io_ins_8(StickySelects_36_io_ins_8),
    .io_ins_9(StickySelects_36_io_ins_9),
    .io_ins_10(StickySelects_36_io_ins_10),
    .io_ins_11(StickySelects_36_io_ins_11),
    .io_ins_12(StickySelects_36_io_ins_12),
    .io_ins_13(StickySelects_36_io_ins_13),
    .io_ins_14(StickySelects_36_io_ins_14),
    .io_outs_0(StickySelects_36_io_outs_0),
    .io_outs_1(StickySelects_36_io_outs_1),
    .io_outs_2(StickySelects_36_io_outs_2),
    .io_outs_3(StickySelects_36_io_outs_3),
    .io_outs_4(StickySelects_36_io_outs_4),
    .io_outs_5(StickySelects_36_io_outs_5),
    .io_outs_6(StickySelects_36_io_outs_6),
    .io_outs_7(StickySelects_36_io_outs_7),
    .io_outs_8(StickySelects_36_io_outs_8),
    .io_outs_9(StickySelects_36_io_outs_9),
    .io_outs_10(StickySelects_36_io_outs_10),
    .io_outs_11(StickySelects_36_io_outs_11),
    .io_outs_12(StickySelects_36_io_outs_12),
    .io_outs_13(StickySelects_36_io_outs_13),
    .io_outs_14(StickySelects_36_io_outs_14)
  );
  StickySelects_1 StickySelects_37 ( // @[MemPrimitives.scala 121:29:@51630.4]
    .clock(StickySelects_37_clock),
    .reset(StickySelects_37_reset),
    .io_ins_0(StickySelects_37_io_ins_0),
    .io_ins_1(StickySelects_37_io_ins_1),
    .io_ins_2(StickySelects_37_io_ins_2),
    .io_ins_3(StickySelects_37_io_ins_3),
    .io_ins_4(StickySelects_37_io_ins_4),
    .io_ins_5(StickySelects_37_io_ins_5),
    .io_ins_6(StickySelects_37_io_ins_6),
    .io_ins_7(StickySelects_37_io_ins_7),
    .io_ins_8(StickySelects_37_io_ins_8),
    .io_ins_9(StickySelects_37_io_ins_9),
    .io_ins_10(StickySelects_37_io_ins_10),
    .io_ins_11(StickySelects_37_io_ins_11),
    .io_ins_12(StickySelects_37_io_ins_12),
    .io_ins_13(StickySelects_37_io_ins_13),
    .io_ins_14(StickySelects_37_io_ins_14),
    .io_outs_0(StickySelects_37_io_outs_0),
    .io_outs_1(StickySelects_37_io_outs_1),
    .io_outs_2(StickySelects_37_io_outs_2),
    .io_outs_3(StickySelects_37_io_outs_3),
    .io_outs_4(StickySelects_37_io_outs_4),
    .io_outs_5(StickySelects_37_io_outs_5),
    .io_outs_6(StickySelects_37_io_outs_6),
    .io_outs_7(StickySelects_37_io_outs_7),
    .io_outs_8(StickySelects_37_io_outs_8),
    .io_outs_9(StickySelects_37_io_outs_9),
    .io_outs_10(StickySelects_37_io_outs_10),
    .io_outs_11(StickySelects_37_io_outs_11),
    .io_outs_12(StickySelects_37_io_outs_12),
    .io_outs_13(StickySelects_37_io_outs_13),
    .io_outs_14(StickySelects_37_io_outs_14)
  );
  StickySelects_1 StickySelects_38 ( // @[MemPrimitives.scala 121:29:@51773.4]
    .clock(StickySelects_38_clock),
    .reset(StickySelects_38_reset),
    .io_ins_0(StickySelects_38_io_ins_0),
    .io_ins_1(StickySelects_38_io_ins_1),
    .io_ins_2(StickySelects_38_io_ins_2),
    .io_ins_3(StickySelects_38_io_ins_3),
    .io_ins_4(StickySelects_38_io_ins_4),
    .io_ins_5(StickySelects_38_io_ins_5),
    .io_ins_6(StickySelects_38_io_ins_6),
    .io_ins_7(StickySelects_38_io_ins_7),
    .io_ins_8(StickySelects_38_io_ins_8),
    .io_ins_9(StickySelects_38_io_ins_9),
    .io_ins_10(StickySelects_38_io_ins_10),
    .io_ins_11(StickySelects_38_io_ins_11),
    .io_ins_12(StickySelects_38_io_ins_12),
    .io_ins_13(StickySelects_38_io_ins_13),
    .io_ins_14(StickySelects_38_io_ins_14),
    .io_outs_0(StickySelects_38_io_outs_0),
    .io_outs_1(StickySelects_38_io_outs_1),
    .io_outs_2(StickySelects_38_io_outs_2),
    .io_outs_3(StickySelects_38_io_outs_3),
    .io_outs_4(StickySelects_38_io_outs_4),
    .io_outs_5(StickySelects_38_io_outs_5),
    .io_outs_6(StickySelects_38_io_outs_6),
    .io_outs_7(StickySelects_38_io_outs_7),
    .io_outs_8(StickySelects_38_io_outs_8),
    .io_outs_9(StickySelects_38_io_outs_9),
    .io_outs_10(StickySelects_38_io_outs_10),
    .io_outs_11(StickySelects_38_io_outs_11),
    .io_outs_12(StickySelects_38_io_outs_12),
    .io_outs_13(StickySelects_38_io_outs_13),
    .io_outs_14(StickySelects_38_io_outs_14)
  );
  StickySelects_1 StickySelects_39 ( // @[MemPrimitives.scala 121:29:@51916.4]
    .clock(StickySelects_39_clock),
    .reset(StickySelects_39_reset),
    .io_ins_0(StickySelects_39_io_ins_0),
    .io_ins_1(StickySelects_39_io_ins_1),
    .io_ins_2(StickySelects_39_io_ins_2),
    .io_ins_3(StickySelects_39_io_ins_3),
    .io_ins_4(StickySelects_39_io_ins_4),
    .io_ins_5(StickySelects_39_io_ins_5),
    .io_ins_6(StickySelects_39_io_ins_6),
    .io_ins_7(StickySelects_39_io_ins_7),
    .io_ins_8(StickySelects_39_io_ins_8),
    .io_ins_9(StickySelects_39_io_ins_9),
    .io_ins_10(StickySelects_39_io_ins_10),
    .io_ins_11(StickySelects_39_io_ins_11),
    .io_ins_12(StickySelects_39_io_ins_12),
    .io_ins_13(StickySelects_39_io_ins_13),
    .io_ins_14(StickySelects_39_io_ins_14),
    .io_outs_0(StickySelects_39_io_outs_0),
    .io_outs_1(StickySelects_39_io_outs_1),
    .io_outs_2(StickySelects_39_io_outs_2),
    .io_outs_3(StickySelects_39_io_outs_3),
    .io_outs_4(StickySelects_39_io_outs_4),
    .io_outs_5(StickySelects_39_io_outs_5),
    .io_outs_6(StickySelects_39_io_outs_6),
    .io_outs_7(StickySelects_39_io_outs_7),
    .io_outs_8(StickySelects_39_io_outs_8),
    .io_outs_9(StickySelects_39_io_outs_9),
    .io_outs_10(StickySelects_39_io_outs_10),
    .io_outs_11(StickySelects_39_io_outs_11),
    .io_outs_12(StickySelects_39_io_outs_12),
    .io_outs_13(StickySelects_39_io_outs_13),
    .io_outs_14(StickySelects_39_io_outs_14)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@52060.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@52068.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@52076.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@52084.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@52092.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@52100.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@52108.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@52116.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@52124.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@52132.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@52140.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@52148.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@52156.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@52164.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@52172.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@52180.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@52188.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@52196.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@52204.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@52212.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@52300.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@52308.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@52316.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@52324.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@52332.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@52340.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@52348.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@52356.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@52364.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@52372.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@52380.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@52388.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@52396.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@52404.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@52412.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@52420.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@52428.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@52436.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@52444.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@52452.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@52540.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@52548.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@52556.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@52564.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@52572.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@52580.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@52588.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@52596.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@52604.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@52612.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@52620.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@52628.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@52636.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@52644.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@52652.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@52660.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@52668.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@52676.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@52684.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@52692.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@52780.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@52788.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@52796.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@52804.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@52812.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@52820.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@52828.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@52836.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@52844.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@52852.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@52860.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@52868.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@52876.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@52884.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@52892.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@52900.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@52908.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@52916.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@52924.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@52932.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@53020.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@53028.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@53036.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@53044.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@53052.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@53060.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@53068.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@53076.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@53084.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@53092.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@53100.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@53108.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@53116.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@53124.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@53132.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@53140.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@53148.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@53156.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@53164.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@53172.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@53260.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@53268.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@53276.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@53284.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@53292.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@53300.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@53308.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@53316.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_108 ( // @[package.scala 93:22:@53324.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_109 ( // @[package.scala 93:22:@53332.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_110 ( // @[package.scala 93:22:@53340.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_111 ( // @[package.scala 93:22:@53348.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_112 ( // @[package.scala 93:22:@53356.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_113 ( // @[package.scala 93:22:@53364.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_114 ( // @[package.scala 93:22:@53372.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_115 ( // @[package.scala 93:22:@53380.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_116 ( // @[package.scala 93:22:@53388.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_117 ( // @[package.scala 93:22:@53396.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_118 ( // @[package.scala 93:22:@53404.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_119 ( // @[package.scala 93:22:@53412.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_120 ( // @[package.scala 93:22:@53500.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_121 ( // @[package.scala 93:22:@53508.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_122 ( // @[package.scala 93:22:@53516.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_123 ( // @[package.scala 93:22:@53524.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_124 ( // @[package.scala 93:22:@53532.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_125 ( // @[package.scala 93:22:@53540.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_126 ( // @[package.scala 93:22:@53548.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_127 ( // @[package.scala 93:22:@53556.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_128 ( // @[package.scala 93:22:@53564.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_129 ( // @[package.scala 93:22:@53572.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_130 ( // @[package.scala 93:22:@53580.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_131 ( // @[package.scala 93:22:@53588.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_132 ( // @[package.scala 93:22:@53596.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_133 ( // @[package.scala 93:22:@53604.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_134 ( // @[package.scala 93:22:@53612.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_135 ( // @[package.scala 93:22:@53620.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_136 ( // @[package.scala 93:22:@53628.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_137 ( // @[package.scala 93:22:@53636.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_138 ( // @[package.scala 93:22:@53644.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_139 ( // @[package.scala 93:22:@53652.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_140 ( // @[package.scala 93:22:@53740.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_141 ( // @[package.scala 93:22:@53748.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_142 ( // @[package.scala 93:22:@53756.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_143 ( // @[package.scala 93:22:@53764.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_144 ( // @[package.scala 93:22:@53772.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_145 ( // @[package.scala 93:22:@53780.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_146 ( // @[package.scala 93:22:@53788.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_147 ( // @[package.scala 93:22:@53796.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_148 ( // @[package.scala 93:22:@53804.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_149 ( // @[package.scala 93:22:@53812.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_150 ( // @[package.scala 93:22:@53820.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_151 ( // @[package.scala 93:22:@53828.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_152 ( // @[package.scala 93:22:@53836.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_153 ( // @[package.scala 93:22:@53844.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_154 ( // @[package.scala 93:22:@53852.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_155 ( // @[package.scala 93:22:@53860.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_156 ( // @[package.scala 93:22:@53868.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_157 ( // @[package.scala 93:22:@53876.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_158 ( // @[package.scala 93:22:@53884.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_159 ( // @[package.scala 93:22:@53892.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_160 ( // @[package.scala 93:22:@53980.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_161 ( // @[package.scala 93:22:@53988.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_162 ( // @[package.scala 93:22:@53996.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_163 ( // @[package.scala 93:22:@54004.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_164 ( // @[package.scala 93:22:@54012.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_165 ( // @[package.scala 93:22:@54020.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_166 ( // @[package.scala 93:22:@54028.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_167 ( // @[package.scala 93:22:@54036.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_168 ( // @[package.scala 93:22:@54044.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_169 ( // @[package.scala 93:22:@54052.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_170 ( // @[package.scala 93:22:@54060.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_171 ( // @[package.scala 93:22:@54068.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_172 ( // @[package.scala 93:22:@54076.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_173 ( // @[package.scala 93:22:@54084.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_174 ( // @[package.scala 93:22:@54092.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_175 ( // @[package.scala 93:22:@54100.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_176 ( // @[package.scala 93:22:@54108.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_177 ( // @[package.scala 93:22:@54116.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_178 ( // @[package.scala 93:22:@54124.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_179 ( // @[package.scala 93:22:@54132.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_180 ( // @[package.scala 93:22:@54220.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_181 ( // @[package.scala 93:22:@54228.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_182 ( // @[package.scala 93:22:@54236.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_183 ( // @[package.scala 93:22:@54244.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_184 ( // @[package.scala 93:22:@54252.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_185 ( // @[package.scala 93:22:@54260.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_186 ( // @[package.scala 93:22:@54268.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_187 ( // @[package.scala 93:22:@54276.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_188 ( // @[package.scala 93:22:@54284.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_189 ( // @[package.scala 93:22:@54292.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_190 ( // @[package.scala 93:22:@54300.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_191 ( // @[package.scala 93:22:@54308.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_192 ( // @[package.scala 93:22:@54316.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_193 ( // @[package.scala 93:22:@54324.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_194 ( // @[package.scala 93:22:@54332.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_195 ( // @[package.scala 93:22:@54340.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_196 ( // @[package.scala 93:22:@54348.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_197 ( // @[package.scala 93:22:@54356.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_198 ( // @[package.scala 93:22:@54364.4]
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_199 ( // @[package.scala 93:22:@54372.4]
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_200 ( // @[package.scala 93:22:@54460.4]
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_201 ( // @[package.scala 93:22:@54468.4]
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_202 ( // @[package.scala 93:22:@54476.4]
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_203 ( // @[package.scala 93:22:@54484.4]
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_204 ( // @[package.scala 93:22:@54492.4]
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_205 ( // @[package.scala 93:22:@54500.4]
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_206 ( // @[package.scala 93:22:@54508.4]
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_207 ( // @[package.scala 93:22:@54516.4]
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_208 ( // @[package.scala 93:22:@54524.4]
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_209 ( // @[package.scala 93:22:@54532.4]
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_210 ( // @[package.scala 93:22:@54540.4]
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_211 ( // @[package.scala 93:22:@54548.4]
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_212 ( // @[package.scala 93:22:@54556.4]
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_213 ( // @[package.scala 93:22:@54564.4]
    .clock(RetimeWrapper_213_clock),
    .reset(RetimeWrapper_213_reset),
    .io_flow(RetimeWrapper_213_io_flow),
    .io_in(RetimeWrapper_213_io_in),
    .io_out(RetimeWrapper_213_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_214 ( // @[package.scala 93:22:@54572.4]
    .clock(RetimeWrapper_214_clock),
    .reset(RetimeWrapper_214_reset),
    .io_flow(RetimeWrapper_214_io_flow),
    .io_in(RetimeWrapper_214_io_in),
    .io_out(RetimeWrapper_214_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_215 ( // @[package.scala 93:22:@54580.4]
    .clock(RetimeWrapper_215_clock),
    .reset(RetimeWrapper_215_reset),
    .io_flow(RetimeWrapper_215_io_flow),
    .io_in(RetimeWrapper_215_io_in),
    .io_out(RetimeWrapper_215_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_216 ( // @[package.scala 93:22:@54588.4]
    .clock(RetimeWrapper_216_clock),
    .reset(RetimeWrapper_216_reset),
    .io_flow(RetimeWrapper_216_io_flow),
    .io_in(RetimeWrapper_216_io_in),
    .io_out(RetimeWrapper_216_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_217 ( // @[package.scala 93:22:@54596.4]
    .clock(RetimeWrapper_217_clock),
    .reset(RetimeWrapper_217_reset),
    .io_flow(RetimeWrapper_217_io_flow),
    .io_in(RetimeWrapper_217_io_in),
    .io_out(RetimeWrapper_217_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_218 ( // @[package.scala 93:22:@54604.4]
    .clock(RetimeWrapper_218_clock),
    .reset(RetimeWrapper_218_reset),
    .io_flow(RetimeWrapper_218_io_flow),
    .io_in(RetimeWrapper_218_io_in),
    .io_out(RetimeWrapper_218_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_219 ( // @[package.scala 93:22:@54612.4]
    .clock(RetimeWrapper_219_clock),
    .reset(RetimeWrapper_219_reset),
    .io_flow(RetimeWrapper_219_io_flow),
    .io_in(RetimeWrapper_219_io_in),
    .io_out(RetimeWrapper_219_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_220 ( // @[package.scala 93:22:@54700.4]
    .clock(RetimeWrapper_220_clock),
    .reset(RetimeWrapper_220_reset),
    .io_flow(RetimeWrapper_220_io_flow),
    .io_in(RetimeWrapper_220_io_in),
    .io_out(RetimeWrapper_220_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_221 ( // @[package.scala 93:22:@54708.4]
    .clock(RetimeWrapper_221_clock),
    .reset(RetimeWrapper_221_reset),
    .io_flow(RetimeWrapper_221_io_flow),
    .io_in(RetimeWrapper_221_io_in),
    .io_out(RetimeWrapper_221_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_222 ( // @[package.scala 93:22:@54716.4]
    .clock(RetimeWrapper_222_clock),
    .reset(RetimeWrapper_222_reset),
    .io_flow(RetimeWrapper_222_io_flow),
    .io_in(RetimeWrapper_222_io_in),
    .io_out(RetimeWrapper_222_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_223 ( // @[package.scala 93:22:@54724.4]
    .clock(RetimeWrapper_223_clock),
    .reset(RetimeWrapper_223_reset),
    .io_flow(RetimeWrapper_223_io_flow),
    .io_in(RetimeWrapper_223_io_in),
    .io_out(RetimeWrapper_223_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_224 ( // @[package.scala 93:22:@54732.4]
    .clock(RetimeWrapper_224_clock),
    .reset(RetimeWrapper_224_reset),
    .io_flow(RetimeWrapper_224_io_flow),
    .io_in(RetimeWrapper_224_io_in),
    .io_out(RetimeWrapper_224_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_225 ( // @[package.scala 93:22:@54740.4]
    .clock(RetimeWrapper_225_clock),
    .reset(RetimeWrapper_225_reset),
    .io_flow(RetimeWrapper_225_io_flow),
    .io_in(RetimeWrapper_225_io_in),
    .io_out(RetimeWrapper_225_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_226 ( // @[package.scala 93:22:@54748.4]
    .clock(RetimeWrapper_226_clock),
    .reset(RetimeWrapper_226_reset),
    .io_flow(RetimeWrapper_226_io_flow),
    .io_in(RetimeWrapper_226_io_in),
    .io_out(RetimeWrapper_226_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_227 ( // @[package.scala 93:22:@54756.4]
    .clock(RetimeWrapper_227_clock),
    .reset(RetimeWrapper_227_reset),
    .io_flow(RetimeWrapper_227_io_flow),
    .io_in(RetimeWrapper_227_io_in),
    .io_out(RetimeWrapper_227_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_228 ( // @[package.scala 93:22:@54764.4]
    .clock(RetimeWrapper_228_clock),
    .reset(RetimeWrapper_228_reset),
    .io_flow(RetimeWrapper_228_io_flow),
    .io_in(RetimeWrapper_228_io_in),
    .io_out(RetimeWrapper_228_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_229 ( // @[package.scala 93:22:@54772.4]
    .clock(RetimeWrapper_229_clock),
    .reset(RetimeWrapper_229_reset),
    .io_flow(RetimeWrapper_229_io_flow),
    .io_in(RetimeWrapper_229_io_in),
    .io_out(RetimeWrapper_229_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_230 ( // @[package.scala 93:22:@54780.4]
    .clock(RetimeWrapper_230_clock),
    .reset(RetimeWrapper_230_reset),
    .io_flow(RetimeWrapper_230_io_flow),
    .io_in(RetimeWrapper_230_io_in),
    .io_out(RetimeWrapper_230_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_231 ( // @[package.scala 93:22:@54788.4]
    .clock(RetimeWrapper_231_clock),
    .reset(RetimeWrapper_231_reset),
    .io_flow(RetimeWrapper_231_io_flow),
    .io_in(RetimeWrapper_231_io_in),
    .io_out(RetimeWrapper_231_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_232 ( // @[package.scala 93:22:@54796.4]
    .clock(RetimeWrapper_232_clock),
    .reset(RetimeWrapper_232_reset),
    .io_flow(RetimeWrapper_232_io_flow),
    .io_in(RetimeWrapper_232_io_in),
    .io_out(RetimeWrapper_232_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_233 ( // @[package.scala 93:22:@54804.4]
    .clock(RetimeWrapper_233_clock),
    .reset(RetimeWrapper_233_reset),
    .io_flow(RetimeWrapper_233_io_flow),
    .io_in(RetimeWrapper_233_io_in),
    .io_out(RetimeWrapper_233_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_234 ( // @[package.scala 93:22:@54812.4]
    .clock(RetimeWrapper_234_clock),
    .reset(RetimeWrapper_234_reset),
    .io_flow(RetimeWrapper_234_io_flow),
    .io_in(RetimeWrapper_234_io_in),
    .io_out(RetimeWrapper_234_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_235 ( // @[package.scala 93:22:@54820.4]
    .clock(RetimeWrapper_235_clock),
    .reset(RetimeWrapper_235_reset),
    .io_flow(RetimeWrapper_235_io_flow),
    .io_in(RetimeWrapper_235_io_in),
    .io_out(RetimeWrapper_235_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_236 ( // @[package.scala 93:22:@54828.4]
    .clock(RetimeWrapper_236_clock),
    .reset(RetimeWrapper_236_reset),
    .io_flow(RetimeWrapper_236_io_flow),
    .io_in(RetimeWrapper_236_io_in),
    .io_out(RetimeWrapper_236_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_237 ( // @[package.scala 93:22:@54836.4]
    .clock(RetimeWrapper_237_clock),
    .reset(RetimeWrapper_237_reset),
    .io_flow(RetimeWrapper_237_io_flow),
    .io_in(RetimeWrapper_237_io_in),
    .io_out(RetimeWrapper_237_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_238 ( // @[package.scala 93:22:@54844.4]
    .clock(RetimeWrapper_238_clock),
    .reset(RetimeWrapper_238_reset),
    .io_flow(RetimeWrapper_238_io_flow),
    .io_in(RetimeWrapper_238_io_in),
    .io_out(RetimeWrapper_238_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_239 ( // @[package.scala 93:22:@54852.4]
    .clock(RetimeWrapper_239_clock),
    .reset(RetimeWrapper_239_reset),
    .io_flow(RetimeWrapper_239_io_flow),
    .io_in(RetimeWrapper_239_io_in),
    .io_out(RetimeWrapper_239_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_240 ( // @[package.scala 93:22:@54940.4]
    .clock(RetimeWrapper_240_clock),
    .reset(RetimeWrapper_240_reset),
    .io_flow(RetimeWrapper_240_io_flow),
    .io_in(RetimeWrapper_240_io_in),
    .io_out(RetimeWrapper_240_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_241 ( // @[package.scala 93:22:@54948.4]
    .clock(RetimeWrapper_241_clock),
    .reset(RetimeWrapper_241_reset),
    .io_flow(RetimeWrapper_241_io_flow),
    .io_in(RetimeWrapper_241_io_in),
    .io_out(RetimeWrapper_241_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_242 ( // @[package.scala 93:22:@54956.4]
    .clock(RetimeWrapper_242_clock),
    .reset(RetimeWrapper_242_reset),
    .io_flow(RetimeWrapper_242_io_flow),
    .io_in(RetimeWrapper_242_io_in),
    .io_out(RetimeWrapper_242_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_243 ( // @[package.scala 93:22:@54964.4]
    .clock(RetimeWrapper_243_clock),
    .reset(RetimeWrapper_243_reset),
    .io_flow(RetimeWrapper_243_io_flow),
    .io_in(RetimeWrapper_243_io_in),
    .io_out(RetimeWrapper_243_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_244 ( // @[package.scala 93:22:@54972.4]
    .clock(RetimeWrapper_244_clock),
    .reset(RetimeWrapper_244_reset),
    .io_flow(RetimeWrapper_244_io_flow),
    .io_in(RetimeWrapper_244_io_in),
    .io_out(RetimeWrapper_244_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_245 ( // @[package.scala 93:22:@54980.4]
    .clock(RetimeWrapper_245_clock),
    .reset(RetimeWrapper_245_reset),
    .io_flow(RetimeWrapper_245_io_flow),
    .io_in(RetimeWrapper_245_io_in),
    .io_out(RetimeWrapper_245_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_246 ( // @[package.scala 93:22:@54988.4]
    .clock(RetimeWrapper_246_clock),
    .reset(RetimeWrapper_246_reset),
    .io_flow(RetimeWrapper_246_io_flow),
    .io_in(RetimeWrapper_246_io_in),
    .io_out(RetimeWrapper_246_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_247 ( // @[package.scala 93:22:@54996.4]
    .clock(RetimeWrapper_247_clock),
    .reset(RetimeWrapper_247_reset),
    .io_flow(RetimeWrapper_247_io_flow),
    .io_in(RetimeWrapper_247_io_in),
    .io_out(RetimeWrapper_247_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_248 ( // @[package.scala 93:22:@55004.4]
    .clock(RetimeWrapper_248_clock),
    .reset(RetimeWrapper_248_reset),
    .io_flow(RetimeWrapper_248_io_flow),
    .io_in(RetimeWrapper_248_io_in),
    .io_out(RetimeWrapper_248_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_249 ( // @[package.scala 93:22:@55012.4]
    .clock(RetimeWrapper_249_clock),
    .reset(RetimeWrapper_249_reset),
    .io_flow(RetimeWrapper_249_io_flow),
    .io_in(RetimeWrapper_249_io_in),
    .io_out(RetimeWrapper_249_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_250 ( // @[package.scala 93:22:@55020.4]
    .clock(RetimeWrapper_250_clock),
    .reset(RetimeWrapper_250_reset),
    .io_flow(RetimeWrapper_250_io_flow),
    .io_in(RetimeWrapper_250_io_in),
    .io_out(RetimeWrapper_250_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_251 ( // @[package.scala 93:22:@55028.4]
    .clock(RetimeWrapper_251_clock),
    .reset(RetimeWrapper_251_reset),
    .io_flow(RetimeWrapper_251_io_flow),
    .io_in(RetimeWrapper_251_io_in),
    .io_out(RetimeWrapper_251_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_252 ( // @[package.scala 93:22:@55036.4]
    .clock(RetimeWrapper_252_clock),
    .reset(RetimeWrapper_252_reset),
    .io_flow(RetimeWrapper_252_io_flow),
    .io_in(RetimeWrapper_252_io_in),
    .io_out(RetimeWrapper_252_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_253 ( // @[package.scala 93:22:@55044.4]
    .clock(RetimeWrapper_253_clock),
    .reset(RetimeWrapper_253_reset),
    .io_flow(RetimeWrapper_253_io_flow),
    .io_in(RetimeWrapper_253_io_in),
    .io_out(RetimeWrapper_253_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_254 ( // @[package.scala 93:22:@55052.4]
    .clock(RetimeWrapper_254_clock),
    .reset(RetimeWrapper_254_reset),
    .io_flow(RetimeWrapper_254_io_flow),
    .io_in(RetimeWrapper_254_io_in),
    .io_out(RetimeWrapper_254_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_255 ( // @[package.scala 93:22:@55060.4]
    .clock(RetimeWrapper_255_clock),
    .reset(RetimeWrapper_255_reset),
    .io_flow(RetimeWrapper_255_io_flow),
    .io_in(RetimeWrapper_255_io_in),
    .io_out(RetimeWrapper_255_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_256 ( // @[package.scala 93:22:@55068.4]
    .clock(RetimeWrapper_256_clock),
    .reset(RetimeWrapper_256_reset),
    .io_flow(RetimeWrapper_256_io_flow),
    .io_in(RetimeWrapper_256_io_in),
    .io_out(RetimeWrapper_256_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_257 ( // @[package.scala 93:22:@55076.4]
    .clock(RetimeWrapper_257_clock),
    .reset(RetimeWrapper_257_reset),
    .io_flow(RetimeWrapper_257_io_flow),
    .io_in(RetimeWrapper_257_io_in),
    .io_out(RetimeWrapper_257_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_258 ( // @[package.scala 93:22:@55084.4]
    .clock(RetimeWrapper_258_clock),
    .reset(RetimeWrapper_258_reset),
    .io_flow(RetimeWrapper_258_io_flow),
    .io_in(RetimeWrapper_258_io_in),
    .io_out(RetimeWrapper_258_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_259 ( // @[package.scala 93:22:@55092.4]
    .clock(RetimeWrapper_259_clock),
    .reset(RetimeWrapper_259_reset),
    .io_flow(RetimeWrapper_259_io_flow),
    .io_in(RetimeWrapper_259_io_in),
    .io_out(RetimeWrapper_259_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_260 ( // @[package.scala 93:22:@55180.4]
    .clock(RetimeWrapper_260_clock),
    .reset(RetimeWrapper_260_reset),
    .io_flow(RetimeWrapper_260_io_flow),
    .io_in(RetimeWrapper_260_io_in),
    .io_out(RetimeWrapper_260_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_261 ( // @[package.scala 93:22:@55188.4]
    .clock(RetimeWrapper_261_clock),
    .reset(RetimeWrapper_261_reset),
    .io_flow(RetimeWrapper_261_io_flow),
    .io_in(RetimeWrapper_261_io_in),
    .io_out(RetimeWrapper_261_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_262 ( // @[package.scala 93:22:@55196.4]
    .clock(RetimeWrapper_262_clock),
    .reset(RetimeWrapper_262_reset),
    .io_flow(RetimeWrapper_262_io_flow),
    .io_in(RetimeWrapper_262_io_in),
    .io_out(RetimeWrapper_262_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_263 ( // @[package.scala 93:22:@55204.4]
    .clock(RetimeWrapper_263_clock),
    .reset(RetimeWrapper_263_reset),
    .io_flow(RetimeWrapper_263_io_flow),
    .io_in(RetimeWrapper_263_io_in),
    .io_out(RetimeWrapper_263_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_264 ( // @[package.scala 93:22:@55212.4]
    .clock(RetimeWrapper_264_clock),
    .reset(RetimeWrapper_264_reset),
    .io_flow(RetimeWrapper_264_io_flow),
    .io_in(RetimeWrapper_264_io_in),
    .io_out(RetimeWrapper_264_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_265 ( // @[package.scala 93:22:@55220.4]
    .clock(RetimeWrapper_265_clock),
    .reset(RetimeWrapper_265_reset),
    .io_flow(RetimeWrapper_265_io_flow),
    .io_in(RetimeWrapper_265_io_in),
    .io_out(RetimeWrapper_265_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_266 ( // @[package.scala 93:22:@55228.4]
    .clock(RetimeWrapper_266_clock),
    .reset(RetimeWrapper_266_reset),
    .io_flow(RetimeWrapper_266_io_flow),
    .io_in(RetimeWrapper_266_io_in),
    .io_out(RetimeWrapper_266_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_267 ( // @[package.scala 93:22:@55236.4]
    .clock(RetimeWrapper_267_clock),
    .reset(RetimeWrapper_267_reset),
    .io_flow(RetimeWrapper_267_io_flow),
    .io_in(RetimeWrapper_267_io_in),
    .io_out(RetimeWrapper_267_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_268 ( // @[package.scala 93:22:@55244.4]
    .clock(RetimeWrapper_268_clock),
    .reset(RetimeWrapper_268_reset),
    .io_flow(RetimeWrapper_268_io_flow),
    .io_in(RetimeWrapper_268_io_in),
    .io_out(RetimeWrapper_268_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_269 ( // @[package.scala 93:22:@55252.4]
    .clock(RetimeWrapper_269_clock),
    .reset(RetimeWrapper_269_reset),
    .io_flow(RetimeWrapper_269_io_flow),
    .io_in(RetimeWrapper_269_io_in),
    .io_out(RetimeWrapper_269_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_270 ( // @[package.scala 93:22:@55260.4]
    .clock(RetimeWrapper_270_clock),
    .reset(RetimeWrapper_270_reset),
    .io_flow(RetimeWrapper_270_io_flow),
    .io_in(RetimeWrapper_270_io_in),
    .io_out(RetimeWrapper_270_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_271 ( // @[package.scala 93:22:@55268.4]
    .clock(RetimeWrapper_271_clock),
    .reset(RetimeWrapper_271_reset),
    .io_flow(RetimeWrapper_271_io_flow),
    .io_in(RetimeWrapper_271_io_in),
    .io_out(RetimeWrapper_271_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_272 ( // @[package.scala 93:22:@55276.4]
    .clock(RetimeWrapper_272_clock),
    .reset(RetimeWrapper_272_reset),
    .io_flow(RetimeWrapper_272_io_flow),
    .io_in(RetimeWrapper_272_io_in),
    .io_out(RetimeWrapper_272_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_273 ( // @[package.scala 93:22:@55284.4]
    .clock(RetimeWrapper_273_clock),
    .reset(RetimeWrapper_273_reset),
    .io_flow(RetimeWrapper_273_io_flow),
    .io_in(RetimeWrapper_273_io_in),
    .io_out(RetimeWrapper_273_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_274 ( // @[package.scala 93:22:@55292.4]
    .clock(RetimeWrapper_274_clock),
    .reset(RetimeWrapper_274_reset),
    .io_flow(RetimeWrapper_274_io_flow),
    .io_in(RetimeWrapper_274_io_in),
    .io_out(RetimeWrapper_274_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_275 ( // @[package.scala 93:22:@55300.4]
    .clock(RetimeWrapper_275_clock),
    .reset(RetimeWrapper_275_reset),
    .io_flow(RetimeWrapper_275_io_flow),
    .io_in(RetimeWrapper_275_io_in),
    .io_out(RetimeWrapper_275_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_276 ( // @[package.scala 93:22:@55308.4]
    .clock(RetimeWrapper_276_clock),
    .reset(RetimeWrapper_276_reset),
    .io_flow(RetimeWrapper_276_io_flow),
    .io_in(RetimeWrapper_276_io_in),
    .io_out(RetimeWrapper_276_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_277 ( // @[package.scala 93:22:@55316.4]
    .clock(RetimeWrapper_277_clock),
    .reset(RetimeWrapper_277_reset),
    .io_flow(RetimeWrapper_277_io_flow),
    .io_in(RetimeWrapper_277_io_in),
    .io_out(RetimeWrapper_277_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_278 ( // @[package.scala 93:22:@55324.4]
    .clock(RetimeWrapper_278_clock),
    .reset(RetimeWrapper_278_reset),
    .io_flow(RetimeWrapper_278_io_flow),
    .io_in(RetimeWrapper_278_io_in),
    .io_out(RetimeWrapper_278_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_279 ( // @[package.scala 93:22:@55332.4]
    .clock(RetimeWrapper_279_clock),
    .reset(RetimeWrapper_279_reset),
    .io_flow(RetimeWrapper_279_io_flow),
    .io_in(RetimeWrapper_279_io_in),
    .io_out(RetimeWrapper_279_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_280 ( // @[package.scala 93:22:@55420.4]
    .clock(RetimeWrapper_280_clock),
    .reset(RetimeWrapper_280_reset),
    .io_flow(RetimeWrapper_280_io_flow),
    .io_in(RetimeWrapper_280_io_in),
    .io_out(RetimeWrapper_280_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_281 ( // @[package.scala 93:22:@55428.4]
    .clock(RetimeWrapper_281_clock),
    .reset(RetimeWrapper_281_reset),
    .io_flow(RetimeWrapper_281_io_flow),
    .io_in(RetimeWrapper_281_io_in),
    .io_out(RetimeWrapper_281_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_282 ( // @[package.scala 93:22:@55436.4]
    .clock(RetimeWrapper_282_clock),
    .reset(RetimeWrapper_282_reset),
    .io_flow(RetimeWrapper_282_io_flow),
    .io_in(RetimeWrapper_282_io_in),
    .io_out(RetimeWrapper_282_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_283 ( // @[package.scala 93:22:@55444.4]
    .clock(RetimeWrapper_283_clock),
    .reset(RetimeWrapper_283_reset),
    .io_flow(RetimeWrapper_283_io_flow),
    .io_in(RetimeWrapper_283_io_in),
    .io_out(RetimeWrapper_283_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_284 ( // @[package.scala 93:22:@55452.4]
    .clock(RetimeWrapper_284_clock),
    .reset(RetimeWrapper_284_reset),
    .io_flow(RetimeWrapper_284_io_flow),
    .io_in(RetimeWrapper_284_io_in),
    .io_out(RetimeWrapper_284_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_285 ( // @[package.scala 93:22:@55460.4]
    .clock(RetimeWrapper_285_clock),
    .reset(RetimeWrapper_285_reset),
    .io_flow(RetimeWrapper_285_io_flow),
    .io_in(RetimeWrapper_285_io_in),
    .io_out(RetimeWrapper_285_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_286 ( // @[package.scala 93:22:@55468.4]
    .clock(RetimeWrapper_286_clock),
    .reset(RetimeWrapper_286_reset),
    .io_flow(RetimeWrapper_286_io_flow),
    .io_in(RetimeWrapper_286_io_in),
    .io_out(RetimeWrapper_286_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_287 ( // @[package.scala 93:22:@55476.4]
    .clock(RetimeWrapper_287_clock),
    .reset(RetimeWrapper_287_reset),
    .io_flow(RetimeWrapper_287_io_flow),
    .io_in(RetimeWrapper_287_io_in),
    .io_out(RetimeWrapper_287_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_288 ( // @[package.scala 93:22:@55484.4]
    .clock(RetimeWrapper_288_clock),
    .reset(RetimeWrapper_288_reset),
    .io_flow(RetimeWrapper_288_io_flow),
    .io_in(RetimeWrapper_288_io_in),
    .io_out(RetimeWrapper_288_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_289 ( // @[package.scala 93:22:@55492.4]
    .clock(RetimeWrapper_289_clock),
    .reset(RetimeWrapper_289_reset),
    .io_flow(RetimeWrapper_289_io_flow),
    .io_in(RetimeWrapper_289_io_in),
    .io_out(RetimeWrapper_289_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_290 ( // @[package.scala 93:22:@55500.4]
    .clock(RetimeWrapper_290_clock),
    .reset(RetimeWrapper_290_reset),
    .io_flow(RetimeWrapper_290_io_flow),
    .io_in(RetimeWrapper_290_io_in),
    .io_out(RetimeWrapper_290_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_291 ( // @[package.scala 93:22:@55508.4]
    .clock(RetimeWrapper_291_clock),
    .reset(RetimeWrapper_291_reset),
    .io_flow(RetimeWrapper_291_io_flow),
    .io_in(RetimeWrapper_291_io_in),
    .io_out(RetimeWrapper_291_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_292 ( // @[package.scala 93:22:@55516.4]
    .clock(RetimeWrapper_292_clock),
    .reset(RetimeWrapper_292_reset),
    .io_flow(RetimeWrapper_292_io_flow),
    .io_in(RetimeWrapper_292_io_in),
    .io_out(RetimeWrapper_292_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_293 ( // @[package.scala 93:22:@55524.4]
    .clock(RetimeWrapper_293_clock),
    .reset(RetimeWrapper_293_reset),
    .io_flow(RetimeWrapper_293_io_flow),
    .io_in(RetimeWrapper_293_io_in),
    .io_out(RetimeWrapper_293_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_294 ( // @[package.scala 93:22:@55532.4]
    .clock(RetimeWrapper_294_clock),
    .reset(RetimeWrapper_294_reset),
    .io_flow(RetimeWrapper_294_io_flow),
    .io_in(RetimeWrapper_294_io_in),
    .io_out(RetimeWrapper_294_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_295 ( // @[package.scala 93:22:@55540.4]
    .clock(RetimeWrapper_295_clock),
    .reset(RetimeWrapper_295_reset),
    .io_flow(RetimeWrapper_295_io_flow),
    .io_in(RetimeWrapper_295_io_in),
    .io_out(RetimeWrapper_295_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_296 ( // @[package.scala 93:22:@55548.4]
    .clock(RetimeWrapper_296_clock),
    .reset(RetimeWrapper_296_reset),
    .io_flow(RetimeWrapper_296_io_flow),
    .io_in(RetimeWrapper_296_io_in),
    .io_out(RetimeWrapper_296_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_297 ( // @[package.scala 93:22:@55556.4]
    .clock(RetimeWrapper_297_clock),
    .reset(RetimeWrapper_297_reset),
    .io_flow(RetimeWrapper_297_io_flow),
    .io_in(RetimeWrapper_297_io_in),
    .io_out(RetimeWrapper_297_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_298 ( // @[package.scala 93:22:@55564.4]
    .clock(RetimeWrapper_298_clock),
    .reset(RetimeWrapper_298_reset),
    .io_flow(RetimeWrapper_298_io_flow),
    .io_in(RetimeWrapper_298_io_in),
    .io_out(RetimeWrapper_298_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_299 ( // @[package.scala 93:22:@55572.4]
    .clock(RetimeWrapper_299_clock),
    .reset(RetimeWrapper_299_reset),
    .io_flow(RetimeWrapper_299_io_flow),
    .io_in(RetimeWrapper_299_io_in),
    .io_out(RetimeWrapper_299_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_300 ( // @[package.scala 93:22:@55660.4]
    .clock(RetimeWrapper_300_clock),
    .reset(RetimeWrapper_300_reset),
    .io_flow(RetimeWrapper_300_io_flow),
    .io_in(RetimeWrapper_300_io_in),
    .io_out(RetimeWrapper_300_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_301 ( // @[package.scala 93:22:@55668.4]
    .clock(RetimeWrapper_301_clock),
    .reset(RetimeWrapper_301_reset),
    .io_flow(RetimeWrapper_301_io_flow),
    .io_in(RetimeWrapper_301_io_in),
    .io_out(RetimeWrapper_301_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_302 ( // @[package.scala 93:22:@55676.4]
    .clock(RetimeWrapper_302_clock),
    .reset(RetimeWrapper_302_reset),
    .io_flow(RetimeWrapper_302_io_flow),
    .io_in(RetimeWrapper_302_io_in),
    .io_out(RetimeWrapper_302_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_303 ( // @[package.scala 93:22:@55684.4]
    .clock(RetimeWrapper_303_clock),
    .reset(RetimeWrapper_303_reset),
    .io_flow(RetimeWrapper_303_io_flow),
    .io_in(RetimeWrapper_303_io_in),
    .io_out(RetimeWrapper_303_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_304 ( // @[package.scala 93:22:@55692.4]
    .clock(RetimeWrapper_304_clock),
    .reset(RetimeWrapper_304_reset),
    .io_flow(RetimeWrapper_304_io_flow),
    .io_in(RetimeWrapper_304_io_in),
    .io_out(RetimeWrapper_304_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_305 ( // @[package.scala 93:22:@55700.4]
    .clock(RetimeWrapper_305_clock),
    .reset(RetimeWrapper_305_reset),
    .io_flow(RetimeWrapper_305_io_flow),
    .io_in(RetimeWrapper_305_io_in),
    .io_out(RetimeWrapper_305_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_306 ( // @[package.scala 93:22:@55708.4]
    .clock(RetimeWrapper_306_clock),
    .reset(RetimeWrapper_306_reset),
    .io_flow(RetimeWrapper_306_io_flow),
    .io_in(RetimeWrapper_306_io_in),
    .io_out(RetimeWrapper_306_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_307 ( // @[package.scala 93:22:@55716.4]
    .clock(RetimeWrapper_307_clock),
    .reset(RetimeWrapper_307_reset),
    .io_flow(RetimeWrapper_307_io_flow),
    .io_in(RetimeWrapper_307_io_in),
    .io_out(RetimeWrapper_307_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_308 ( // @[package.scala 93:22:@55724.4]
    .clock(RetimeWrapper_308_clock),
    .reset(RetimeWrapper_308_reset),
    .io_flow(RetimeWrapper_308_io_flow),
    .io_in(RetimeWrapper_308_io_in),
    .io_out(RetimeWrapper_308_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_309 ( // @[package.scala 93:22:@55732.4]
    .clock(RetimeWrapper_309_clock),
    .reset(RetimeWrapper_309_reset),
    .io_flow(RetimeWrapper_309_io_flow),
    .io_in(RetimeWrapper_309_io_in),
    .io_out(RetimeWrapper_309_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_310 ( // @[package.scala 93:22:@55740.4]
    .clock(RetimeWrapper_310_clock),
    .reset(RetimeWrapper_310_reset),
    .io_flow(RetimeWrapper_310_io_flow),
    .io_in(RetimeWrapper_310_io_in),
    .io_out(RetimeWrapper_310_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_311 ( // @[package.scala 93:22:@55748.4]
    .clock(RetimeWrapper_311_clock),
    .reset(RetimeWrapper_311_reset),
    .io_flow(RetimeWrapper_311_io_flow),
    .io_in(RetimeWrapper_311_io_in),
    .io_out(RetimeWrapper_311_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_312 ( // @[package.scala 93:22:@55756.4]
    .clock(RetimeWrapper_312_clock),
    .reset(RetimeWrapper_312_reset),
    .io_flow(RetimeWrapper_312_io_flow),
    .io_in(RetimeWrapper_312_io_in),
    .io_out(RetimeWrapper_312_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_313 ( // @[package.scala 93:22:@55764.4]
    .clock(RetimeWrapper_313_clock),
    .reset(RetimeWrapper_313_reset),
    .io_flow(RetimeWrapper_313_io_flow),
    .io_in(RetimeWrapper_313_io_in),
    .io_out(RetimeWrapper_313_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_314 ( // @[package.scala 93:22:@55772.4]
    .clock(RetimeWrapper_314_clock),
    .reset(RetimeWrapper_314_reset),
    .io_flow(RetimeWrapper_314_io_flow),
    .io_in(RetimeWrapper_314_io_in),
    .io_out(RetimeWrapper_314_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_315 ( // @[package.scala 93:22:@55780.4]
    .clock(RetimeWrapper_315_clock),
    .reset(RetimeWrapper_315_reset),
    .io_flow(RetimeWrapper_315_io_flow),
    .io_in(RetimeWrapper_315_io_in),
    .io_out(RetimeWrapper_315_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_316 ( // @[package.scala 93:22:@55788.4]
    .clock(RetimeWrapper_316_clock),
    .reset(RetimeWrapper_316_reset),
    .io_flow(RetimeWrapper_316_io_flow),
    .io_in(RetimeWrapper_316_io_in),
    .io_out(RetimeWrapper_316_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_317 ( // @[package.scala 93:22:@55796.4]
    .clock(RetimeWrapper_317_clock),
    .reset(RetimeWrapper_317_reset),
    .io_flow(RetimeWrapper_317_io_flow),
    .io_in(RetimeWrapper_317_io_in),
    .io_out(RetimeWrapper_317_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_318 ( // @[package.scala 93:22:@55804.4]
    .clock(RetimeWrapper_318_clock),
    .reset(RetimeWrapper_318_reset),
    .io_flow(RetimeWrapper_318_io_flow),
    .io_in(RetimeWrapper_318_io_in),
    .io_out(RetimeWrapper_318_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_319 ( // @[package.scala 93:22:@55812.4]
    .clock(RetimeWrapper_319_clock),
    .reset(RetimeWrapper_319_reset),
    .io_flow(RetimeWrapper_319_io_flow),
    .io_in(RetimeWrapper_319_io_in),
    .io_out(RetimeWrapper_319_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_320 ( // @[package.scala 93:22:@55900.4]
    .clock(RetimeWrapper_320_clock),
    .reset(RetimeWrapper_320_reset),
    .io_flow(RetimeWrapper_320_io_flow),
    .io_in(RetimeWrapper_320_io_in),
    .io_out(RetimeWrapper_320_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_321 ( // @[package.scala 93:22:@55908.4]
    .clock(RetimeWrapper_321_clock),
    .reset(RetimeWrapper_321_reset),
    .io_flow(RetimeWrapper_321_io_flow),
    .io_in(RetimeWrapper_321_io_in),
    .io_out(RetimeWrapper_321_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_322 ( // @[package.scala 93:22:@55916.4]
    .clock(RetimeWrapper_322_clock),
    .reset(RetimeWrapper_322_reset),
    .io_flow(RetimeWrapper_322_io_flow),
    .io_in(RetimeWrapper_322_io_in),
    .io_out(RetimeWrapper_322_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_323 ( // @[package.scala 93:22:@55924.4]
    .clock(RetimeWrapper_323_clock),
    .reset(RetimeWrapper_323_reset),
    .io_flow(RetimeWrapper_323_io_flow),
    .io_in(RetimeWrapper_323_io_in),
    .io_out(RetimeWrapper_323_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_324 ( // @[package.scala 93:22:@55932.4]
    .clock(RetimeWrapper_324_clock),
    .reset(RetimeWrapper_324_reset),
    .io_flow(RetimeWrapper_324_io_flow),
    .io_in(RetimeWrapper_324_io_in),
    .io_out(RetimeWrapper_324_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_325 ( // @[package.scala 93:22:@55940.4]
    .clock(RetimeWrapper_325_clock),
    .reset(RetimeWrapper_325_reset),
    .io_flow(RetimeWrapper_325_io_flow),
    .io_in(RetimeWrapper_325_io_in),
    .io_out(RetimeWrapper_325_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_326 ( // @[package.scala 93:22:@55948.4]
    .clock(RetimeWrapper_326_clock),
    .reset(RetimeWrapper_326_reset),
    .io_flow(RetimeWrapper_326_io_flow),
    .io_in(RetimeWrapper_326_io_in),
    .io_out(RetimeWrapper_326_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_327 ( // @[package.scala 93:22:@55956.4]
    .clock(RetimeWrapper_327_clock),
    .reset(RetimeWrapper_327_reset),
    .io_flow(RetimeWrapper_327_io_flow),
    .io_in(RetimeWrapper_327_io_in),
    .io_out(RetimeWrapper_327_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_328 ( // @[package.scala 93:22:@55964.4]
    .clock(RetimeWrapper_328_clock),
    .reset(RetimeWrapper_328_reset),
    .io_flow(RetimeWrapper_328_io_flow),
    .io_in(RetimeWrapper_328_io_in),
    .io_out(RetimeWrapper_328_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_329 ( // @[package.scala 93:22:@55972.4]
    .clock(RetimeWrapper_329_clock),
    .reset(RetimeWrapper_329_reset),
    .io_flow(RetimeWrapper_329_io_flow),
    .io_in(RetimeWrapper_329_io_in),
    .io_out(RetimeWrapper_329_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_330 ( // @[package.scala 93:22:@55980.4]
    .clock(RetimeWrapper_330_clock),
    .reset(RetimeWrapper_330_reset),
    .io_flow(RetimeWrapper_330_io_flow),
    .io_in(RetimeWrapper_330_io_in),
    .io_out(RetimeWrapper_330_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_331 ( // @[package.scala 93:22:@55988.4]
    .clock(RetimeWrapper_331_clock),
    .reset(RetimeWrapper_331_reset),
    .io_flow(RetimeWrapper_331_io_flow),
    .io_in(RetimeWrapper_331_io_in),
    .io_out(RetimeWrapper_331_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_332 ( // @[package.scala 93:22:@55996.4]
    .clock(RetimeWrapper_332_clock),
    .reset(RetimeWrapper_332_reset),
    .io_flow(RetimeWrapper_332_io_flow),
    .io_in(RetimeWrapper_332_io_in),
    .io_out(RetimeWrapper_332_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_333 ( // @[package.scala 93:22:@56004.4]
    .clock(RetimeWrapper_333_clock),
    .reset(RetimeWrapper_333_reset),
    .io_flow(RetimeWrapper_333_io_flow),
    .io_in(RetimeWrapper_333_io_in),
    .io_out(RetimeWrapper_333_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_334 ( // @[package.scala 93:22:@56012.4]
    .clock(RetimeWrapper_334_clock),
    .reset(RetimeWrapper_334_reset),
    .io_flow(RetimeWrapper_334_io_flow),
    .io_in(RetimeWrapper_334_io_in),
    .io_out(RetimeWrapper_334_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_335 ( // @[package.scala 93:22:@56020.4]
    .clock(RetimeWrapper_335_clock),
    .reset(RetimeWrapper_335_reset),
    .io_flow(RetimeWrapper_335_io_flow),
    .io_in(RetimeWrapper_335_io_in),
    .io_out(RetimeWrapper_335_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_336 ( // @[package.scala 93:22:@56028.4]
    .clock(RetimeWrapper_336_clock),
    .reset(RetimeWrapper_336_reset),
    .io_flow(RetimeWrapper_336_io_flow),
    .io_in(RetimeWrapper_336_io_in),
    .io_out(RetimeWrapper_336_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_337 ( // @[package.scala 93:22:@56036.4]
    .clock(RetimeWrapper_337_clock),
    .reset(RetimeWrapper_337_reset),
    .io_flow(RetimeWrapper_337_io_flow),
    .io_in(RetimeWrapper_337_io_in),
    .io_out(RetimeWrapper_337_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_338 ( // @[package.scala 93:22:@56044.4]
    .clock(RetimeWrapper_338_clock),
    .reset(RetimeWrapper_338_reset),
    .io_flow(RetimeWrapper_338_io_flow),
    .io_in(RetimeWrapper_338_io_in),
    .io_out(RetimeWrapper_338_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_339 ( // @[package.scala 93:22:@56052.4]
    .clock(RetimeWrapper_339_clock),
    .reset(RetimeWrapper_339_reset),
    .io_flow(RetimeWrapper_339_io_flow),
    .io_in(RetimeWrapper_339_io_in),
    .io_out(RetimeWrapper_339_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_340 ( // @[package.scala 93:22:@56140.4]
    .clock(RetimeWrapper_340_clock),
    .reset(RetimeWrapper_340_reset),
    .io_flow(RetimeWrapper_340_io_flow),
    .io_in(RetimeWrapper_340_io_in),
    .io_out(RetimeWrapper_340_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_341 ( // @[package.scala 93:22:@56148.4]
    .clock(RetimeWrapper_341_clock),
    .reset(RetimeWrapper_341_reset),
    .io_flow(RetimeWrapper_341_io_flow),
    .io_in(RetimeWrapper_341_io_in),
    .io_out(RetimeWrapper_341_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_342 ( // @[package.scala 93:22:@56156.4]
    .clock(RetimeWrapper_342_clock),
    .reset(RetimeWrapper_342_reset),
    .io_flow(RetimeWrapper_342_io_flow),
    .io_in(RetimeWrapper_342_io_in),
    .io_out(RetimeWrapper_342_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_343 ( // @[package.scala 93:22:@56164.4]
    .clock(RetimeWrapper_343_clock),
    .reset(RetimeWrapper_343_reset),
    .io_flow(RetimeWrapper_343_io_flow),
    .io_in(RetimeWrapper_343_io_in),
    .io_out(RetimeWrapper_343_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_344 ( // @[package.scala 93:22:@56172.4]
    .clock(RetimeWrapper_344_clock),
    .reset(RetimeWrapper_344_reset),
    .io_flow(RetimeWrapper_344_io_flow),
    .io_in(RetimeWrapper_344_io_in),
    .io_out(RetimeWrapper_344_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_345 ( // @[package.scala 93:22:@56180.4]
    .clock(RetimeWrapper_345_clock),
    .reset(RetimeWrapper_345_reset),
    .io_flow(RetimeWrapper_345_io_flow),
    .io_in(RetimeWrapper_345_io_in),
    .io_out(RetimeWrapper_345_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_346 ( // @[package.scala 93:22:@56188.4]
    .clock(RetimeWrapper_346_clock),
    .reset(RetimeWrapper_346_reset),
    .io_flow(RetimeWrapper_346_io_flow),
    .io_in(RetimeWrapper_346_io_in),
    .io_out(RetimeWrapper_346_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_347 ( // @[package.scala 93:22:@56196.4]
    .clock(RetimeWrapper_347_clock),
    .reset(RetimeWrapper_347_reset),
    .io_flow(RetimeWrapper_347_io_flow),
    .io_in(RetimeWrapper_347_io_in),
    .io_out(RetimeWrapper_347_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_348 ( // @[package.scala 93:22:@56204.4]
    .clock(RetimeWrapper_348_clock),
    .reset(RetimeWrapper_348_reset),
    .io_flow(RetimeWrapper_348_io_flow),
    .io_in(RetimeWrapper_348_io_in),
    .io_out(RetimeWrapper_348_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_349 ( // @[package.scala 93:22:@56212.4]
    .clock(RetimeWrapper_349_clock),
    .reset(RetimeWrapper_349_reset),
    .io_flow(RetimeWrapper_349_io_flow),
    .io_in(RetimeWrapper_349_io_in),
    .io_out(RetimeWrapper_349_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_350 ( // @[package.scala 93:22:@56220.4]
    .clock(RetimeWrapper_350_clock),
    .reset(RetimeWrapper_350_reset),
    .io_flow(RetimeWrapper_350_io_flow),
    .io_in(RetimeWrapper_350_io_in),
    .io_out(RetimeWrapper_350_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_351 ( // @[package.scala 93:22:@56228.4]
    .clock(RetimeWrapper_351_clock),
    .reset(RetimeWrapper_351_reset),
    .io_flow(RetimeWrapper_351_io_flow),
    .io_in(RetimeWrapper_351_io_in),
    .io_out(RetimeWrapper_351_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_352 ( // @[package.scala 93:22:@56236.4]
    .clock(RetimeWrapper_352_clock),
    .reset(RetimeWrapper_352_reset),
    .io_flow(RetimeWrapper_352_io_flow),
    .io_in(RetimeWrapper_352_io_in),
    .io_out(RetimeWrapper_352_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_353 ( // @[package.scala 93:22:@56244.4]
    .clock(RetimeWrapper_353_clock),
    .reset(RetimeWrapper_353_reset),
    .io_flow(RetimeWrapper_353_io_flow),
    .io_in(RetimeWrapper_353_io_in),
    .io_out(RetimeWrapper_353_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_354 ( // @[package.scala 93:22:@56252.4]
    .clock(RetimeWrapper_354_clock),
    .reset(RetimeWrapper_354_reset),
    .io_flow(RetimeWrapper_354_io_flow),
    .io_in(RetimeWrapper_354_io_in),
    .io_out(RetimeWrapper_354_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_355 ( // @[package.scala 93:22:@56260.4]
    .clock(RetimeWrapper_355_clock),
    .reset(RetimeWrapper_355_reset),
    .io_flow(RetimeWrapper_355_io_flow),
    .io_in(RetimeWrapper_355_io_in),
    .io_out(RetimeWrapper_355_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_356 ( // @[package.scala 93:22:@56268.4]
    .clock(RetimeWrapper_356_clock),
    .reset(RetimeWrapper_356_reset),
    .io_flow(RetimeWrapper_356_io_flow),
    .io_in(RetimeWrapper_356_io_in),
    .io_out(RetimeWrapper_356_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_357 ( // @[package.scala 93:22:@56276.4]
    .clock(RetimeWrapper_357_clock),
    .reset(RetimeWrapper_357_reset),
    .io_flow(RetimeWrapper_357_io_flow),
    .io_in(RetimeWrapper_357_io_in),
    .io_out(RetimeWrapper_357_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_358 ( // @[package.scala 93:22:@56284.4]
    .clock(RetimeWrapper_358_clock),
    .reset(RetimeWrapper_358_reset),
    .io_flow(RetimeWrapper_358_io_flow),
    .io_in(RetimeWrapper_358_io_in),
    .io_out(RetimeWrapper_358_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_359 ( // @[package.scala 93:22:@56292.4]
    .clock(RetimeWrapper_359_clock),
    .reset(RetimeWrapper_359_reset),
    .io_flow(RetimeWrapper_359_io_flow),
    .io_in(RetimeWrapper_359_io_in),
    .io_out(RetimeWrapper_359_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_360 ( // @[package.scala 93:22:@56380.4]
    .clock(RetimeWrapper_360_clock),
    .reset(RetimeWrapper_360_reset),
    .io_flow(RetimeWrapper_360_io_flow),
    .io_in(RetimeWrapper_360_io_in),
    .io_out(RetimeWrapper_360_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_361 ( // @[package.scala 93:22:@56388.4]
    .clock(RetimeWrapper_361_clock),
    .reset(RetimeWrapper_361_reset),
    .io_flow(RetimeWrapper_361_io_flow),
    .io_in(RetimeWrapper_361_io_in),
    .io_out(RetimeWrapper_361_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_362 ( // @[package.scala 93:22:@56396.4]
    .clock(RetimeWrapper_362_clock),
    .reset(RetimeWrapper_362_reset),
    .io_flow(RetimeWrapper_362_io_flow),
    .io_in(RetimeWrapper_362_io_in),
    .io_out(RetimeWrapper_362_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_363 ( // @[package.scala 93:22:@56404.4]
    .clock(RetimeWrapper_363_clock),
    .reset(RetimeWrapper_363_reset),
    .io_flow(RetimeWrapper_363_io_flow),
    .io_in(RetimeWrapper_363_io_in),
    .io_out(RetimeWrapper_363_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_364 ( // @[package.scala 93:22:@56412.4]
    .clock(RetimeWrapper_364_clock),
    .reset(RetimeWrapper_364_reset),
    .io_flow(RetimeWrapper_364_io_flow),
    .io_in(RetimeWrapper_364_io_in),
    .io_out(RetimeWrapper_364_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_365 ( // @[package.scala 93:22:@56420.4]
    .clock(RetimeWrapper_365_clock),
    .reset(RetimeWrapper_365_reset),
    .io_flow(RetimeWrapper_365_io_flow),
    .io_in(RetimeWrapper_365_io_in),
    .io_out(RetimeWrapper_365_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_366 ( // @[package.scala 93:22:@56428.4]
    .clock(RetimeWrapper_366_clock),
    .reset(RetimeWrapper_366_reset),
    .io_flow(RetimeWrapper_366_io_flow),
    .io_in(RetimeWrapper_366_io_in),
    .io_out(RetimeWrapper_366_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_367 ( // @[package.scala 93:22:@56436.4]
    .clock(RetimeWrapper_367_clock),
    .reset(RetimeWrapper_367_reset),
    .io_flow(RetimeWrapper_367_io_flow),
    .io_in(RetimeWrapper_367_io_in),
    .io_out(RetimeWrapper_367_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_368 ( // @[package.scala 93:22:@56444.4]
    .clock(RetimeWrapper_368_clock),
    .reset(RetimeWrapper_368_reset),
    .io_flow(RetimeWrapper_368_io_flow),
    .io_in(RetimeWrapper_368_io_in),
    .io_out(RetimeWrapper_368_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_369 ( // @[package.scala 93:22:@56452.4]
    .clock(RetimeWrapper_369_clock),
    .reset(RetimeWrapper_369_reset),
    .io_flow(RetimeWrapper_369_io_flow),
    .io_in(RetimeWrapper_369_io_in),
    .io_out(RetimeWrapper_369_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_370 ( // @[package.scala 93:22:@56460.4]
    .clock(RetimeWrapper_370_clock),
    .reset(RetimeWrapper_370_reset),
    .io_flow(RetimeWrapper_370_io_flow),
    .io_in(RetimeWrapper_370_io_in),
    .io_out(RetimeWrapper_370_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_371 ( // @[package.scala 93:22:@56468.4]
    .clock(RetimeWrapper_371_clock),
    .reset(RetimeWrapper_371_reset),
    .io_flow(RetimeWrapper_371_io_flow),
    .io_in(RetimeWrapper_371_io_in),
    .io_out(RetimeWrapper_371_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_372 ( // @[package.scala 93:22:@56476.4]
    .clock(RetimeWrapper_372_clock),
    .reset(RetimeWrapper_372_reset),
    .io_flow(RetimeWrapper_372_io_flow),
    .io_in(RetimeWrapper_372_io_in),
    .io_out(RetimeWrapper_372_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_373 ( // @[package.scala 93:22:@56484.4]
    .clock(RetimeWrapper_373_clock),
    .reset(RetimeWrapper_373_reset),
    .io_flow(RetimeWrapper_373_io_flow),
    .io_in(RetimeWrapper_373_io_in),
    .io_out(RetimeWrapper_373_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_374 ( // @[package.scala 93:22:@56492.4]
    .clock(RetimeWrapper_374_clock),
    .reset(RetimeWrapper_374_reset),
    .io_flow(RetimeWrapper_374_io_flow),
    .io_in(RetimeWrapper_374_io_in),
    .io_out(RetimeWrapper_374_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_375 ( // @[package.scala 93:22:@56500.4]
    .clock(RetimeWrapper_375_clock),
    .reset(RetimeWrapper_375_reset),
    .io_flow(RetimeWrapper_375_io_flow),
    .io_in(RetimeWrapper_375_io_in),
    .io_out(RetimeWrapper_375_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_376 ( // @[package.scala 93:22:@56508.4]
    .clock(RetimeWrapper_376_clock),
    .reset(RetimeWrapper_376_reset),
    .io_flow(RetimeWrapper_376_io_flow),
    .io_in(RetimeWrapper_376_io_in),
    .io_out(RetimeWrapper_376_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_377 ( // @[package.scala 93:22:@56516.4]
    .clock(RetimeWrapper_377_clock),
    .reset(RetimeWrapper_377_reset),
    .io_flow(RetimeWrapper_377_io_flow),
    .io_in(RetimeWrapper_377_io_in),
    .io_out(RetimeWrapper_377_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_378 ( // @[package.scala 93:22:@56524.4]
    .clock(RetimeWrapper_378_clock),
    .reset(RetimeWrapper_378_reset),
    .io_flow(RetimeWrapper_378_io_flow),
    .io_in(RetimeWrapper_378_io_in),
    .io_out(RetimeWrapper_378_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_379 ( // @[package.scala 93:22:@56532.4]
    .clock(RetimeWrapper_379_clock),
    .reset(RetimeWrapper_379_reset),
    .io_flow(RetimeWrapper_379_io_flow),
    .io_in(RetimeWrapper_379_io_in),
    .io_out(RetimeWrapper_379_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_380 ( // @[package.scala 93:22:@56620.4]
    .clock(RetimeWrapper_380_clock),
    .reset(RetimeWrapper_380_reset),
    .io_flow(RetimeWrapper_380_io_flow),
    .io_in(RetimeWrapper_380_io_in),
    .io_out(RetimeWrapper_380_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_381 ( // @[package.scala 93:22:@56628.4]
    .clock(RetimeWrapper_381_clock),
    .reset(RetimeWrapper_381_reset),
    .io_flow(RetimeWrapper_381_io_flow),
    .io_in(RetimeWrapper_381_io_in),
    .io_out(RetimeWrapper_381_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_382 ( // @[package.scala 93:22:@56636.4]
    .clock(RetimeWrapper_382_clock),
    .reset(RetimeWrapper_382_reset),
    .io_flow(RetimeWrapper_382_io_flow),
    .io_in(RetimeWrapper_382_io_in),
    .io_out(RetimeWrapper_382_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_383 ( // @[package.scala 93:22:@56644.4]
    .clock(RetimeWrapper_383_clock),
    .reset(RetimeWrapper_383_reset),
    .io_flow(RetimeWrapper_383_io_flow),
    .io_in(RetimeWrapper_383_io_in),
    .io_out(RetimeWrapper_383_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_384 ( // @[package.scala 93:22:@56652.4]
    .clock(RetimeWrapper_384_clock),
    .reset(RetimeWrapper_384_reset),
    .io_flow(RetimeWrapper_384_io_flow),
    .io_in(RetimeWrapper_384_io_in),
    .io_out(RetimeWrapper_384_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_385 ( // @[package.scala 93:22:@56660.4]
    .clock(RetimeWrapper_385_clock),
    .reset(RetimeWrapper_385_reset),
    .io_flow(RetimeWrapper_385_io_flow),
    .io_in(RetimeWrapper_385_io_in),
    .io_out(RetimeWrapper_385_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_386 ( // @[package.scala 93:22:@56668.4]
    .clock(RetimeWrapper_386_clock),
    .reset(RetimeWrapper_386_reset),
    .io_flow(RetimeWrapper_386_io_flow),
    .io_in(RetimeWrapper_386_io_in),
    .io_out(RetimeWrapper_386_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_387 ( // @[package.scala 93:22:@56676.4]
    .clock(RetimeWrapper_387_clock),
    .reset(RetimeWrapper_387_reset),
    .io_flow(RetimeWrapper_387_io_flow),
    .io_in(RetimeWrapper_387_io_in),
    .io_out(RetimeWrapper_387_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_388 ( // @[package.scala 93:22:@56684.4]
    .clock(RetimeWrapper_388_clock),
    .reset(RetimeWrapper_388_reset),
    .io_flow(RetimeWrapper_388_io_flow),
    .io_in(RetimeWrapper_388_io_in),
    .io_out(RetimeWrapper_388_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_389 ( // @[package.scala 93:22:@56692.4]
    .clock(RetimeWrapper_389_clock),
    .reset(RetimeWrapper_389_reset),
    .io_flow(RetimeWrapper_389_io_flow),
    .io_in(RetimeWrapper_389_io_in),
    .io_out(RetimeWrapper_389_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_390 ( // @[package.scala 93:22:@56700.4]
    .clock(RetimeWrapper_390_clock),
    .reset(RetimeWrapper_390_reset),
    .io_flow(RetimeWrapper_390_io_flow),
    .io_in(RetimeWrapper_390_io_in),
    .io_out(RetimeWrapper_390_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_391 ( // @[package.scala 93:22:@56708.4]
    .clock(RetimeWrapper_391_clock),
    .reset(RetimeWrapper_391_reset),
    .io_flow(RetimeWrapper_391_io_flow),
    .io_in(RetimeWrapper_391_io_in),
    .io_out(RetimeWrapper_391_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_392 ( // @[package.scala 93:22:@56716.4]
    .clock(RetimeWrapper_392_clock),
    .reset(RetimeWrapper_392_reset),
    .io_flow(RetimeWrapper_392_io_flow),
    .io_in(RetimeWrapper_392_io_in),
    .io_out(RetimeWrapper_392_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_393 ( // @[package.scala 93:22:@56724.4]
    .clock(RetimeWrapper_393_clock),
    .reset(RetimeWrapper_393_reset),
    .io_flow(RetimeWrapper_393_io_flow),
    .io_in(RetimeWrapper_393_io_in),
    .io_out(RetimeWrapper_393_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_394 ( // @[package.scala 93:22:@56732.4]
    .clock(RetimeWrapper_394_clock),
    .reset(RetimeWrapper_394_reset),
    .io_flow(RetimeWrapper_394_io_flow),
    .io_in(RetimeWrapper_394_io_in),
    .io_out(RetimeWrapper_394_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_395 ( // @[package.scala 93:22:@56740.4]
    .clock(RetimeWrapper_395_clock),
    .reset(RetimeWrapper_395_reset),
    .io_flow(RetimeWrapper_395_io_flow),
    .io_in(RetimeWrapper_395_io_in),
    .io_out(RetimeWrapper_395_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_396 ( // @[package.scala 93:22:@56748.4]
    .clock(RetimeWrapper_396_clock),
    .reset(RetimeWrapper_396_reset),
    .io_flow(RetimeWrapper_396_io_flow),
    .io_in(RetimeWrapper_396_io_in),
    .io_out(RetimeWrapper_396_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_397 ( // @[package.scala 93:22:@56756.4]
    .clock(RetimeWrapper_397_clock),
    .reset(RetimeWrapper_397_reset),
    .io_flow(RetimeWrapper_397_io_flow),
    .io_in(RetimeWrapper_397_io_in),
    .io_out(RetimeWrapper_397_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_398 ( // @[package.scala 93:22:@56764.4]
    .clock(RetimeWrapper_398_clock),
    .reset(RetimeWrapper_398_reset),
    .io_flow(RetimeWrapper_398_io_flow),
    .io_in(RetimeWrapper_398_io_in),
    .io_out(RetimeWrapper_398_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_399 ( // @[package.scala 93:22:@56772.4]
    .clock(RetimeWrapper_399_clock),
    .reset(RetimeWrapper_399_reset),
    .io_flow(RetimeWrapper_399_io_flow),
    .io_in(RetimeWrapper_399_io_in),
    .io_out(RetimeWrapper_399_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_400 ( // @[package.scala 93:22:@56860.4]
    .clock(RetimeWrapper_400_clock),
    .reset(RetimeWrapper_400_reset),
    .io_flow(RetimeWrapper_400_io_flow),
    .io_in(RetimeWrapper_400_io_in),
    .io_out(RetimeWrapper_400_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_401 ( // @[package.scala 93:22:@56868.4]
    .clock(RetimeWrapper_401_clock),
    .reset(RetimeWrapper_401_reset),
    .io_flow(RetimeWrapper_401_io_flow),
    .io_in(RetimeWrapper_401_io_in),
    .io_out(RetimeWrapper_401_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_402 ( // @[package.scala 93:22:@56876.4]
    .clock(RetimeWrapper_402_clock),
    .reset(RetimeWrapper_402_reset),
    .io_flow(RetimeWrapper_402_io_flow),
    .io_in(RetimeWrapper_402_io_in),
    .io_out(RetimeWrapper_402_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_403 ( // @[package.scala 93:22:@56884.4]
    .clock(RetimeWrapper_403_clock),
    .reset(RetimeWrapper_403_reset),
    .io_flow(RetimeWrapper_403_io_flow),
    .io_in(RetimeWrapper_403_io_in),
    .io_out(RetimeWrapper_403_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_404 ( // @[package.scala 93:22:@56892.4]
    .clock(RetimeWrapper_404_clock),
    .reset(RetimeWrapper_404_reset),
    .io_flow(RetimeWrapper_404_io_flow),
    .io_in(RetimeWrapper_404_io_in),
    .io_out(RetimeWrapper_404_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_405 ( // @[package.scala 93:22:@56900.4]
    .clock(RetimeWrapper_405_clock),
    .reset(RetimeWrapper_405_reset),
    .io_flow(RetimeWrapper_405_io_flow),
    .io_in(RetimeWrapper_405_io_in),
    .io_out(RetimeWrapper_405_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_406 ( // @[package.scala 93:22:@56908.4]
    .clock(RetimeWrapper_406_clock),
    .reset(RetimeWrapper_406_reset),
    .io_flow(RetimeWrapper_406_io_flow),
    .io_in(RetimeWrapper_406_io_in),
    .io_out(RetimeWrapper_406_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_407 ( // @[package.scala 93:22:@56916.4]
    .clock(RetimeWrapper_407_clock),
    .reset(RetimeWrapper_407_reset),
    .io_flow(RetimeWrapper_407_io_flow),
    .io_in(RetimeWrapper_407_io_in),
    .io_out(RetimeWrapper_407_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_408 ( // @[package.scala 93:22:@56924.4]
    .clock(RetimeWrapper_408_clock),
    .reset(RetimeWrapper_408_reset),
    .io_flow(RetimeWrapper_408_io_flow),
    .io_in(RetimeWrapper_408_io_in),
    .io_out(RetimeWrapper_408_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_409 ( // @[package.scala 93:22:@56932.4]
    .clock(RetimeWrapper_409_clock),
    .reset(RetimeWrapper_409_reset),
    .io_flow(RetimeWrapper_409_io_flow),
    .io_in(RetimeWrapper_409_io_in),
    .io_out(RetimeWrapper_409_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_410 ( // @[package.scala 93:22:@56940.4]
    .clock(RetimeWrapper_410_clock),
    .reset(RetimeWrapper_410_reset),
    .io_flow(RetimeWrapper_410_io_flow),
    .io_in(RetimeWrapper_410_io_in),
    .io_out(RetimeWrapper_410_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_411 ( // @[package.scala 93:22:@56948.4]
    .clock(RetimeWrapper_411_clock),
    .reset(RetimeWrapper_411_reset),
    .io_flow(RetimeWrapper_411_io_flow),
    .io_in(RetimeWrapper_411_io_in),
    .io_out(RetimeWrapper_411_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_412 ( // @[package.scala 93:22:@56956.4]
    .clock(RetimeWrapper_412_clock),
    .reset(RetimeWrapper_412_reset),
    .io_flow(RetimeWrapper_412_io_flow),
    .io_in(RetimeWrapper_412_io_in),
    .io_out(RetimeWrapper_412_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_413 ( // @[package.scala 93:22:@56964.4]
    .clock(RetimeWrapper_413_clock),
    .reset(RetimeWrapper_413_reset),
    .io_flow(RetimeWrapper_413_io_flow),
    .io_in(RetimeWrapper_413_io_in),
    .io_out(RetimeWrapper_413_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_414 ( // @[package.scala 93:22:@56972.4]
    .clock(RetimeWrapper_414_clock),
    .reset(RetimeWrapper_414_reset),
    .io_flow(RetimeWrapper_414_io_flow),
    .io_in(RetimeWrapper_414_io_in),
    .io_out(RetimeWrapper_414_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_415 ( // @[package.scala 93:22:@56980.4]
    .clock(RetimeWrapper_415_clock),
    .reset(RetimeWrapper_415_reset),
    .io_flow(RetimeWrapper_415_io_flow),
    .io_in(RetimeWrapper_415_io_in),
    .io_out(RetimeWrapper_415_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_416 ( // @[package.scala 93:22:@56988.4]
    .clock(RetimeWrapper_416_clock),
    .reset(RetimeWrapper_416_reset),
    .io_flow(RetimeWrapper_416_io_flow),
    .io_in(RetimeWrapper_416_io_in),
    .io_out(RetimeWrapper_416_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_417 ( // @[package.scala 93:22:@56996.4]
    .clock(RetimeWrapper_417_clock),
    .reset(RetimeWrapper_417_reset),
    .io_flow(RetimeWrapper_417_io_flow),
    .io_in(RetimeWrapper_417_io_in),
    .io_out(RetimeWrapper_417_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_418 ( // @[package.scala 93:22:@57004.4]
    .clock(RetimeWrapper_418_clock),
    .reset(RetimeWrapper_418_reset),
    .io_flow(RetimeWrapper_418_io_flow),
    .io_in(RetimeWrapper_418_io_in),
    .io_out(RetimeWrapper_418_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_419 ( // @[package.scala 93:22:@57012.4]
    .clock(RetimeWrapper_419_clock),
    .reset(RetimeWrapper_419_reset),
    .io_flow(RetimeWrapper_419_io_flow),
    .io_in(RetimeWrapper_419_io_in),
    .io_out(RetimeWrapper_419_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_420 ( // @[package.scala 93:22:@57100.4]
    .clock(RetimeWrapper_420_clock),
    .reset(RetimeWrapper_420_reset),
    .io_flow(RetimeWrapper_420_io_flow),
    .io_in(RetimeWrapper_420_io_in),
    .io_out(RetimeWrapper_420_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_421 ( // @[package.scala 93:22:@57108.4]
    .clock(RetimeWrapper_421_clock),
    .reset(RetimeWrapper_421_reset),
    .io_flow(RetimeWrapper_421_io_flow),
    .io_in(RetimeWrapper_421_io_in),
    .io_out(RetimeWrapper_421_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_422 ( // @[package.scala 93:22:@57116.4]
    .clock(RetimeWrapper_422_clock),
    .reset(RetimeWrapper_422_reset),
    .io_flow(RetimeWrapper_422_io_flow),
    .io_in(RetimeWrapper_422_io_in),
    .io_out(RetimeWrapper_422_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_423 ( // @[package.scala 93:22:@57124.4]
    .clock(RetimeWrapper_423_clock),
    .reset(RetimeWrapper_423_reset),
    .io_flow(RetimeWrapper_423_io_flow),
    .io_in(RetimeWrapper_423_io_in),
    .io_out(RetimeWrapper_423_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_424 ( // @[package.scala 93:22:@57132.4]
    .clock(RetimeWrapper_424_clock),
    .reset(RetimeWrapper_424_reset),
    .io_flow(RetimeWrapper_424_io_flow),
    .io_in(RetimeWrapper_424_io_in),
    .io_out(RetimeWrapper_424_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_425 ( // @[package.scala 93:22:@57140.4]
    .clock(RetimeWrapper_425_clock),
    .reset(RetimeWrapper_425_reset),
    .io_flow(RetimeWrapper_425_io_flow),
    .io_in(RetimeWrapper_425_io_in),
    .io_out(RetimeWrapper_425_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_426 ( // @[package.scala 93:22:@57148.4]
    .clock(RetimeWrapper_426_clock),
    .reset(RetimeWrapper_426_reset),
    .io_flow(RetimeWrapper_426_io_flow),
    .io_in(RetimeWrapper_426_io_in),
    .io_out(RetimeWrapper_426_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_427 ( // @[package.scala 93:22:@57156.4]
    .clock(RetimeWrapper_427_clock),
    .reset(RetimeWrapper_427_reset),
    .io_flow(RetimeWrapper_427_io_flow),
    .io_in(RetimeWrapper_427_io_in),
    .io_out(RetimeWrapper_427_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_428 ( // @[package.scala 93:22:@57164.4]
    .clock(RetimeWrapper_428_clock),
    .reset(RetimeWrapper_428_reset),
    .io_flow(RetimeWrapper_428_io_flow),
    .io_in(RetimeWrapper_428_io_in),
    .io_out(RetimeWrapper_428_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_429 ( // @[package.scala 93:22:@57172.4]
    .clock(RetimeWrapper_429_clock),
    .reset(RetimeWrapper_429_reset),
    .io_flow(RetimeWrapper_429_io_flow),
    .io_in(RetimeWrapper_429_io_in),
    .io_out(RetimeWrapper_429_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_430 ( // @[package.scala 93:22:@57180.4]
    .clock(RetimeWrapper_430_clock),
    .reset(RetimeWrapper_430_reset),
    .io_flow(RetimeWrapper_430_io_flow),
    .io_in(RetimeWrapper_430_io_in),
    .io_out(RetimeWrapper_430_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_431 ( // @[package.scala 93:22:@57188.4]
    .clock(RetimeWrapper_431_clock),
    .reset(RetimeWrapper_431_reset),
    .io_flow(RetimeWrapper_431_io_flow),
    .io_in(RetimeWrapper_431_io_in),
    .io_out(RetimeWrapper_431_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_432 ( // @[package.scala 93:22:@57196.4]
    .clock(RetimeWrapper_432_clock),
    .reset(RetimeWrapper_432_reset),
    .io_flow(RetimeWrapper_432_io_flow),
    .io_in(RetimeWrapper_432_io_in),
    .io_out(RetimeWrapper_432_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_433 ( // @[package.scala 93:22:@57204.4]
    .clock(RetimeWrapper_433_clock),
    .reset(RetimeWrapper_433_reset),
    .io_flow(RetimeWrapper_433_io_flow),
    .io_in(RetimeWrapper_433_io_in),
    .io_out(RetimeWrapper_433_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_434 ( // @[package.scala 93:22:@57212.4]
    .clock(RetimeWrapper_434_clock),
    .reset(RetimeWrapper_434_reset),
    .io_flow(RetimeWrapper_434_io_flow),
    .io_in(RetimeWrapper_434_io_in),
    .io_out(RetimeWrapper_434_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_435 ( // @[package.scala 93:22:@57220.4]
    .clock(RetimeWrapper_435_clock),
    .reset(RetimeWrapper_435_reset),
    .io_flow(RetimeWrapper_435_io_flow),
    .io_in(RetimeWrapper_435_io_in),
    .io_out(RetimeWrapper_435_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_436 ( // @[package.scala 93:22:@57228.4]
    .clock(RetimeWrapper_436_clock),
    .reset(RetimeWrapper_436_reset),
    .io_flow(RetimeWrapper_436_io_flow),
    .io_in(RetimeWrapper_436_io_in),
    .io_out(RetimeWrapper_436_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_437 ( // @[package.scala 93:22:@57236.4]
    .clock(RetimeWrapper_437_clock),
    .reset(RetimeWrapper_437_reset),
    .io_flow(RetimeWrapper_437_io_flow),
    .io_in(RetimeWrapper_437_io_in),
    .io_out(RetimeWrapper_437_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_438 ( // @[package.scala 93:22:@57244.4]
    .clock(RetimeWrapper_438_clock),
    .reset(RetimeWrapper_438_reset),
    .io_flow(RetimeWrapper_438_io_flow),
    .io_in(RetimeWrapper_438_io_in),
    .io_out(RetimeWrapper_438_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_439 ( // @[package.scala 93:22:@57252.4]
    .clock(RetimeWrapper_439_clock),
    .reset(RetimeWrapper_439_reset),
    .io_flow(RetimeWrapper_439_io_flow),
    .io_in(RetimeWrapper_439_io_in),
    .io_out(RetimeWrapper_439_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_440 ( // @[package.scala 93:22:@57340.4]
    .clock(RetimeWrapper_440_clock),
    .reset(RetimeWrapper_440_reset),
    .io_flow(RetimeWrapper_440_io_flow),
    .io_in(RetimeWrapper_440_io_in),
    .io_out(RetimeWrapper_440_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_441 ( // @[package.scala 93:22:@57348.4]
    .clock(RetimeWrapper_441_clock),
    .reset(RetimeWrapper_441_reset),
    .io_flow(RetimeWrapper_441_io_flow),
    .io_in(RetimeWrapper_441_io_in),
    .io_out(RetimeWrapper_441_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_442 ( // @[package.scala 93:22:@57356.4]
    .clock(RetimeWrapper_442_clock),
    .reset(RetimeWrapper_442_reset),
    .io_flow(RetimeWrapper_442_io_flow),
    .io_in(RetimeWrapper_442_io_in),
    .io_out(RetimeWrapper_442_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_443 ( // @[package.scala 93:22:@57364.4]
    .clock(RetimeWrapper_443_clock),
    .reset(RetimeWrapper_443_reset),
    .io_flow(RetimeWrapper_443_io_flow),
    .io_in(RetimeWrapper_443_io_in),
    .io_out(RetimeWrapper_443_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_444 ( // @[package.scala 93:22:@57372.4]
    .clock(RetimeWrapper_444_clock),
    .reset(RetimeWrapper_444_reset),
    .io_flow(RetimeWrapper_444_io_flow),
    .io_in(RetimeWrapper_444_io_in),
    .io_out(RetimeWrapper_444_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_445 ( // @[package.scala 93:22:@57380.4]
    .clock(RetimeWrapper_445_clock),
    .reset(RetimeWrapper_445_reset),
    .io_flow(RetimeWrapper_445_io_flow),
    .io_in(RetimeWrapper_445_io_in),
    .io_out(RetimeWrapper_445_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_446 ( // @[package.scala 93:22:@57388.4]
    .clock(RetimeWrapper_446_clock),
    .reset(RetimeWrapper_446_reset),
    .io_flow(RetimeWrapper_446_io_flow),
    .io_in(RetimeWrapper_446_io_in),
    .io_out(RetimeWrapper_446_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_447 ( // @[package.scala 93:22:@57396.4]
    .clock(RetimeWrapper_447_clock),
    .reset(RetimeWrapper_447_reset),
    .io_flow(RetimeWrapper_447_io_flow),
    .io_in(RetimeWrapper_447_io_in),
    .io_out(RetimeWrapper_447_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_448 ( // @[package.scala 93:22:@57404.4]
    .clock(RetimeWrapper_448_clock),
    .reset(RetimeWrapper_448_reset),
    .io_flow(RetimeWrapper_448_io_flow),
    .io_in(RetimeWrapper_448_io_in),
    .io_out(RetimeWrapper_448_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_449 ( // @[package.scala 93:22:@57412.4]
    .clock(RetimeWrapper_449_clock),
    .reset(RetimeWrapper_449_reset),
    .io_flow(RetimeWrapper_449_io_flow),
    .io_in(RetimeWrapper_449_io_in),
    .io_out(RetimeWrapper_449_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_450 ( // @[package.scala 93:22:@57420.4]
    .clock(RetimeWrapper_450_clock),
    .reset(RetimeWrapper_450_reset),
    .io_flow(RetimeWrapper_450_io_flow),
    .io_in(RetimeWrapper_450_io_in),
    .io_out(RetimeWrapper_450_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_451 ( // @[package.scala 93:22:@57428.4]
    .clock(RetimeWrapper_451_clock),
    .reset(RetimeWrapper_451_reset),
    .io_flow(RetimeWrapper_451_io_flow),
    .io_in(RetimeWrapper_451_io_in),
    .io_out(RetimeWrapper_451_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_452 ( // @[package.scala 93:22:@57436.4]
    .clock(RetimeWrapper_452_clock),
    .reset(RetimeWrapper_452_reset),
    .io_flow(RetimeWrapper_452_io_flow),
    .io_in(RetimeWrapper_452_io_in),
    .io_out(RetimeWrapper_452_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_453 ( // @[package.scala 93:22:@57444.4]
    .clock(RetimeWrapper_453_clock),
    .reset(RetimeWrapper_453_reset),
    .io_flow(RetimeWrapper_453_io_flow),
    .io_in(RetimeWrapper_453_io_in),
    .io_out(RetimeWrapper_453_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_454 ( // @[package.scala 93:22:@57452.4]
    .clock(RetimeWrapper_454_clock),
    .reset(RetimeWrapper_454_reset),
    .io_flow(RetimeWrapper_454_io_flow),
    .io_in(RetimeWrapper_454_io_in),
    .io_out(RetimeWrapper_454_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_455 ( // @[package.scala 93:22:@57460.4]
    .clock(RetimeWrapper_455_clock),
    .reset(RetimeWrapper_455_reset),
    .io_flow(RetimeWrapper_455_io_flow),
    .io_in(RetimeWrapper_455_io_in),
    .io_out(RetimeWrapper_455_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_456 ( // @[package.scala 93:22:@57468.4]
    .clock(RetimeWrapper_456_clock),
    .reset(RetimeWrapper_456_reset),
    .io_flow(RetimeWrapper_456_io_flow),
    .io_in(RetimeWrapper_456_io_in),
    .io_out(RetimeWrapper_456_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_457 ( // @[package.scala 93:22:@57476.4]
    .clock(RetimeWrapper_457_clock),
    .reset(RetimeWrapper_457_reset),
    .io_flow(RetimeWrapper_457_io_flow),
    .io_in(RetimeWrapper_457_io_in),
    .io_out(RetimeWrapper_457_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_458 ( // @[package.scala 93:22:@57484.4]
    .clock(RetimeWrapper_458_clock),
    .reset(RetimeWrapper_458_reset),
    .io_flow(RetimeWrapper_458_io_flow),
    .io_in(RetimeWrapper_458_io_in),
    .io_out(RetimeWrapper_458_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_459 ( // @[package.scala 93:22:@57492.4]
    .clock(RetimeWrapper_459_clock),
    .reset(RetimeWrapper_459_reset),
    .io_flow(RetimeWrapper_459_io_flow),
    .io_in(RetimeWrapper_459_io_in),
    .io_out(RetimeWrapper_459_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_460 ( // @[package.scala 93:22:@57580.4]
    .clock(RetimeWrapper_460_clock),
    .reset(RetimeWrapper_460_reset),
    .io_flow(RetimeWrapper_460_io_flow),
    .io_in(RetimeWrapper_460_io_in),
    .io_out(RetimeWrapper_460_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_461 ( // @[package.scala 93:22:@57588.4]
    .clock(RetimeWrapper_461_clock),
    .reset(RetimeWrapper_461_reset),
    .io_flow(RetimeWrapper_461_io_flow),
    .io_in(RetimeWrapper_461_io_in),
    .io_out(RetimeWrapper_461_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_462 ( // @[package.scala 93:22:@57596.4]
    .clock(RetimeWrapper_462_clock),
    .reset(RetimeWrapper_462_reset),
    .io_flow(RetimeWrapper_462_io_flow),
    .io_in(RetimeWrapper_462_io_in),
    .io_out(RetimeWrapper_462_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_463 ( // @[package.scala 93:22:@57604.4]
    .clock(RetimeWrapper_463_clock),
    .reset(RetimeWrapper_463_reset),
    .io_flow(RetimeWrapper_463_io_flow),
    .io_in(RetimeWrapper_463_io_in),
    .io_out(RetimeWrapper_463_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_464 ( // @[package.scala 93:22:@57612.4]
    .clock(RetimeWrapper_464_clock),
    .reset(RetimeWrapper_464_reset),
    .io_flow(RetimeWrapper_464_io_flow),
    .io_in(RetimeWrapper_464_io_in),
    .io_out(RetimeWrapper_464_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_465 ( // @[package.scala 93:22:@57620.4]
    .clock(RetimeWrapper_465_clock),
    .reset(RetimeWrapper_465_reset),
    .io_flow(RetimeWrapper_465_io_flow),
    .io_in(RetimeWrapper_465_io_in),
    .io_out(RetimeWrapper_465_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_466 ( // @[package.scala 93:22:@57628.4]
    .clock(RetimeWrapper_466_clock),
    .reset(RetimeWrapper_466_reset),
    .io_flow(RetimeWrapper_466_io_flow),
    .io_in(RetimeWrapper_466_io_in),
    .io_out(RetimeWrapper_466_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_467 ( // @[package.scala 93:22:@57636.4]
    .clock(RetimeWrapper_467_clock),
    .reset(RetimeWrapper_467_reset),
    .io_flow(RetimeWrapper_467_io_flow),
    .io_in(RetimeWrapper_467_io_in),
    .io_out(RetimeWrapper_467_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_468 ( // @[package.scala 93:22:@57644.4]
    .clock(RetimeWrapper_468_clock),
    .reset(RetimeWrapper_468_reset),
    .io_flow(RetimeWrapper_468_io_flow),
    .io_in(RetimeWrapper_468_io_in),
    .io_out(RetimeWrapper_468_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_469 ( // @[package.scala 93:22:@57652.4]
    .clock(RetimeWrapper_469_clock),
    .reset(RetimeWrapper_469_reset),
    .io_flow(RetimeWrapper_469_io_flow),
    .io_in(RetimeWrapper_469_io_in),
    .io_out(RetimeWrapper_469_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_470 ( // @[package.scala 93:22:@57660.4]
    .clock(RetimeWrapper_470_clock),
    .reset(RetimeWrapper_470_reset),
    .io_flow(RetimeWrapper_470_io_flow),
    .io_in(RetimeWrapper_470_io_in),
    .io_out(RetimeWrapper_470_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_471 ( // @[package.scala 93:22:@57668.4]
    .clock(RetimeWrapper_471_clock),
    .reset(RetimeWrapper_471_reset),
    .io_flow(RetimeWrapper_471_io_flow),
    .io_in(RetimeWrapper_471_io_in),
    .io_out(RetimeWrapper_471_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_472 ( // @[package.scala 93:22:@57676.4]
    .clock(RetimeWrapper_472_clock),
    .reset(RetimeWrapper_472_reset),
    .io_flow(RetimeWrapper_472_io_flow),
    .io_in(RetimeWrapper_472_io_in),
    .io_out(RetimeWrapper_472_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_473 ( // @[package.scala 93:22:@57684.4]
    .clock(RetimeWrapper_473_clock),
    .reset(RetimeWrapper_473_reset),
    .io_flow(RetimeWrapper_473_io_flow),
    .io_in(RetimeWrapper_473_io_in),
    .io_out(RetimeWrapper_473_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_474 ( // @[package.scala 93:22:@57692.4]
    .clock(RetimeWrapper_474_clock),
    .reset(RetimeWrapper_474_reset),
    .io_flow(RetimeWrapper_474_io_flow),
    .io_in(RetimeWrapper_474_io_in),
    .io_out(RetimeWrapper_474_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_475 ( // @[package.scala 93:22:@57700.4]
    .clock(RetimeWrapper_475_clock),
    .reset(RetimeWrapper_475_reset),
    .io_flow(RetimeWrapper_475_io_flow),
    .io_in(RetimeWrapper_475_io_in),
    .io_out(RetimeWrapper_475_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_476 ( // @[package.scala 93:22:@57708.4]
    .clock(RetimeWrapper_476_clock),
    .reset(RetimeWrapper_476_reset),
    .io_flow(RetimeWrapper_476_io_flow),
    .io_in(RetimeWrapper_476_io_in),
    .io_out(RetimeWrapper_476_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_477 ( // @[package.scala 93:22:@57716.4]
    .clock(RetimeWrapper_477_clock),
    .reset(RetimeWrapper_477_reset),
    .io_flow(RetimeWrapper_477_io_flow),
    .io_in(RetimeWrapper_477_io_in),
    .io_out(RetimeWrapper_477_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_478 ( // @[package.scala 93:22:@57724.4]
    .clock(RetimeWrapper_478_clock),
    .reset(RetimeWrapper_478_reset),
    .io_flow(RetimeWrapper_478_io_flow),
    .io_in(RetimeWrapper_478_io_in),
    .io_out(RetimeWrapper_478_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_479 ( // @[package.scala 93:22:@57732.4]
    .clock(RetimeWrapper_479_clock),
    .reset(RetimeWrapper_479_reset),
    .io_flow(RetimeWrapper_479_io_flow),
    .io_in(RetimeWrapper_479_io_in),
    .io_out(RetimeWrapper_479_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_480 ( // @[package.scala 93:22:@57820.4]
    .clock(RetimeWrapper_480_clock),
    .reset(RetimeWrapper_480_reset),
    .io_flow(RetimeWrapper_480_io_flow),
    .io_in(RetimeWrapper_480_io_in),
    .io_out(RetimeWrapper_480_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_481 ( // @[package.scala 93:22:@57828.4]
    .clock(RetimeWrapper_481_clock),
    .reset(RetimeWrapper_481_reset),
    .io_flow(RetimeWrapper_481_io_flow),
    .io_in(RetimeWrapper_481_io_in),
    .io_out(RetimeWrapper_481_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_482 ( // @[package.scala 93:22:@57836.4]
    .clock(RetimeWrapper_482_clock),
    .reset(RetimeWrapper_482_reset),
    .io_flow(RetimeWrapper_482_io_flow),
    .io_in(RetimeWrapper_482_io_in),
    .io_out(RetimeWrapper_482_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_483 ( // @[package.scala 93:22:@57844.4]
    .clock(RetimeWrapper_483_clock),
    .reset(RetimeWrapper_483_reset),
    .io_flow(RetimeWrapper_483_io_flow),
    .io_in(RetimeWrapper_483_io_in),
    .io_out(RetimeWrapper_483_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_484 ( // @[package.scala 93:22:@57852.4]
    .clock(RetimeWrapper_484_clock),
    .reset(RetimeWrapper_484_reset),
    .io_flow(RetimeWrapper_484_io_flow),
    .io_in(RetimeWrapper_484_io_in),
    .io_out(RetimeWrapper_484_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_485 ( // @[package.scala 93:22:@57860.4]
    .clock(RetimeWrapper_485_clock),
    .reset(RetimeWrapper_485_reset),
    .io_flow(RetimeWrapper_485_io_flow),
    .io_in(RetimeWrapper_485_io_in),
    .io_out(RetimeWrapper_485_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_486 ( // @[package.scala 93:22:@57868.4]
    .clock(RetimeWrapper_486_clock),
    .reset(RetimeWrapper_486_reset),
    .io_flow(RetimeWrapper_486_io_flow),
    .io_in(RetimeWrapper_486_io_in),
    .io_out(RetimeWrapper_486_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_487 ( // @[package.scala 93:22:@57876.4]
    .clock(RetimeWrapper_487_clock),
    .reset(RetimeWrapper_487_reset),
    .io_flow(RetimeWrapper_487_io_flow),
    .io_in(RetimeWrapper_487_io_in),
    .io_out(RetimeWrapper_487_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_488 ( // @[package.scala 93:22:@57884.4]
    .clock(RetimeWrapper_488_clock),
    .reset(RetimeWrapper_488_reset),
    .io_flow(RetimeWrapper_488_io_flow),
    .io_in(RetimeWrapper_488_io_in),
    .io_out(RetimeWrapper_488_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_489 ( // @[package.scala 93:22:@57892.4]
    .clock(RetimeWrapper_489_clock),
    .reset(RetimeWrapper_489_reset),
    .io_flow(RetimeWrapper_489_io_flow),
    .io_in(RetimeWrapper_489_io_in),
    .io_out(RetimeWrapper_489_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_490 ( // @[package.scala 93:22:@57900.4]
    .clock(RetimeWrapper_490_clock),
    .reset(RetimeWrapper_490_reset),
    .io_flow(RetimeWrapper_490_io_flow),
    .io_in(RetimeWrapper_490_io_in),
    .io_out(RetimeWrapper_490_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_491 ( // @[package.scala 93:22:@57908.4]
    .clock(RetimeWrapper_491_clock),
    .reset(RetimeWrapper_491_reset),
    .io_flow(RetimeWrapper_491_io_flow),
    .io_in(RetimeWrapper_491_io_in),
    .io_out(RetimeWrapper_491_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_492 ( // @[package.scala 93:22:@57916.4]
    .clock(RetimeWrapper_492_clock),
    .reset(RetimeWrapper_492_reset),
    .io_flow(RetimeWrapper_492_io_flow),
    .io_in(RetimeWrapper_492_io_in),
    .io_out(RetimeWrapper_492_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_493 ( // @[package.scala 93:22:@57924.4]
    .clock(RetimeWrapper_493_clock),
    .reset(RetimeWrapper_493_reset),
    .io_flow(RetimeWrapper_493_io_flow),
    .io_in(RetimeWrapper_493_io_in),
    .io_out(RetimeWrapper_493_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_494 ( // @[package.scala 93:22:@57932.4]
    .clock(RetimeWrapper_494_clock),
    .reset(RetimeWrapper_494_reset),
    .io_flow(RetimeWrapper_494_io_flow),
    .io_in(RetimeWrapper_494_io_in),
    .io_out(RetimeWrapper_494_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_495 ( // @[package.scala 93:22:@57940.4]
    .clock(RetimeWrapper_495_clock),
    .reset(RetimeWrapper_495_reset),
    .io_flow(RetimeWrapper_495_io_flow),
    .io_in(RetimeWrapper_495_io_in),
    .io_out(RetimeWrapper_495_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_496 ( // @[package.scala 93:22:@57948.4]
    .clock(RetimeWrapper_496_clock),
    .reset(RetimeWrapper_496_reset),
    .io_flow(RetimeWrapper_496_io_flow),
    .io_in(RetimeWrapper_496_io_in),
    .io_out(RetimeWrapper_496_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_497 ( // @[package.scala 93:22:@57956.4]
    .clock(RetimeWrapper_497_clock),
    .reset(RetimeWrapper_497_reset),
    .io_flow(RetimeWrapper_497_io_flow),
    .io_in(RetimeWrapper_497_io_in),
    .io_out(RetimeWrapper_497_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_498 ( // @[package.scala 93:22:@57964.4]
    .clock(RetimeWrapper_498_clock),
    .reset(RetimeWrapper_498_reset),
    .io_flow(RetimeWrapper_498_io_flow),
    .io_in(RetimeWrapper_498_io_in),
    .io_out(RetimeWrapper_498_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_499 ( // @[package.scala 93:22:@57972.4]
    .clock(RetimeWrapper_499_clock),
    .reset(RetimeWrapper_499_reset),
    .io_flow(RetimeWrapper_499_io_flow),
    .io_in(RetimeWrapper_499_io_in),
    .io_out(RetimeWrapper_499_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_500 ( // @[package.scala 93:22:@58060.4]
    .clock(RetimeWrapper_500_clock),
    .reset(RetimeWrapper_500_reset),
    .io_flow(RetimeWrapper_500_io_flow),
    .io_in(RetimeWrapper_500_io_in),
    .io_out(RetimeWrapper_500_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_501 ( // @[package.scala 93:22:@58068.4]
    .clock(RetimeWrapper_501_clock),
    .reset(RetimeWrapper_501_reset),
    .io_flow(RetimeWrapper_501_io_flow),
    .io_in(RetimeWrapper_501_io_in),
    .io_out(RetimeWrapper_501_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_502 ( // @[package.scala 93:22:@58076.4]
    .clock(RetimeWrapper_502_clock),
    .reset(RetimeWrapper_502_reset),
    .io_flow(RetimeWrapper_502_io_flow),
    .io_in(RetimeWrapper_502_io_in),
    .io_out(RetimeWrapper_502_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_503 ( // @[package.scala 93:22:@58084.4]
    .clock(RetimeWrapper_503_clock),
    .reset(RetimeWrapper_503_reset),
    .io_flow(RetimeWrapper_503_io_flow),
    .io_in(RetimeWrapper_503_io_in),
    .io_out(RetimeWrapper_503_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_504 ( // @[package.scala 93:22:@58092.4]
    .clock(RetimeWrapper_504_clock),
    .reset(RetimeWrapper_504_reset),
    .io_flow(RetimeWrapper_504_io_flow),
    .io_in(RetimeWrapper_504_io_in),
    .io_out(RetimeWrapper_504_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_505 ( // @[package.scala 93:22:@58100.4]
    .clock(RetimeWrapper_505_clock),
    .reset(RetimeWrapper_505_reset),
    .io_flow(RetimeWrapper_505_io_flow),
    .io_in(RetimeWrapper_505_io_in),
    .io_out(RetimeWrapper_505_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_506 ( // @[package.scala 93:22:@58108.4]
    .clock(RetimeWrapper_506_clock),
    .reset(RetimeWrapper_506_reset),
    .io_flow(RetimeWrapper_506_io_flow),
    .io_in(RetimeWrapper_506_io_in),
    .io_out(RetimeWrapper_506_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_507 ( // @[package.scala 93:22:@58116.4]
    .clock(RetimeWrapper_507_clock),
    .reset(RetimeWrapper_507_reset),
    .io_flow(RetimeWrapper_507_io_flow),
    .io_in(RetimeWrapper_507_io_in),
    .io_out(RetimeWrapper_507_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_508 ( // @[package.scala 93:22:@58124.4]
    .clock(RetimeWrapper_508_clock),
    .reset(RetimeWrapper_508_reset),
    .io_flow(RetimeWrapper_508_io_flow),
    .io_in(RetimeWrapper_508_io_in),
    .io_out(RetimeWrapper_508_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_509 ( // @[package.scala 93:22:@58132.4]
    .clock(RetimeWrapper_509_clock),
    .reset(RetimeWrapper_509_reset),
    .io_flow(RetimeWrapper_509_io_flow),
    .io_in(RetimeWrapper_509_io_in),
    .io_out(RetimeWrapper_509_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_510 ( // @[package.scala 93:22:@58140.4]
    .clock(RetimeWrapper_510_clock),
    .reset(RetimeWrapper_510_reset),
    .io_flow(RetimeWrapper_510_io_flow),
    .io_in(RetimeWrapper_510_io_in),
    .io_out(RetimeWrapper_510_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_511 ( // @[package.scala 93:22:@58148.4]
    .clock(RetimeWrapper_511_clock),
    .reset(RetimeWrapper_511_reset),
    .io_flow(RetimeWrapper_511_io_flow),
    .io_in(RetimeWrapper_511_io_in),
    .io_out(RetimeWrapper_511_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_512 ( // @[package.scala 93:22:@58156.4]
    .clock(RetimeWrapper_512_clock),
    .reset(RetimeWrapper_512_reset),
    .io_flow(RetimeWrapper_512_io_flow),
    .io_in(RetimeWrapper_512_io_in),
    .io_out(RetimeWrapper_512_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_513 ( // @[package.scala 93:22:@58164.4]
    .clock(RetimeWrapper_513_clock),
    .reset(RetimeWrapper_513_reset),
    .io_flow(RetimeWrapper_513_io_flow),
    .io_in(RetimeWrapper_513_io_in),
    .io_out(RetimeWrapper_513_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_514 ( // @[package.scala 93:22:@58172.4]
    .clock(RetimeWrapper_514_clock),
    .reset(RetimeWrapper_514_reset),
    .io_flow(RetimeWrapper_514_io_flow),
    .io_in(RetimeWrapper_514_io_in),
    .io_out(RetimeWrapper_514_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_515 ( // @[package.scala 93:22:@58180.4]
    .clock(RetimeWrapper_515_clock),
    .reset(RetimeWrapper_515_reset),
    .io_flow(RetimeWrapper_515_io_flow),
    .io_in(RetimeWrapper_515_io_in),
    .io_out(RetimeWrapper_515_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_516 ( // @[package.scala 93:22:@58188.4]
    .clock(RetimeWrapper_516_clock),
    .reset(RetimeWrapper_516_reset),
    .io_flow(RetimeWrapper_516_io_flow),
    .io_in(RetimeWrapper_516_io_in),
    .io_out(RetimeWrapper_516_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_517 ( // @[package.scala 93:22:@58196.4]
    .clock(RetimeWrapper_517_clock),
    .reset(RetimeWrapper_517_reset),
    .io_flow(RetimeWrapper_517_io_flow),
    .io_in(RetimeWrapper_517_io_in),
    .io_out(RetimeWrapper_517_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_518 ( // @[package.scala 93:22:@58204.4]
    .clock(RetimeWrapper_518_clock),
    .reset(RetimeWrapper_518_reset),
    .io_flow(RetimeWrapper_518_io_flow),
    .io_in(RetimeWrapper_518_io_in),
    .io_out(RetimeWrapper_518_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_519 ( // @[package.scala 93:22:@58212.4]
    .clock(RetimeWrapper_519_clock),
    .reset(RetimeWrapper_519_reset),
    .io_flow(RetimeWrapper_519_io_flow),
    .io_in(RetimeWrapper_519_io_in),
    .io_out(RetimeWrapper_519_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_520 ( // @[package.scala 93:22:@58300.4]
    .clock(RetimeWrapper_520_clock),
    .reset(RetimeWrapper_520_reset),
    .io_flow(RetimeWrapper_520_io_flow),
    .io_in(RetimeWrapper_520_io_in),
    .io_out(RetimeWrapper_520_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_521 ( // @[package.scala 93:22:@58308.4]
    .clock(RetimeWrapper_521_clock),
    .reset(RetimeWrapper_521_reset),
    .io_flow(RetimeWrapper_521_io_flow),
    .io_in(RetimeWrapper_521_io_in),
    .io_out(RetimeWrapper_521_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_522 ( // @[package.scala 93:22:@58316.4]
    .clock(RetimeWrapper_522_clock),
    .reset(RetimeWrapper_522_reset),
    .io_flow(RetimeWrapper_522_io_flow),
    .io_in(RetimeWrapper_522_io_in),
    .io_out(RetimeWrapper_522_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_523 ( // @[package.scala 93:22:@58324.4]
    .clock(RetimeWrapper_523_clock),
    .reset(RetimeWrapper_523_reset),
    .io_flow(RetimeWrapper_523_io_flow),
    .io_in(RetimeWrapper_523_io_in),
    .io_out(RetimeWrapper_523_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_524 ( // @[package.scala 93:22:@58332.4]
    .clock(RetimeWrapper_524_clock),
    .reset(RetimeWrapper_524_reset),
    .io_flow(RetimeWrapper_524_io_flow),
    .io_in(RetimeWrapper_524_io_in),
    .io_out(RetimeWrapper_524_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_525 ( // @[package.scala 93:22:@58340.4]
    .clock(RetimeWrapper_525_clock),
    .reset(RetimeWrapper_525_reset),
    .io_flow(RetimeWrapper_525_io_flow),
    .io_in(RetimeWrapper_525_io_in),
    .io_out(RetimeWrapper_525_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_526 ( // @[package.scala 93:22:@58348.4]
    .clock(RetimeWrapper_526_clock),
    .reset(RetimeWrapper_526_reset),
    .io_flow(RetimeWrapper_526_io_flow),
    .io_in(RetimeWrapper_526_io_in),
    .io_out(RetimeWrapper_526_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_527 ( // @[package.scala 93:22:@58356.4]
    .clock(RetimeWrapper_527_clock),
    .reset(RetimeWrapper_527_reset),
    .io_flow(RetimeWrapper_527_io_flow),
    .io_in(RetimeWrapper_527_io_in),
    .io_out(RetimeWrapper_527_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_528 ( // @[package.scala 93:22:@58364.4]
    .clock(RetimeWrapper_528_clock),
    .reset(RetimeWrapper_528_reset),
    .io_flow(RetimeWrapper_528_io_flow),
    .io_in(RetimeWrapper_528_io_in),
    .io_out(RetimeWrapper_528_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_529 ( // @[package.scala 93:22:@58372.4]
    .clock(RetimeWrapper_529_clock),
    .reset(RetimeWrapper_529_reset),
    .io_flow(RetimeWrapper_529_io_flow),
    .io_in(RetimeWrapper_529_io_in),
    .io_out(RetimeWrapper_529_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_530 ( // @[package.scala 93:22:@58380.4]
    .clock(RetimeWrapper_530_clock),
    .reset(RetimeWrapper_530_reset),
    .io_flow(RetimeWrapper_530_io_flow),
    .io_in(RetimeWrapper_530_io_in),
    .io_out(RetimeWrapper_530_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_531 ( // @[package.scala 93:22:@58388.4]
    .clock(RetimeWrapper_531_clock),
    .reset(RetimeWrapper_531_reset),
    .io_flow(RetimeWrapper_531_io_flow),
    .io_in(RetimeWrapper_531_io_in),
    .io_out(RetimeWrapper_531_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_532 ( // @[package.scala 93:22:@58396.4]
    .clock(RetimeWrapper_532_clock),
    .reset(RetimeWrapper_532_reset),
    .io_flow(RetimeWrapper_532_io_flow),
    .io_in(RetimeWrapper_532_io_in),
    .io_out(RetimeWrapper_532_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_533 ( // @[package.scala 93:22:@58404.4]
    .clock(RetimeWrapper_533_clock),
    .reset(RetimeWrapper_533_reset),
    .io_flow(RetimeWrapper_533_io_flow),
    .io_in(RetimeWrapper_533_io_in),
    .io_out(RetimeWrapper_533_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_534 ( // @[package.scala 93:22:@58412.4]
    .clock(RetimeWrapper_534_clock),
    .reset(RetimeWrapper_534_reset),
    .io_flow(RetimeWrapper_534_io_flow),
    .io_in(RetimeWrapper_534_io_in),
    .io_out(RetimeWrapper_534_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_535 ( // @[package.scala 93:22:@58420.4]
    .clock(RetimeWrapper_535_clock),
    .reset(RetimeWrapper_535_reset),
    .io_flow(RetimeWrapper_535_io_flow),
    .io_in(RetimeWrapper_535_io_in),
    .io_out(RetimeWrapper_535_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_536 ( // @[package.scala 93:22:@58428.4]
    .clock(RetimeWrapper_536_clock),
    .reset(RetimeWrapper_536_reset),
    .io_flow(RetimeWrapper_536_io_flow),
    .io_in(RetimeWrapper_536_io_in),
    .io_out(RetimeWrapper_536_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_537 ( // @[package.scala 93:22:@58436.4]
    .clock(RetimeWrapper_537_clock),
    .reset(RetimeWrapper_537_reset),
    .io_flow(RetimeWrapper_537_io_flow),
    .io_in(RetimeWrapper_537_io_in),
    .io_out(RetimeWrapper_537_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_538 ( // @[package.scala 93:22:@58444.4]
    .clock(RetimeWrapper_538_clock),
    .reset(RetimeWrapper_538_reset),
    .io_flow(RetimeWrapper_538_io_flow),
    .io_in(RetimeWrapper_538_io_in),
    .io_out(RetimeWrapper_538_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_539 ( // @[package.scala 93:22:@58452.4]
    .clock(RetimeWrapper_539_clock),
    .reset(RetimeWrapper_539_reset),
    .io_flow(RetimeWrapper_539_io_flow),
    .io_in(RetimeWrapper_539_io_in),
    .io_out(RetimeWrapper_539_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_540 ( // @[package.scala 93:22:@58540.4]
    .clock(RetimeWrapper_540_clock),
    .reset(RetimeWrapper_540_reset),
    .io_flow(RetimeWrapper_540_io_flow),
    .io_in(RetimeWrapper_540_io_in),
    .io_out(RetimeWrapper_540_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_541 ( // @[package.scala 93:22:@58548.4]
    .clock(RetimeWrapper_541_clock),
    .reset(RetimeWrapper_541_reset),
    .io_flow(RetimeWrapper_541_io_flow),
    .io_in(RetimeWrapper_541_io_in),
    .io_out(RetimeWrapper_541_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_542 ( // @[package.scala 93:22:@58556.4]
    .clock(RetimeWrapper_542_clock),
    .reset(RetimeWrapper_542_reset),
    .io_flow(RetimeWrapper_542_io_flow),
    .io_in(RetimeWrapper_542_io_in),
    .io_out(RetimeWrapper_542_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_543 ( // @[package.scala 93:22:@58564.4]
    .clock(RetimeWrapper_543_clock),
    .reset(RetimeWrapper_543_reset),
    .io_flow(RetimeWrapper_543_io_flow),
    .io_in(RetimeWrapper_543_io_in),
    .io_out(RetimeWrapper_543_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_544 ( // @[package.scala 93:22:@58572.4]
    .clock(RetimeWrapper_544_clock),
    .reset(RetimeWrapper_544_reset),
    .io_flow(RetimeWrapper_544_io_flow),
    .io_in(RetimeWrapper_544_io_in),
    .io_out(RetimeWrapper_544_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_545 ( // @[package.scala 93:22:@58580.4]
    .clock(RetimeWrapper_545_clock),
    .reset(RetimeWrapper_545_reset),
    .io_flow(RetimeWrapper_545_io_flow),
    .io_in(RetimeWrapper_545_io_in),
    .io_out(RetimeWrapper_545_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_546 ( // @[package.scala 93:22:@58588.4]
    .clock(RetimeWrapper_546_clock),
    .reset(RetimeWrapper_546_reset),
    .io_flow(RetimeWrapper_546_io_flow),
    .io_in(RetimeWrapper_546_io_in),
    .io_out(RetimeWrapper_546_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_547 ( // @[package.scala 93:22:@58596.4]
    .clock(RetimeWrapper_547_clock),
    .reset(RetimeWrapper_547_reset),
    .io_flow(RetimeWrapper_547_io_flow),
    .io_in(RetimeWrapper_547_io_in),
    .io_out(RetimeWrapper_547_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_548 ( // @[package.scala 93:22:@58604.4]
    .clock(RetimeWrapper_548_clock),
    .reset(RetimeWrapper_548_reset),
    .io_flow(RetimeWrapper_548_io_flow),
    .io_in(RetimeWrapper_548_io_in),
    .io_out(RetimeWrapper_548_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_549 ( // @[package.scala 93:22:@58612.4]
    .clock(RetimeWrapper_549_clock),
    .reset(RetimeWrapper_549_reset),
    .io_flow(RetimeWrapper_549_io_flow),
    .io_in(RetimeWrapper_549_io_in),
    .io_out(RetimeWrapper_549_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_550 ( // @[package.scala 93:22:@58620.4]
    .clock(RetimeWrapper_550_clock),
    .reset(RetimeWrapper_550_reset),
    .io_flow(RetimeWrapper_550_io_flow),
    .io_in(RetimeWrapper_550_io_in),
    .io_out(RetimeWrapper_550_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_551 ( // @[package.scala 93:22:@58628.4]
    .clock(RetimeWrapper_551_clock),
    .reset(RetimeWrapper_551_reset),
    .io_flow(RetimeWrapper_551_io_flow),
    .io_in(RetimeWrapper_551_io_in),
    .io_out(RetimeWrapper_551_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_552 ( // @[package.scala 93:22:@58636.4]
    .clock(RetimeWrapper_552_clock),
    .reset(RetimeWrapper_552_reset),
    .io_flow(RetimeWrapper_552_io_flow),
    .io_in(RetimeWrapper_552_io_in),
    .io_out(RetimeWrapper_552_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_553 ( // @[package.scala 93:22:@58644.4]
    .clock(RetimeWrapper_553_clock),
    .reset(RetimeWrapper_553_reset),
    .io_flow(RetimeWrapper_553_io_flow),
    .io_in(RetimeWrapper_553_io_in),
    .io_out(RetimeWrapper_553_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_554 ( // @[package.scala 93:22:@58652.4]
    .clock(RetimeWrapper_554_clock),
    .reset(RetimeWrapper_554_reset),
    .io_flow(RetimeWrapper_554_io_flow),
    .io_in(RetimeWrapper_554_io_in),
    .io_out(RetimeWrapper_554_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_555 ( // @[package.scala 93:22:@58660.4]
    .clock(RetimeWrapper_555_clock),
    .reset(RetimeWrapper_555_reset),
    .io_flow(RetimeWrapper_555_io_flow),
    .io_in(RetimeWrapper_555_io_in),
    .io_out(RetimeWrapper_555_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_556 ( // @[package.scala 93:22:@58668.4]
    .clock(RetimeWrapper_556_clock),
    .reset(RetimeWrapper_556_reset),
    .io_flow(RetimeWrapper_556_io_flow),
    .io_in(RetimeWrapper_556_io_in),
    .io_out(RetimeWrapper_556_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_557 ( // @[package.scala 93:22:@58676.4]
    .clock(RetimeWrapper_557_clock),
    .reset(RetimeWrapper_557_reset),
    .io_flow(RetimeWrapper_557_io_flow),
    .io_in(RetimeWrapper_557_io_in),
    .io_out(RetimeWrapper_557_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_558 ( // @[package.scala 93:22:@58684.4]
    .clock(RetimeWrapper_558_clock),
    .reset(RetimeWrapper_558_reset),
    .io_flow(RetimeWrapper_558_io_flow),
    .io_in(RetimeWrapper_558_io_in),
    .io_out(RetimeWrapper_558_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_559 ( // @[package.scala 93:22:@58692.4]
    .clock(RetimeWrapper_559_clock),
    .reset(RetimeWrapper_559_reset),
    .io_flow(RetimeWrapper_559_io_flow),
    .io_in(RetimeWrapper_559_io_in),
    .io_out(RetimeWrapper_559_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_560 ( // @[package.scala 93:22:@58780.4]
    .clock(RetimeWrapper_560_clock),
    .reset(RetimeWrapper_560_reset),
    .io_flow(RetimeWrapper_560_io_flow),
    .io_in(RetimeWrapper_560_io_in),
    .io_out(RetimeWrapper_560_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_561 ( // @[package.scala 93:22:@58788.4]
    .clock(RetimeWrapper_561_clock),
    .reset(RetimeWrapper_561_reset),
    .io_flow(RetimeWrapper_561_io_flow),
    .io_in(RetimeWrapper_561_io_in),
    .io_out(RetimeWrapper_561_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_562 ( // @[package.scala 93:22:@58796.4]
    .clock(RetimeWrapper_562_clock),
    .reset(RetimeWrapper_562_reset),
    .io_flow(RetimeWrapper_562_io_flow),
    .io_in(RetimeWrapper_562_io_in),
    .io_out(RetimeWrapper_562_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_563 ( // @[package.scala 93:22:@58804.4]
    .clock(RetimeWrapper_563_clock),
    .reset(RetimeWrapper_563_reset),
    .io_flow(RetimeWrapper_563_io_flow),
    .io_in(RetimeWrapper_563_io_in),
    .io_out(RetimeWrapper_563_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_564 ( // @[package.scala 93:22:@58812.4]
    .clock(RetimeWrapper_564_clock),
    .reset(RetimeWrapper_564_reset),
    .io_flow(RetimeWrapper_564_io_flow),
    .io_in(RetimeWrapper_564_io_in),
    .io_out(RetimeWrapper_564_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_565 ( // @[package.scala 93:22:@58820.4]
    .clock(RetimeWrapper_565_clock),
    .reset(RetimeWrapper_565_reset),
    .io_flow(RetimeWrapper_565_io_flow),
    .io_in(RetimeWrapper_565_io_in),
    .io_out(RetimeWrapper_565_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_566 ( // @[package.scala 93:22:@58828.4]
    .clock(RetimeWrapper_566_clock),
    .reset(RetimeWrapper_566_reset),
    .io_flow(RetimeWrapper_566_io_flow),
    .io_in(RetimeWrapper_566_io_in),
    .io_out(RetimeWrapper_566_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_567 ( // @[package.scala 93:22:@58836.4]
    .clock(RetimeWrapper_567_clock),
    .reset(RetimeWrapper_567_reset),
    .io_flow(RetimeWrapper_567_io_flow),
    .io_in(RetimeWrapper_567_io_in),
    .io_out(RetimeWrapper_567_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_568 ( // @[package.scala 93:22:@58844.4]
    .clock(RetimeWrapper_568_clock),
    .reset(RetimeWrapper_568_reset),
    .io_flow(RetimeWrapper_568_io_flow),
    .io_in(RetimeWrapper_568_io_in),
    .io_out(RetimeWrapper_568_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_569 ( // @[package.scala 93:22:@58852.4]
    .clock(RetimeWrapper_569_clock),
    .reset(RetimeWrapper_569_reset),
    .io_flow(RetimeWrapper_569_io_flow),
    .io_in(RetimeWrapper_569_io_in),
    .io_out(RetimeWrapper_569_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_570 ( // @[package.scala 93:22:@58860.4]
    .clock(RetimeWrapper_570_clock),
    .reset(RetimeWrapper_570_reset),
    .io_flow(RetimeWrapper_570_io_flow),
    .io_in(RetimeWrapper_570_io_in),
    .io_out(RetimeWrapper_570_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_571 ( // @[package.scala 93:22:@58868.4]
    .clock(RetimeWrapper_571_clock),
    .reset(RetimeWrapper_571_reset),
    .io_flow(RetimeWrapper_571_io_flow),
    .io_in(RetimeWrapper_571_io_in),
    .io_out(RetimeWrapper_571_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_572 ( // @[package.scala 93:22:@58876.4]
    .clock(RetimeWrapper_572_clock),
    .reset(RetimeWrapper_572_reset),
    .io_flow(RetimeWrapper_572_io_flow),
    .io_in(RetimeWrapper_572_io_in),
    .io_out(RetimeWrapper_572_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_573 ( // @[package.scala 93:22:@58884.4]
    .clock(RetimeWrapper_573_clock),
    .reset(RetimeWrapper_573_reset),
    .io_flow(RetimeWrapper_573_io_flow),
    .io_in(RetimeWrapper_573_io_in),
    .io_out(RetimeWrapper_573_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_574 ( // @[package.scala 93:22:@58892.4]
    .clock(RetimeWrapper_574_clock),
    .reset(RetimeWrapper_574_reset),
    .io_flow(RetimeWrapper_574_io_flow),
    .io_in(RetimeWrapper_574_io_in),
    .io_out(RetimeWrapper_574_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_575 ( // @[package.scala 93:22:@58900.4]
    .clock(RetimeWrapper_575_clock),
    .reset(RetimeWrapper_575_reset),
    .io_flow(RetimeWrapper_575_io_flow),
    .io_in(RetimeWrapper_575_io_in),
    .io_out(RetimeWrapper_575_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_576 ( // @[package.scala 93:22:@58908.4]
    .clock(RetimeWrapper_576_clock),
    .reset(RetimeWrapper_576_reset),
    .io_flow(RetimeWrapper_576_io_flow),
    .io_in(RetimeWrapper_576_io_in),
    .io_out(RetimeWrapper_576_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_577 ( // @[package.scala 93:22:@58916.4]
    .clock(RetimeWrapper_577_clock),
    .reset(RetimeWrapper_577_reset),
    .io_flow(RetimeWrapper_577_io_flow),
    .io_in(RetimeWrapper_577_io_in),
    .io_out(RetimeWrapper_577_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_578 ( // @[package.scala 93:22:@58924.4]
    .clock(RetimeWrapper_578_clock),
    .reset(RetimeWrapper_578_reset),
    .io_flow(RetimeWrapper_578_io_flow),
    .io_in(RetimeWrapper_578_io_in),
    .io_out(RetimeWrapper_578_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_579 ( // @[package.scala 93:22:@58932.4]
    .clock(RetimeWrapper_579_clock),
    .reset(RetimeWrapper_579_reset),
    .io_flow(RetimeWrapper_579_io_flow),
    .io_in(RetimeWrapper_579_io_in),
    .io_out(RetimeWrapper_579_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_580 ( // @[package.scala 93:22:@59020.4]
    .clock(RetimeWrapper_580_clock),
    .reset(RetimeWrapper_580_reset),
    .io_flow(RetimeWrapper_580_io_flow),
    .io_in(RetimeWrapper_580_io_in),
    .io_out(RetimeWrapper_580_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_581 ( // @[package.scala 93:22:@59028.4]
    .clock(RetimeWrapper_581_clock),
    .reset(RetimeWrapper_581_reset),
    .io_flow(RetimeWrapper_581_io_flow),
    .io_in(RetimeWrapper_581_io_in),
    .io_out(RetimeWrapper_581_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_582 ( // @[package.scala 93:22:@59036.4]
    .clock(RetimeWrapper_582_clock),
    .reset(RetimeWrapper_582_reset),
    .io_flow(RetimeWrapper_582_io_flow),
    .io_in(RetimeWrapper_582_io_in),
    .io_out(RetimeWrapper_582_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_583 ( // @[package.scala 93:22:@59044.4]
    .clock(RetimeWrapper_583_clock),
    .reset(RetimeWrapper_583_reset),
    .io_flow(RetimeWrapper_583_io_flow),
    .io_in(RetimeWrapper_583_io_in),
    .io_out(RetimeWrapper_583_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_584 ( // @[package.scala 93:22:@59052.4]
    .clock(RetimeWrapper_584_clock),
    .reset(RetimeWrapper_584_reset),
    .io_flow(RetimeWrapper_584_io_flow),
    .io_in(RetimeWrapper_584_io_in),
    .io_out(RetimeWrapper_584_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_585 ( // @[package.scala 93:22:@59060.4]
    .clock(RetimeWrapper_585_clock),
    .reset(RetimeWrapper_585_reset),
    .io_flow(RetimeWrapper_585_io_flow),
    .io_in(RetimeWrapper_585_io_in),
    .io_out(RetimeWrapper_585_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_586 ( // @[package.scala 93:22:@59068.4]
    .clock(RetimeWrapper_586_clock),
    .reset(RetimeWrapper_586_reset),
    .io_flow(RetimeWrapper_586_io_flow),
    .io_in(RetimeWrapper_586_io_in),
    .io_out(RetimeWrapper_586_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_587 ( // @[package.scala 93:22:@59076.4]
    .clock(RetimeWrapper_587_clock),
    .reset(RetimeWrapper_587_reset),
    .io_flow(RetimeWrapper_587_io_flow),
    .io_in(RetimeWrapper_587_io_in),
    .io_out(RetimeWrapper_587_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_588 ( // @[package.scala 93:22:@59084.4]
    .clock(RetimeWrapper_588_clock),
    .reset(RetimeWrapper_588_reset),
    .io_flow(RetimeWrapper_588_io_flow),
    .io_in(RetimeWrapper_588_io_in),
    .io_out(RetimeWrapper_588_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_589 ( // @[package.scala 93:22:@59092.4]
    .clock(RetimeWrapper_589_clock),
    .reset(RetimeWrapper_589_reset),
    .io_flow(RetimeWrapper_589_io_flow),
    .io_in(RetimeWrapper_589_io_in),
    .io_out(RetimeWrapper_589_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_590 ( // @[package.scala 93:22:@59100.4]
    .clock(RetimeWrapper_590_clock),
    .reset(RetimeWrapper_590_reset),
    .io_flow(RetimeWrapper_590_io_flow),
    .io_in(RetimeWrapper_590_io_in),
    .io_out(RetimeWrapper_590_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_591 ( // @[package.scala 93:22:@59108.4]
    .clock(RetimeWrapper_591_clock),
    .reset(RetimeWrapper_591_reset),
    .io_flow(RetimeWrapper_591_io_flow),
    .io_in(RetimeWrapper_591_io_in),
    .io_out(RetimeWrapper_591_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_592 ( // @[package.scala 93:22:@59116.4]
    .clock(RetimeWrapper_592_clock),
    .reset(RetimeWrapper_592_reset),
    .io_flow(RetimeWrapper_592_io_flow),
    .io_in(RetimeWrapper_592_io_in),
    .io_out(RetimeWrapper_592_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_593 ( // @[package.scala 93:22:@59124.4]
    .clock(RetimeWrapper_593_clock),
    .reset(RetimeWrapper_593_reset),
    .io_flow(RetimeWrapper_593_io_flow),
    .io_in(RetimeWrapper_593_io_in),
    .io_out(RetimeWrapper_593_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_594 ( // @[package.scala 93:22:@59132.4]
    .clock(RetimeWrapper_594_clock),
    .reset(RetimeWrapper_594_reset),
    .io_flow(RetimeWrapper_594_io_flow),
    .io_in(RetimeWrapper_594_io_in),
    .io_out(RetimeWrapper_594_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_595 ( // @[package.scala 93:22:@59140.4]
    .clock(RetimeWrapper_595_clock),
    .reset(RetimeWrapper_595_reset),
    .io_flow(RetimeWrapper_595_io_flow),
    .io_in(RetimeWrapper_595_io_in),
    .io_out(RetimeWrapper_595_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_596 ( // @[package.scala 93:22:@59148.4]
    .clock(RetimeWrapper_596_clock),
    .reset(RetimeWrapper_596_reset),
    .io_flow(RetimeWrapper_596_io_flow),
    .io_in(RetimeWrapper_596_io_in),
    .io_out(RetimeWrapper_596_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_597 ( // @[package.scala 93:22:@59156.4]
    .clock(RetimeWrapper_597_clock),
    .reset(RetimeWrapper_597_reset),
    .io_flow(RetimeWrapper_597_io_flow),
    .io_in(RetimeWrapper_597_io_in),
    .io_out(RetimeWrapper_597_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_598 ( // @[package.scala 93:22:@59164.4]
    .clock(RetimeWrapper_598_clock),
    .reset(RetimeWrapper_598_reset),
    .io_flow(RetimeWrapper_598_io_flow),
    .io_in(RetimeWrapper_598_io_in),
    .io_out(RetimeWrapper_598_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_599 ( // @[package.scala 93:22:@59172.4]
    .clock(RetimeWrapper_599_clock),
    .reset(RetimeWrapper_599_reset),
    .io_flow(RetimeWrapper_599_io_flow),
    .io_in(RetimeWrapper_599_io_in),
    .io_out(RetimeWrapper_599_io_out)
  );
  assign _T_1212 = io_wPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@44959.4]
  assign _T_1214 = io_wPort_4_banks_1 == 4'h0; // @[MemPrimitives.scala 82:210:@44960.4]
  assign _T_1215 = _T_1212 & _T_1214; // @[MemPrimitives.scala 82:228:@44961.4]
  assign _T_1216 = io_wPort_4_en_0 & _T_1215; // @[MemPrimitives.scala 83:102:@44962.4]
  assign _T_1218 = io_wPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@44963.4]
  assign _T_1220 = io_wPort_5_banks_1 == 4'h0; // @[MemPrimitives.scala 82:210:@44964.4]
  assign _T_1221 = _T_1218 & _T_1220; // @[MemPrimitives.scala 82:228:@44965.4]
  assign _T_1222 = io_wPort_5_en_0 & _T_1221; // @[MemPrimitives.scala 83:102:@44966.4]
  assign _T_1224 = io_wPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@44967.4]
  assign _T_1226 = io_wPort_6_banks_1 == 4'h0; // @[MemPrimitives.scala 82:210:@44968.4]
  assign _T_1227 = _T_1224 & _T_1226; // @[MemPrimitives.scala 82:228:@44969.4]
  assign _T_1228 = io_wPort_6_en_0 & _T_1227; // @[MemPrimitives.scala 83:102:@44970.4]
  assign _T_1230 = io_wPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@44971.4]
  assign _T_1232 = io_wPort_7_banks_1 == 4'h0; // @[MemPrimitives.scala 82:210:@44972.4]
  assign _T_1233 = _T_1230 & _T_1232; // @[MemPrimitives.scala 82:228:@44973.4]
  assign _T_1234 = io_wPort_7_en_0 & _T_1233; // @[MemPrimitives.scala 83:102:@44974.4]
  assign _T_1236 = {_T_1216,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@44976.4]
  assign _T_1238 = {_T_1222,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@44978.4]
  assign _T_1240 = {_T_1228,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@44980.4]
  assign _T_1242 = {_T_1234,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@44982.4]
  assign _T_1243 = _T_1228 ? _T_1240 : _T_1242; // @[Mux.scala 31:69:@44983.4]
  assign _T_1244 = _T_1222 ? _T_1238 : _T_1243; // @[Mux.scala 31:69:@44984.4]
  assign _T_1245 = _T_1216 ? _T_1236 : _T_1244; // @[Mux.scala 31:69:@44985.4]
  assign _T_1250 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@44992.4]
  assign _T_1252 = io_wPort_0_banks_1 == 4'h1; // @[MemPrimitives.scala 82:210:@44993.4]
  assign _T_1253 = _T_1250 & _T_1252; // @[MemPrimitives.scala 82:228:@44994.4]
  assign _T_1254 = io_wPort_0_en_0 & _T_1253; // @[MemPrimitives.scala 83:102:@44995.4]
  assign _T_1256 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@44996.4]
  assign _T_1258 = io_wPort_1_banks_1 == 4'h1; // @[MemPrimitives.scala 82:210:@44997.4]
  assign _T_1259 = _T_1256 & _T_1258; // @[MemPrimitives.scala 82:228:@44998.4]
  assign _T_1260 = io_wPort_1_en_0 & _T_1259; // @[MemPrimitives.scala 83:102:@44999.4]
  assign _T_1262 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@45000.4]
  assign _T_1264 = io_wPort_2_banks_1 == 4'h1; // @[MemPrimitives.scala 82:210:@45001.4]
  assign _T_1265 = _T_1262 & _T_1264; // @[MemPrimitives.scala 82:228:@45002.4]
  assign _T_1266 = io_wPort_2_en_0 & _T_1265; // @[MemPrimitives.scala 83:102:@45003.4]
  assign _T_1268 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@45004.4]
  assign _T_1270 = io_wPort_3_banks_1 == 4'h1; // @[MemPrimitives.scala 82:210:@45005.4]
  assign _T_1271 = _T_1268 & _T_1270; // @[MemPrimitives.scala 82:228:@45006.4]
  assign _T_1272 = io_wPort_3_en_0 & _T_1271; // @[MemPrimitives.scala 83:102:@45007.4]
  assign _T_1274 = {_T_1254,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45009.4]
  assign _T_1276 = {_T_1260,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45011.4]
  assign _T_1278 = {_T_1266,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45013.4]
  assign _T_1280 = {_T_1272,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45015.4]
  assign _T_1281 = _T_1266 ? _T_1278 : _T_1280; // @[Mux.scala 31:69:@45016.4]
  assign _T_1282 = _T_1260 ? _T_1276 : _T_1281; // @[Mux.scala 31:69:@45017.4]
  assign _T_1283 = _T_1254 ? _T_1274 : _T_1282; // @[Mux.scala 31:69:@45018.4]
  assign _T_1290 = io_wPort_4_banks_1 == 4'h2; // @[MemPrimitives.scala 82:210:@45026.4]
  assign _T_1291 = _T_1212 & _T_1290; // @[MemPrimitives.scala 82:228:@45027.4]
  assign _T_1292 = io_wPort_4_en_0 & _T_1291; // @[MemPrimitives.scala 83:102:@45028.4]
  assign _T_1296 = io_wPort_5_banks_1 == 4'h2; // @[MemPrimitives.scala 82:210:@45030.4]
  assign _T_1297 = _T_1218 & _T_1296; // @[MemPrimitives.scala 82:228:@45031.4]
  assign _T_1298 = io_wPort_5_en_0 & _T_1297; // @[MemPrimitives.scala 83:102:@45032.4]
  assign _T_1302 = io_wPort_6_banks_1 == 4'h2; // @[MemPrimitives.scala 82:210:@45034.4]
  assign _T_1303 = _T_1224 & _T_1302; // @[MemPrimitives.scala 82:228:@45035.4]
  assign _T_1304 = io_wPort_6_en_0 & _T_1303; // @[MemPrimitives.scala 83:102:@45036.4]
  assign _T_1308 = io_wPort_7_banks_1 == 4'h2; // @[MemPrimitives.scala 82:210:@45038.4]
  assign _T_1309 = _T_1230 & _T_1308; // @[MemPrimitives.scala 82:228:@45039.4]
  assign _T_1310 = io_wPort_7_en_0 & _T_1309; // @[MemPrimitives.scala 83:102:@45040.4]
  assign _T_1312 = {_T_1292,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45042.4]
  assign _T_1314 = {_T_1298,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45044.4]
  assign _T_1316 = {_T_1304,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45046.4]
  assign _T_1318 = {_T_1310,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45048.4]
  assign _T_1319 = _T_1304 ? _T_1316 : _T_1318; // @[Mux.scala 31:69:@45049.4]
  assign _T_1320 = _T_1298 ? _T_1314 : _T_1319; // @[Mux.scala 31:69:@45050.4]
  assign _T_1321 = _T_1292 ? _T_1312 : _T_1320; // @[Mux.scala 31:69:@45051.4]
  assign _T_1328 = io_wPort_0_banks_1 == 4'h3; // @[MemPrimitives.scala 82:210:@45059.4]
  assign _T_1329 = _T_1250 & _T_1328; // @[MemPrimitives.scala 82:228:@45060.4]
  assign _T_1330 = io_wPort_0_en_0 & _T_1329; // @[MemPrimitives.scala 83:102:@45061.4]
  assign _T_1334 = io_wPort_1_banks_1 == 4'h3; // @[MemPrimitives.scala 82:210:@45063.4]
  assign _T_1335 = _T_1256 & _T_1334; // @[MemPrimitives.scala 82:228:@45064.4]
  assign _T_1336 = io_wPort_1_en_0 & _T_1335; // @[MemPrimitives.scala 83:102:@45065.4]
  assign _T_1340 = io_wPort_2_banks_1 == 4'h3; // @[MemPrimitives.scala 82:210:@45067.4]
  assign _T_1341 = _T_1262 & _T_1340; // @[MemPrimitives.scala 82:228:@45068.4]
  assign _T_1342 = io_wPort_2_en_0 & _T_1341; // @[MemPrimitives.scala 83:102:@45069.4]
  assign _T_1346 = io_wPort_3_banks_1 == 4'h3; // @[MemPrimitives.scala 82:210:@45071.4]
  assign _T_1347 = _T_1268 & _T_1346; // @[MemPrimitives.scala 82:228:@45072.4]
  assign _T_1348 = io_wPort_3_en_0 & _T_1347; // @[MemPrimitives.scala 83:102:@45073.4]
  assign _T_1350 = {_T_1330,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45075.4]
  assign _T_1352 = {_T_1336,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45077.4]
  assign _T_1354 = {_T_1342,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45079.4]
  assign _T_1356 = {_T_1348,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45081.4]
  assign _T_1357 = _T_1342 ? _T_1354 : _T_1356; // @[Mux.scala 31:69:@45082.4]
  assign _T_1358 = _T_1336 ? _T_1352 : _T_1357; // @[Mux.scala 31:69:@45083.4]
  assign _T_1359 = _T_1330 ? _T_1350 : _T_1358; // @[Mux.scala 31:69:@45084.4]
  assign _T_1366 = io_wPort_4_banks_1 == 4'h4; // @[MemPrimitives.scala 82:210:@45092.4]
  assign _T_1367 = _T_1212 & _T_1366; // @[MemPrimitives.scala 82:228:@45093.4]
  assign _T_1368 = io_wPort_4_en_0 & _T_1367; // @[MemPrimitives.scala 83:102:@45094.4]
  assign _T_1372 = io_wPort_5_banks_1 == 4'h4; // @[MemPrimitives.scala 82:210:@45096.4]
  assign _T_1373 = _T_1218 & _T_1372; // @[MemPrimitives.scala 82:228:@45097.4]
  assign _T_1374 = io_wPort_5_en_0 & _T_1373; // @[MemPrimitives.scala 83:102:@45098.4]
  assign _T_1378 = io_wPort_6_banks_1 == 4'h4; // @[MemPrimitives.scala 82:210:@45100.4]
  assign _T_1379 = _T_1224 & _T_1378; // @[MemPrimitives.scala 82:228:@45101.4]
  assign _T_1380 = io_wPort_6_en_0 & _T_1379; // @[MemPrimitives.scala 83:102:@45102.4]
  assign _T_1384 = io_wPort_7_banks_1 == 4'h4; // @[MemPrimitives.scala 82:210:@45104.4]
  assign _T_1385 = _T_1230 & _T_1384; // @[MemPrimitives.scala 82:228:@45105.4]
  assign _T_1386 = io_wPort_7_en_0 & _T_1385; // @[MemPrimitives.scala 83:102:@45106.4]
  assign _T_1388 = {_T_1368,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45108.4]
  assign _T_1390 = {_T_1374,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45110.4]
  assign _T_1392 = {_T_1380,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45112.4]
  assign _T_1394 = {_T_1386,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45114.4]
  assign _T_1395 = _T_1380 ? _T_1392 : _T_1394; // @[Mux.scala 31:69:@45115.4]
  assign _T_1396 = _T_1374 ? _T_1390 : _T_1395; // @[Mux.scala 31:69:@45116.4]
  assign _T_1397 = _T_1368 ? _T_1388 : _T_1396; // @[Mux.scala 31:69:@45117.4]
  assign _T_1404 = io_wPort_0_banks_1 == 4'h5; // @[MemPrimitives.scala 82:210:@45125.4]
  assign _T_1405 = _T_1250 & _T_1404; // @[MemPrimitives.scala 82:228:@45126.4]
  assign _T_1406 = io_wPort_0_en_0 & _T_1405; // @[MemPrimitives.scala 83:102:@45127.4]
  assign _T_1410 = io_wPort_1_banks_1 == 4'h5; // @[MemPrimitives.scala 82:210:@45129.4]
  assign _T_1411 = _T_1256 & _T_1410; // @[MemPrimitives.scala 82:228:@45130.4]
  assign _T_1412 = io_wPort_1_en_0 & _T_1411; // @[MemPrimitives.scala 83:102:@45131.4]
  assign _T_1416 = io_wPort_2_banks_1 == 4'h5; // @[MemPrimitives.scala 82:210:@45133.4]
  assign _T_1417 = _T_1262 & _T_1416; // @[MemPrimitives.scala 82:228:@45134.4]
  assign _T_1418 = io_wPort_2_en_0 & _T_1417; // @[MemPrimitives.scala 83:102:@45135.4]
  assign _T_1422 = io_wPort_3_banks_1 == 4'h5; // @[MemPrimitives.scala 82:210:@45137.4]
  assign _T_1423 = _T_1268 & _T_1422; // @[MemPrimitives.scala 82:228:@45138.4]
  assign _T_1424 = io_wPort_3_en_0 & _T_1423; // @[MemPrimitives.scala 83:102:@45139.4]
  assign _T_1426 = {_T_1406,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45141.4]
  assign _T_1428 = {_T_1412,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45143.4]
  assign _T_1430 = {_T_1418,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45145.4]
  assign _T_1432 = {_T_1424,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45147.4]
  assign _T_1433 = _T_1418 ? _T_1430 : _T_1432; // @[Mux.scala 31:69:@45148.4]
  assign _T_1434 = _T_1412 ? _T_1428 : _T_1433; // @[Mux.scala 31:69:@45149.4]
  assign _T_1435 = _T_1406 ? _T_1426 : _T_1434; // @[Mux.scala 31:69:@45150.4]
  assign _T_1442 = io_wPort_4_banks_1 == 4'h6; // @[MemPrimitives.scala 82:210:@45158.4]
  assign _T_1443 = _T_1212 & _T_1442; // @[MemPrimitives.scala 82:228:@45159.4]
  assign _T_1444 = io_wPort_4_en_0 & _T_1443; // @[MemPrimitives.scala 83:102:@45160.4]
  assign _T_1448 = io_wPort_5_banks_1 == 4'h6; // @[MemPrimitives.scala 82:210:@45162.4]
  assign _T_1449 = _T_1218 & _T_1448; // @[MemPrimitives.scala 82:228:@45163.4]
  assign _T_1450 = io_wPort_5_en_0 & _T_1449; // @[MemPrimitives.scala 83:102:@45164.4]
  assign _T_1454 = io_wPort_6_banks_1 == 4'h6; // @[MemPrimitives.scala 82:210:@45166.4]
  assign _T_1455 = _T_1224 & _T_1454; // @[MemPrimitives.scala 82:228:@45167.4]
  assign _T_1456 = io_wPort_6_en_0 & _T_1455; // @[MemPrimitives.scala 83:102:@45168.4]
  assign _T_1460 = io_wPort_7_banks_1 == 4'h6; // @[MemPrimitives.scala 82:210:@45170.4]
  assign _T_1461 = _T_1230 & _T_1460; // @[MemPrimitives.scala 82:228:@45171.4]
  assign _T_1462 = io_wPort_7_en_0 & _T_1461; // @[MemPrimitives.scala 83:102:@45172.4]
  assign _T_1464 = {_T_1444,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45174.4]
  assign _T_1466 = {_T_1450,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45176.4]
  assign _T_1468 = {_T_1456,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45178.4]
  assign _T_1470 = {_T_1462,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45180.4]
  assign _T_1471 = _T_1456 ? _T_1468 : _T_1470; // @[Mux.scala 31:69:@45181.4]
  assign _T_1472 = _T_1450 ? _T_1466 : _T_1471; // @[Mux.scala 31:69:@45182.4]
  assign _T_1473 = _T_1444 ? _T_1464 : _T_1472; // @[Mux.scala 31:69:@45183.4]
  assign _T_1480 = io_wPort_0_banks_1 == 4'h7; // @[MemPrimitives.scala 82:210:@45191.4]
  assign _T_1481 = _T_1250 & _T_1480; // @[MemPrimitives.scala 82:228:@45192.4]
  assign _T_1482 = io_wPort_0_en_0 & _T_1481; // @[MemPrimitives.scala 83:102:@45193.4]
  assign _T_1486 = io_wPort_1_banks_1 == 4'h7; // @[MemPrimitives.scala 82:210:@45195.4]
  assign _T_1487 = _T_1256 & _T_1486; // @[MemPrimitives.scala 82:228:@45196.4]
  assign _T_1488 = io_wPort_1_en_0 & _T_1487; // @[MemPrimitives.scala 83:102:@45197.4]
  assign _T_1492 = io_wPort_2_banks_1 == 4'h7; // @[MemPrimitives.scala 82:210:@45199.4]
  assign _T_1493 = _T_1262 & _T_1492; // @[MemPrimitives.scala 82:228:@45200.4]
  assign _T_1494 = io_wPort_2_en_0 & _T_1493; // @[MemPrimitives.scala 83:102:@45201.4]
  assign _T_1498 = io_wPort_3_banks_1 == 4'h7; // @[MemPrimitives.scala 82:210:@45203.4]
  assign _T_1499 = _T_1268 & _T_1498; // @[MemPrimitives.scala 82:228:@45204.4]
  assign _T_1500 = io_wPort_3_en_0 & _T_1499; // @[MemPrimitives.scala 83:102:@45205.4]
  assign _T_1502 = {_T_1482,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45207.4]
  assign _T_1504 = {_T_1488,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45209.4]
  assign _T_1506 = {_T_1494,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45211.4]
  assign _T_1508 = {_T_1500,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45213.4]
  assign _T_1509 = _T_1494 ? _T_1506 : _T_1508; // @[Mux.scala 31:69:@45214.4]
  assign _T_1510 = _T_1488 ? _T_1504 : _T_1509; // @[Mux.scala 31:69:@45215.4]
  assign _T_1511 = _T_1482 ? _T_1502 : _T_1510; // @[Mux.scala 31:69:@45216.4]
  assign _T_1518 = io_wPort_4_banks_1 == 4'h8; // @[MemPrimitives.scala 82:210:@45224.4]
  assign _T_1519 = _T_1212 & _T_1518; // @[MemPrimitives.scala 82:228:@45225.4]
  assign _T_1520 = io_wPort_4_en_0 & _T_1519; // @[MemPrimitives.scala 83:102:@45226.4]
  assign _T_1524 = io_wPort_5_banks_1 == 4'h8; // @[MemPrimitives.scala 82:210:@45228.4]
  assign _T_1525 = _T_1218 & _T_1524; // @[MemPrimitives.scala 82:228:@45229.4]
  assign _T_1526 = io_wPort_5_en_0 & _T_1525; // @[MemPrimitives.scala 83:102:@45230.4]
  assign _T_1530 = io_wPort_6_banks_1 == 4'h8; // @[MemPrimitives.scala 82:210:@45232.4]
  assign _T_1531 = _T_1224 & _T_1530; // @[MemPrimitives.scala 82:228:@45233.4]
  assign _T_1532 = io_wPort_6_en_0 & _T_1531; // @[MemPrimitives.scala 83:102:@45234.4]
  assign _T_1536 = io_wPort_7_banks_1 == 4'h8; // @[MemPrimitives.scala 82:210:@45236.4]
  assign _T_1537 = _T_1230 & _T_1536; // @[MemPrimitives.scala 82:228:@45237.4]
  assign _T_1538 = io_wPort_7_en_0 & _T_1537; // @[MemPrimitives.scala 83:102:@45238.4]
  assign _T_1540 = {_T_1520,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45240.4]
  assign _T_1542 = {_T_1526,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45242.4]
  assign _T_1544 = {_T_1532,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45244.4]
  assign _T_1546 = {_T_1538,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45246.4]
  assign _T_1547 = _T_1532 ? _T_1544 : _T_1546; // @[Mux.scala 31:69:@45247.4]
  assign _T_1548 = _T_1526 ? _T_1542 : _T_1547; // @[Mux.scala 31:69:@45248.4]
  assign _T_1549 = _T_1520 ? _T_1540 : _T_1548; // @[Mux.scala 31:69:@45249.4]
  assign _T_1556 = io_wPort_0_banks_1 == 4'h9; // @[MemPrimitives.scala 82:210:@45257.4]
  assign _T_1557 = _T_1250 & _T_1556; // @[MemPrimitives.scala 82:228:@45258.4]
  assign _T_1558 = io_wPort_0_en_0 & _T_1557; // @[MemPrimitives.scala 83:102:@45259.4]
  assign _T_1562 = io_wPort_1_banks_1 == 4'h9; // @[MemPrimitives.scala 82:210:@45261.4]
  assign _T_1563 = _T_1256 & _T_1562; // @[MemPrimitives.scala 82:228:@45262.4]
  assign _T_1564 = io_wPort_1_en_0 & _T_1563; // @[MemPrimitives.scala 83:102:@45263.4]
  assign _T_1568 = io_wPort_2_banks_1 == 4'h9; // @[MemPrimitives.scala 82:210:@45265.4]
  assign _T_1569 = _T_1262 & _T_1568; // @[MemPrimitives.scala 82:228:@45266.4]
  assign _T_1570 = io_wPort_2_en_0 & _T_1569; // @[MemPrimitives.scala 83:102:@45267.4]
  assign _T_1574 = io_wPort_3_banks_1 == 4'h9; // @[MemPrimitives.scala 82:210:@45269.4]
  assign _T_1575 = _T_1268 & _T_1574; // @[MemPrimitives.scala 82:228:@45270.4]
  assign _T_1576 = io_wPort_3_en_0 & _T_1575; // @[MemPrimitives.scala 83:102:@45271.4]
  assign _T_1578 = {_T_1558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45273.4]
  assign _T_1580 = {_T_1564,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45275.4]
  assign _T_1582 = {_T_1570,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45277.4]
  assign _T_1584 = {_T_1576,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45279.4]
  assign _T_1585 = _T_1570 ? _T_1582 : _T_1584; // @[Mux.scala 31:69:@45280.4]
  assign _T_1586 = _T_1564 ? _T_1580 : _T_1585; // @[Mux.scala 31:69:@45281.4]
  assign _T_1587 = _T_1558 ? _T_1578 : _T_1586; // @[Mux.scala 31:69:@45282.4]
  assign _T_1592 = io_wPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45289.4]
  assign _T_1595 = _T_1592 & _T_1214; // @[MemPrimitives.scala 82:228:@45291.4]
  assign _T_1596 = io_wPort_4_en_0 & _T_1595; // @[MemPrimitives.scala 83:102:@45292.4]
  assign _T_1598 = io_wPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45293.4]
  assign _T_1601 = _T_1598 & _T_1220; // @[MemPrimitives.scala 82:228:@45295.4]
  assign _T_1602 = io_wPort_5_en_0 & _T_1601; // @[MemPrimitives.scala 83:102:@45296.4]
  assign _T_1604 = io_wPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45297.4]
  assign _T_1607 = _T_1604 & _T_1226; // @[MemPrimitives.scala 82:228:@45299.4]
  assign _T_1608 = io_wPort_6_en_0 & _T_1607; // @[MemPrimitives.scala 83:102:@45300.4]
  assign _T_1610 = io_wPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45301.4]
  assign _T_1613 = _T_1610 & _T_1232; // @[MemPrimitives.scala 82:228:@45303.4]
  assign _T_1614 = io_wPort_7_en_0 & _T_1613; // @[MemPrimitives.scala 83:102:@45304.4]
  assign _T_1616 = {_T_1596,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45306.4]
  assign _T_1618 = {_T_1602,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45308.4]
  assign _T_1620 = {_T_1608,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45310.4]
  assign _T_1622 = {_T_1614,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45312.4]
  assign _T_1623 = _T_1608 ? _T_1620 : _T_1622; // @[Mux.scala 31:69:@45313.4]
  assign _T_1624 = _T_1602 ? _T_1618 : _T_1623; // @[Mux.scala 31:69:@45314.4]
  assign _T_1625 = _T_1596 ? _T_1616 : _T_1624; // @[Mux.scala 31:69:@45315.4]
  assign _T_1630 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45322.4]
  assign _T_1633 = _T_1630 & _T_1252; // @[MemPrimitives.scala 82:228:@45324.4]
  assign _T_1634 = io_wPort_0_en_0 & _T_1633; // @[MemPrimitives.scala 83:102:@45325.4]
  assign _T_1636 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45326.4]
  assign _T_1639 = _T_1636 & _T_1258; // @[MemPrimitives.scala 82:228:@45328.4]
  assign _T_1640 = io_wPort_1_en_0 & _T_1639; // @[MemPrimitives.scala 83:102:@45329.4]
  assign _T_1642 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45330.4]
  assign _T_1645 = _T_1642 & _T_1264; // @[MemPrimitives.scala 82:228:@45332.4]
  assign _T_1646 = io_wPort_2_en_0 & _T_1645; // @[MemPrimitives.scala 83:102:@45333.4]
  assign _T_1648 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@45334.4]
  assign _T_1651 = _T_1648 & _T_1270; // @[MemPrimitives.scala 82:228:@45336.4]
  assign _T_1652 = io_wPort_3_en_0 & _T_1651; // @[MemPrimitives.scala 83:102:@45337.4]
  assign _T_1654 = {_T_1634,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45339.4]
  assign _T_1656 = {_T_1640,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45341.4]
  assign _T_1658 = {_T_1646,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45343.4]
  assign _T_1660 = {_T_1652,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45345.4]
  assign _T_1661 = _T_1646 ? _T_1658 : _T_1660; // @[Mux.scala 31:69:@45346.4]
  assign _T_1662 = _T_1640 ? _T_1656 : _T_1661; // @[Mux.scala 31:69:@45347.4]
  assign _T_1663 = _T_1634 ? _T_1654 : _T_1662; // @[Mux.scala 31:69:@45348.4]
  assign _T_1671 = _T_1592 & _T_1290; // @[MemPrimitives.scala 82:228:@45357.4]
  assign _T_1672 = io_wPort_4_en_0 & _T_1671; // @[MemPrimitives.scala 83:102:@45358.4]
  assign _T_1677 = _T_1598 & _T_1296; // @[MemPrimitives.scala 82:228:@45361.4]
  assign _T_1678 = io_wPort_5_en_0 & _T_1677; // @[MemPrimitives.scala 83:102:@45362.4]
  assign _T_1683 = _T_1604 & _T_1302; // @[MemPrimitives.scala 82:228:@45365.4]
  assign _T_1684 = io_wPort_6_en_0 & _T_1683; // @[MemPrimitives.scala 83:102:@45366.4]
  assign _T_1689 = _T_1610 & _T_1308; // @[MemPrimitives.scala 82:228:@45369.4]
  assign _T_1690 = io_wPort_7_en_0 & _T_1689; // @[MemPrimitives.scala 83:102:@45370.4]
  assign _T_1692 = {_T_1672,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45372.4]
  assign _T_1694 = {_T_1678,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45374.4]
  assign _T_1696 = {_T_1684,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45376.4]
  assign _T_1698 = {_T_1690,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45378.4]
  assign _T_1699 = _T_1684 ? _T_1696 : _T_1698; // @[Mux.scala 31:69:@45379.4]
  assign _T_1700 = _T_1678 ? _T_1694 : _T_1699; // @[Mux.scala 31:69:@45380.4]
  assign _T_1701 = _T_1672 ? _T_1692 : _T_1700; // @[Mux.scala 31:69:@45381.4]
  assign _T_1709 = _T_1630 & _T_1328; // @[MemPrimitives.scala 82:228:@45390.4]
  assign _T_1710 = io_wPort_0_en_0 & _T_1709; // @[MemPrimitives.scala 83:102:@45391.4]
  assign _T_1715 = _T_1636 & _T_1334; // @[MemPrimitives.scala 82:228:@45394.4]
  assign _T_1716 = io_wPort_1_en_0 & _T_1715; // @[MemPrimitives.scala 83:102:@45395.4]
  assign _T_1721 = _T_1642 & _T_1340; // @[MemPrimitives.scala 82:228:@45398.4]
  assign _T_1722 = io_wPort_2_en_0 & _T_1721; // @[MemPrimitives.scala 83:102:@45399.4]
  assign _T_1727 = _T_1648 & _T_1346; // @[MemPrimitives.scala 82:228:@45402.4]
  assign _T_1728 = io_wPort_3_en_0 & _T_1727; // @[MemPrimitives.scala 83:102:@45403.4]
  assign _T_1730 = {_T_1710,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45405.4]
  assign _T_1732 = {_T_1716,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45407.4]
  assign _T_1734 = {_T_1722,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45409.4]
  assign _T_1736 = {_T_1728,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45411.4]
  assign _T_1737 = _T_1722 ? _T_1734 : _T_1736; // @[Mux.scala 31:69:@45412.4]
  assign _T_1738 = _T_1716 ? _T_1732 : _T_1737; // @[Mux.scala 31:69:@45413.4]
  assign _T_1739 = _T_1710 ? _T_1730 : _T_1738; // @[Mux.scala 31:69:@45414.4]
  assign _T_1747 = _T_1592 & _T_1366; // @[MemPrimitives.scala 82:228:@45423.4]
  assign _T_1748 = io_wPort_4_en_0 & _T_1747; // @[MemPrimitives.scala 83:102:@45424.4]
  assign _T_1753 = _T_1598 & _T_1372; // @[MemPrimitives.scala 82:228:@45427.4]
  assign _T_1754 = io_wPort_5_en_0 & _T_1753; // @[MemPrimitives.scala 83:102:@45428.4]
  assign _T_1759 = _T_1604 & _T_1378; // @[MemPrimitives.scala 82:228:@45431.4]
  assign _T_1760 = io_wPort_6_en_0 & _T_1759; // @[MemPrimitives.scala 83:102:@45432.4]
  assign _T_1765 = _T_1610 & _T_1384; // @[MemPrimitives.scala 82:228:@45435.4]
  assign _T_1766 = io_wPort_7_en_0 & _T_1765; // @[MemPrimitives.scala 83:102:@45436.4]
  assign _T_1768 = {_T_1748,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45438.4]
  assign _T_1770 = {_T_1754,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45440.4]
  assign _T_1772 = {_T_1760,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45442.4]
  assign _T_1774 = {_T_1766,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45444.4]
  assign _T_1775 = _T_1760 ? _T_1772 : _T_1774; // @[Mux.scala 31:69:@45445.4]
  assign _T_1776 = _T_1754 ? _T_1770 : _T_1775; // @[Mux.scala 31:69:@45446.4]
  assign _T_1777 = _T_1748 ? _T_1768 : _T_1776; // @[Mux.scala 31:69:@45447.4]
  assign _T_1785 = _T_1630 & _T_1404; // @[MemPrimitives.scala 82:228:@45456.4]
  assign _T_1786 = io_wPort_0_en_0 & _T_1785; // @[MemPrimitives.scala 83:102:@45457.4]
  assign _T_1791 = _T_1636 & _T_1410; // @[MemPrimitives.scala 82:228:@45460.4]
  assign _T_1792 = io_wPort_1_en_0 & _T_1791; // @[MemPrimitives.scala 83:102:@45461.4]
  assign _T_1797 = _T_1642 & _T_1416; // @[MemPrimitives.scala 82:228:@45464.4]
  assign _T_1798 = io_wPort_2_en_0 & _T_1797; // @[MemPrimitives.scala 83:102:@45465.4]
  assign _T_1803 = _T_1648 & _T_1422; // @[MemPrimitives.scala 82:228:@45468.4]
  assign _T_1804 = io_wPort_3_en_0 & _T_1803; // @[MemPrimitives.scala 83:102:@45469.4]
  assign _T_1806 = {_T_1786,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45471.4]
  assign _T_1808 = {_T_1792,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45473.4]
  assign _T_1810 = {_T_1798,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45475.4]
  assign _T_1812 = {_T_1804,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45477.4]
  assign _T_1813 = _T_1798 ? _T_1810 : _T_1812; // @[Mux.scala 31:69:@45478.4]
  assign _T_1814 = _T_1792 ? _T_1808 : _T_1813; // @[Mux.scala 31:69:@45479.4]
  assign _T_1815 = _T_1786 ? _T_1806 : _T_1814; // @[Mux.scala 31:69:@45480.4]
  assign _T_1823 = _T_1592 & _T_1442; // @[MemPrimitives.scala 82:228:@45489.4]
  assign _T_1824 = io_wPort_4_en_0 & _T_1823; // @[MemPrimitives.scala 83:102:@45490.4]
  assign _T_1829 = _T_1598 & _T_1448; // @[MemPrimitives.scala 82:228:@45493.4]
  assign _T_1830 = io_wPort_5_en_0 & _T_1829; // @[MemPrimitives.scala 83:102:@45494.4]
  assign _T_1835 = _T_1604 & _T_1454; // @[MemPrimitives.scala 82:228:@45497.4]
  assign _T_1836 = io_wPort_6_en_0 & _T_1835; // @[MemPrimitives.scala 83:102:@45498.4]
  assign _T_1841 = _T_1610 & _T_1460; // @[MemPrimitives.scala 82:228:@45501.4]
  assign _T_1842 = io_wPort_7_en_0 & _T_1841; // @[MemPrimitives.scala 83:102:@45502.4]
  assign _T_1844 = {_T_1824,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45504.4]
  assign _T_1846 = {_T_1830,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45506.4]
  assign _T_1848 = {_T_1836,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45508.4]
  assign _T_1850 = {_T_1842,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45510.4]
  assign _T_1851 = _T_1836 ? _T_1848 : _T_1850; // @[Mux.scala 31:69:@45511.4]
  assign _T_1852 = _T_1830 ? _T_1846 : _T_1851; // @[Mux.scala 31:69:@45512.4]
  assign _T_1853 = _T_1824 ? _T_1844 : _T_1852; // @[Mux.scala 31:69:@45513.4]
  assign _T_1861 = _T_1630 & _T_1480; // @[MemPrimitives.scala 82:228:@45522.4]
  assign _T_1862 = io_wPort_0_en_0 & _T_1861; // @[MemPrimitives.scala 83:102:@45523.4]
  assign _T_1867 = _T_1636 & _T_1486; // @[MemPrimitives.scala 82:228:@45526.4]
  assign _T_1868 = io_wPort_1_en_0 & _T_1867; // @[MemPrimitives.scala 83:102:@45527.4]
  assign _T_1873 = _T_1642 & _T_1492; // @[MemPrimitives.scala 82:228:@45530.4]
  assign _T_1874 = io_wPort_2_en_0 & _T_1873; // @[MemPrimitives.scala 83:102:@45531.4]
  assign _T_1879 = _T_1648 & _T_1498; // @[MemPrimitives.scala 82:228:@45534.4]
  assign _T_1880 = io_wPort_3_en_0 & _T_1879; // @[MemPrimitives.scala 83:102:@45535.4]
  assign _T_1882 = {_T_1862,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45537.4]
  assign _T_1884 = {_T_1868,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45539.4]
  assign _T_1886 = {_T_1874,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45541.4]
  assign _T_1888 = {_T_1880,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45543.4]
  assign _T_1889 = _T_1874 ? _T_1886 : _T_1888; // @[Mux.scala 31:69:@45544.4]
  assign _T_1890 = _T_1868 ? _T_1884 : _T_1889; // @[Mux.scala 31:69:@45545.4]
  assign _T_1891 = _T_1862 ? _T_1882 : _T_1890; // @[Mux.scala 31:69:@45546.4]
  assign _T_1899 = _T_1592 & _T_1518; // @[MemPrimitives.scala 82:228:@45555.4]
  assign _T_1900 = io_wPort_4_en_0 & _T_1899; // @[MemPrimitives.scala 83:102:@45556.4]
  assign _T_1905 = _T_1598 & _T_1524; // @[MemPrimitives.scala 82:228:@45559.4]
  assign _T_1906 = io_wPort_5_en_0 & _T_1905; // @[MemPrimitives.scala 83:102:@45560.4]
  assign _T_1911 = _T_1604 & _T_1530; // @[MemPrimitives.scala 82:228:@45563.4]
  assign _T_1912 = io_wPort_6_en_0 & _T_1911; // @[MemPrimitives.scala 83:102:@45564.4]
  assign _T_1917 = _T_1610 & _T_1536; // @[MemPrimitives.scala 82:228:@45567.4]
  assign _T_1918 = io_wPort_7_en_0 & _T_1917; // @[MemPrimitives.scala 83:102:@45568.4]
  assign _T_1920 = {_T_1900,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45570.4]
  assign _T_1922 = {_T_1906,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45572.4]
  assign _T_1924 = {_T_1912,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45574.4]
  assign _T_1926 = {_T_1918,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45576.4]
  assign _T_1927 = _T_1912 ? _T_1924 : _T_1926; // @[Mux.scala 31:69:@45577.4]
  assign _T_1928 = _T_1906 ? _T_1922 : _T_1927; // @[Mux.scala 31:69:@45578.4]
  assign _T_1929 = _T_1900 ? _T_1920 : _T_1928; // @[Mux.scala 31:69:@45579.4]
  assign _T_1937 = _T_1630 & _T_1556; // @[MemPrimitives.scala 82:228:@45588.4]
  assign _T_1938 = io_wPort_0_en_0 & _T_1937; // @[MemPrimitives.scala 83:102:@45589.4]
  assign _T_1943 = _T_1636 & _T_1562; // @[MemPrimitives.scala 82:228:@45592.4]
  assign _T_1944 = io_wPort_1_en_0 & _T_1943; // @[MemPrimitives.scala 83:102:@45593.4]
  assign _T_1949 = _T_1642 & _T_1568; // @[MemPrimitives.scala 82:228:@45596.4]
  assign _T_1950 = io_wPort_2_en_0 & _T_1949; // @[MemPrimitives.scala 83:102:@45597.4]
  assign _T_1955 = _T_1648 & _T_1574; // @[MemPrimitives.scala 82:228:@45600.4]
  assign _T_1956 = io_wPort_3_en_0 & _T_1955; // @[MemPrimitives.scala 83:102:@45601.4]
  assign _T_1958 = {_T_1938,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45603.4]
  assign _T_1960 = {_T_1944,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45605.4]
  assign _T_1962 = {_T_1950,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45607.4]
  assign _T_1964 = {_T_1956,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45609.4]
  assign _T_1965 = _T_1950 ? _T_1962 : _T_1964; // @[Mux.scala 31:69:@45610.4]
  assign _T_1966 = _T_1944 ? _T_1960 : _T_1965; // @[Mux.scala 31:69:@45611.4]
  assign _T_1967 = _T_1938 ? _T_1958 : _T_1966; // @[Mux.scala 31:69:@45612.4]
  assign _T_1972 = io_wPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45619.4]
  assign _T_1975 = _T_1972 & _T_1214; // @[MemPrimitives.scala 82:228:@45621.4]
  assign _T_1976 = io_wPort_4_en_0 & _T_1975; // @[MemPrimitives.scala 83:102:@45622.4]
  assign _T_1978 = io_wPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45623.4]
  assign _T_1981 = _T_1978 & _T_1220; // @[MemPrimitives.scala 82:228:@45625.4]
  assign _T_1982 = io_wPort_5_en_0 & _T_1981; // @[MemPrimitives.scala 83:102:@45626.4]
  assign _T_1984 = io_wPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45627.4]
  assign _T_1987 = _T_1984 & _T_1226; // @[MemPrimitives.scala 82:228:@45629.4]
  assign _T_1988 = io_wPort_6_en_0 & _T_1987; // @[MemPrimitives.scala 83:102:@45630.4]
  assign _T_1990 = io_wPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45631.4]
  assign _T_1993 = _T_1990 & _T_1232; // @[MemPrimitives.scala 82:228:@45633.4]
  assign _T_1994 = io_wPort_7_en_0 & _T_1993; // @[MemPrimitives.scala 83:102:@45634.4]
  assign _T_1996 = {_T_1976,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45636.4]
  assign _T_1998 = {_T_1982,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45638.4]
  assign _T_2000 = {_T_1988,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45640.4]
  assign _T_2002 = {_T_1994,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45642.4]
  assign _T_2003 = _T_1988 ? _T_2000 : _T_2002; // @[Mux.scala 31:69:@45643.4]
  assign _T_2004 = _T_1982 ? _T_1998 : _T_2003; // @[Mux.scala 31:69:@45644.4]
  assign _T_2005 = _T_1976 ? _T_1996 : _T_2004; // @[Mux.scala 31:69:@45645.4]
  assign _T_2010 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45652.4]
  assign _T_2013 = _T_2010 & _T_1252; // @[MemPrimitives.scala 82:228:@45654.4]
  assign _T_2014 = io_wPort_0_en_0 & _T_2013; // @[MemPrimitives.scala 83:102:@45655.4]
  assign _T_2016 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45656.4]
  assign _T_2019 = _T_2016 & _T_1258; // @[MemPrimitives.scala 82:228:@45658.4]
  assign _T_2020 = io_wPort_1_en_0 & _T_2019; // @[MemPrimitives.scala 83:102:@45659.4]
  assign _T_2022 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45660.4]
  assign _T_2025 = _T_2022 & _T_1264; // @[MemPrimitives.scala 82:228:@45662.4]
  assign _T_2026 = io_wPort_2_en_0 & _T_2025; // @[MemPrimitives.scala 83:102:@45663.4]
  assign _T_2028 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@45664.4]
  assign _T_2031 = _T_2028 & _T_1270; // @[MemPrimitives.scala 82:228:@45666.4]
  assign _T_2032 = io_wPort_3_en_0 & _T_2031; // @[MemPrimitives.scala 83:102:@45667.4]
  assign _T_2034 = {_T_2014,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45669.4]
  assign _T_2036 = {_T_2020,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45671.4]
  assign _T_2038 = {_T_2026,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45673.4]
  assign _T_2040 = {_T_2032,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45675.4]
  assign _T_2041 = _T_2026 ? _T_2038 : _T_2040; // @[Mux.scala 31:69:@45676.4]
  assign _T_2042 = _T_2020 ? _T_2036 : _T_2041; // @[Mux.scala 31:69:@45677.4]
  assign _T_2043 = _T_2014 ? _T_2034 : _T_2042; // @[Mux.scala 31:69:@45678.4]
  assign _T_2051 = _T_1972 & _T_1290; // @[MemPrimitives.scala 82:228:@45687.4]
  assign _T_2052 = io_wPort_4_en_0 & _T_2051; // @[MemPrimitives.scala 83:102:@45688.4]
  assign _T_2057 = _T_1978 & _T_1296; // @[MemPrimitives.scala 82:228:@45691.4]
  assign _T_2058 = io_wPort_5_en_0 & _T_2057; // @[MemPrimitives.scala 83:102:@45692.4]
  assign _T_2063 = _T_1984 & _T_1302; // @[MemPrimitives.scala 82:228:@45695.4]
  assign _T_2064 = io_wPort_6_en_0 & _T_2063; // @[MemPrimitives.scala 83:102:@45696.4]
  assign _T_2069 = _T_1990 & _T_1308; // @[MemPrimitives.scala 82:228:@45699.4]
  assign _T_2070 = io_wPort_7_en_0 & _T_2069; // @[MemPrimitives.scala 83:102:@45700.4]
  assign _T_2072 = {_T_2052,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45702.4]
  assign _T_2074 = {_T_2058,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45704.4]
  assign _T_2076 = {_T_2064,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45706.4]
  assign _T_2078 = {_T_2070,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45708.4]
  assign _T_2079 = _T_2064 ? _T_2076 : _T_2078; // @[Mux.scala 31:69:@45709.4]
  assign _T_2080 = _T_2058 ? _T_2074 : _T_2079; // @[Mux.scala 31:69:@45710.4]
  assign _T_2081 = _T_2052 ? _T_2072 : _T_2080; // @[Mux.scala 31:69:@45711.4]
  assign _T_2089 = _T_2010 & _T_1328; // @[MemPrimitives.scala 82:228:@45720.4]
  assign _T_2090 = io_wPort_0_en_0 & _T_2089; // @[MemPrimitives.scala 83:102:@45721.4]
  assign _T_2095 = _T_2016 & _T_1334; // @[MemPrimitives.scala 82:228:@45724.4]
  assign _T_2096 = io_wPort_1_en_0 & _T_2095; // @[MemPrimitives.scala 83:102:@45725.4]
  assign _T_2101 = _T_2022 & _T_1340; // @[MemPrimitives.scala 82:228:@45728.4]
  assign _T_2102 = io_wPort_2_en_0 & _T_2101; // @[MemPrimitives.scala 83:102:@45729.4]
  assign _T_2107 = _T_2028 & _T_1346; // @[MemPrimitives.scala 82:228:@45732.4]
  assign _T_2108 = io_wPort_3_en_0 & _T_2107; // @[MemPrimitives.scala 83:102:@45733.4]
  assign _T_2110 = {_T_2090,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45735.4]
  assign _T_2112 = {_T_2096,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45737.4]
  assign _T_2114 = {_T_2102,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45739.4]
  assign _T_2116 = {_T_2108,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45741.4]
  assign _T_2117 = _T_2102 ? _T_2114 : _T_2116; // @[Mux.scala 31:69:@45742.4]
  assign _T_2118 = _T_2096 ? _T_2112 : _T_2117; // @[Mux.scala 31:69:@45743.4]
  assign _T_2119 = _T_2090 ? _T_2110 : _T_2118; // @[Mux.scala 31:69:@45744.4]
  assign _T_2127 = _T_1972 & _T_1366; // @[MemPrimitives.scala 82:228:@45753.4]
  assign _T_2128 = io_wPort_4_en_0 & _T_2127; // @[MemPrimitives.scala 83:102:@45754.4]
  assign _T_2133 = _T_1978 & _T_1372; // @[MemPrimitives.scala 82:228:@45757.4]
  assign _T_2134 = io_wPort_5_en_0 & _T_2133; // @[MemPrimitives.scala 83:102:@45758.4]
  assign _T_2139 = _T_1984 & _T_1378; // @[MemPrimitives.scala 82:228:@45761.4]
  assign _T_2140 = io_wPort_6_en_0 & _T_2139; // @[MemPrimitives.scala 83:102:@45762.4]
  assign _T_2145 = _T_1990 & _T_1384; // @[MemPrimitives.scala 82:228:@45765.4]
  assign _T_2146 = io_wPort_7_en_0 & _T_2145; // @[MemPrimitives.scala 83:102:@45766.4]
  assign _T_2148 = {_T_2128,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45768.4]
  assign _T_2150 = {_T_2134,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45770.4]
  assign _T_2152 = {_T_2140,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45772.4]
  assign _T_2154 = {_T_2146,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45774.4]
  assign _T_2155 = _T_2140 ? _T_2152 : _T_2154; // @[Mux.scala 31:69:@45775.4]
  assign _T_2156 = _T_2134 ? _T_2150 : _T_2155; // @[Mux.scala 31:69:@45776.4]
  assign _T_2157 = _T_2128 ? _T_2148 : _T_2156; // @[Mux.scala 31:69:@45777.4]
  assign _T_2165 = _T_2010 & _T_1404; // @[MemPrimitives.scala 82:228:@45786.4]
  assign _T_2166 = io_wPort_0_en_0 & _T_2165; // @[MemPrimitives.scala 83:102:@45787.4]
  assign _T_2171 = _T_2016 & _T_1410; // @[MemPrimitives.scala 82:228:@45790.4]
  assign _T_2172 = io_wPort_1_en_0 & _T_2171; // @[MemPrimitives.scala 83:102:@45791.4]
  assign _T_2177 = _T_2022 & _T_1416; // @[MemPrimitives.scala 82:228:@45794.4]
  assign _T_2178 = io_wPort_2_en_0 & _T_2177; // @[MemPrimitives.scala 83:102:@45795.4]
  assign _T_2183 = _T_2028 & _T_1422; // @[MemPrimitives.scala 82:228:@45798.4]
  assign _T_2184 = io_wPort_3_en_0 & _T_2183; // @[MemPrimitives.scala 83:102:@45799.4]
  assign _T_2186 = {_T_2166,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45801.4]
  assign _T_2188 = {_T_2172,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45803.4]
  assign _T_2190 = {_T_2178,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45805.4]
  assign _T_2192 = {_T_2184,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45807.4]
  assign _T_2193 = _T_2178 ? _T_2190 : _T_2192; // @[Mux.scala 31:69:@45808.4]
  assign _T_2194 = _T_2172 ? _T_2188 : _T_2193; // @[Mux.scala 31:69:@45809.4]
  assign _T_2195 = _T_2166 ? _T_2186 : _T_2194; // @[Mux.scala 31:69:@45810.4]
  assign _T_2203 = _T_1972 & _T_1442; // @[MemPrimitives.scala 82:228:@45819.4]
  assign _T_2204 = io_wPort_4_en_0 & _T_2203; // @[MemPrimitives.scala 83:102:@45820.4]
  assign _T_2209 = _T_1978 & _T_1448; // @[MemPrimitives.scala 82:228:@45823.4]
  assign _T_2210 = io_wPort_5_en_0 & _T_2209; // @[MemPrimitives.scala 83:102:@45824.4]
  assign _T_2215 = _T_1984 & _T_1454; // @[MemPrimitives.scala 82:228:@45827.4]
  assign _T_2216 = io_wPort_6_en_0 & _T_2215; // @[MemPrimitives.scala 83:102:@45828.4]
  assign _T_2221 = _T_1990 & _T_1460; // @[MemPrimitives.scala 82:228:@45831.4]
  assign _T_2222 = io_wPort_7_en_0 & _T_2221; // @[MemPrimitives.scala 83:102:@45832.4]
  assign _T_2224 = {_T_2204,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45834.4]
  assign _T_2226 = {_T_2210,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45836.4]
  assign _T_2228 = {_T_2216,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45838.4]
  assign _T_2230 = {_T_2222,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45840.4]
  assign _T_2231 = _T_2216 ? _T_2228 : _T_2230; // @[Mux.scala 31:69:@45841.4]
  assign _T_2232 = _T_2210 ? _T_2226 : _T_2231; // @[Mux.scala 31:69:@45842.4]
  assign _T_2233 = _T_2204 ? _T_2224 : _T_2232; // @[Mux.scala 31:69:@45843.4]
  assign _T_2241 = _T_2010 & _T_1480; // @[MemPrimitives.scala 82:228:@45852.4]
  assign _T_2242 = io_wPort_0_en_0 & _T_2241; // @[MemPrimitives.scala 83:102:@45853.4]
  assign _T_2247 = _T_2016 & _T_1486; // @[MemPrimitives.scala 82:228:@45856.4]
  assign _T_2248 = io_wPort_1_en_0 & _T_2247; // @[MemPrimitives.scala 83:102:@45857.4]
  assign _T_2253 = _T_2022 & _T_1492; // @[MemPrimitives.scala 82:228:@45860.4]
  assign _T_2254 = io_wPort_2_en_0 & _T_2253; // @[MemPrimitives.scala 83:102:@45861.4]
  assign _T_2259 = _T_2028 & _T_1498; // @[MemPrimitives.scala 82:228:@45864.4]
  assign _T_2260 = io_wPort_3_en_0 & _T_2259; // @[MemPrimitives.scala 83:102:@45865.4]
  assign _T_2262 = {_T_2242,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45867.4]
  assign _T_2264 = {_T_2248,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45869.4]
  assign _T_2266 = {_T_2254,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45871.4]
  assign _T_2268 = {_T_2260,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45873.4]
  assign _T_2269 = _T_2254 ? _T_2266 : _T_2268; // @[Mux.scala 31:69:@45874.4]
  assign _T_2270 = _T_2248 ? _T_2264 : _T_2269; // @[Mux.scala 31:69:@45875.4]
  assign _T_2271 = _T_2242 ? _T_2262 : _T_2270; // @[Mux.scala 31:69:@45876.4]
  assign _T_2279 = _T_1972 & _T_1518; // @[MemPrimitives.scala 82:228:@45885.4]
  assign _T_2280 = io_wPort_4_en_0 & _T_2279; // @[MemPrimitives.scala 83:102:@45886.4]
  assign _T_2285 = _T_1978 & _T_1524; // @[MemPrimitives.scala 82:228:@45889.4]
  assign _T_2286 = io_wPort_5_en_0 & _T_2285; // @[MemPrimitives.scala 83:102:@45890.4]
  assign _T_2291 = _T_1984 & _T_1530; // @[MemPrimitives.scala 82:228:@45893.4]
  assign _T_2292 = io_wPort_6_en_0 & _T_2291; // @[MemPrimitives.scala 83:102:@45894.4]
  assign _T_2297 = _T_1990 & _T_1536; // @[MemPrimitives.scala 82:228:@45897.4]
  assign _T_2298 = io_wPort_7_en_0 & _T_2297; // @[MemPrimitives.scala 83:102:@45898.4]
  assign _T_2300 = {_T_2280,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45900.4]
  assign _T_2302 = {_T_2286,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45902.4]
  assign _T_2304 = {_T_2292,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45904.4]
  assign _T_2306 = {_T_2298,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45906.4]
  assign _T_2307 = _T_2292 ? _T_2304 : _T_2306; // @[Mux.scala 31:69:@45907.4]
  assign _T_2308 = _T_2286 ? _T_2302 : _T_2307; // @[Mux.scala 31:69:@45908.4]
  assign _T_2309 = _T_2280 ? _T_2300 : _T_2308; // @[Mux.scala 31:69:@45909.4]
  assign _T_2317 = _T_2010 & _T_1556; // @[MemPrimitives.scala 82:228:@45918.4]
  assign _T_2318 = io_wPort_0_en_0 & _T_2317; // @[MemPrimitives.scala 83:102:@45919.4]
  assign _T_2323 = _T_2016 & _T_1562; // @[MemPrimitives.scala 82:228:@45922.4]
  assign _T_2324 = io_wPort_1_en_0 & _T_2323; // @[MemPrimitives.scala 83:102:@45923.4]
  assign _T_2329 = _T_2022 & _T_1568; // @[MemPrimitives.scala 82:228:@45926.4]
  assign _T_2330 = io_wPort_2_en_0 & _T_2329; // @[MemPrimitives.scala 83:102:@45927.4]
  assign _T_2335 = _T_2028 & _T_1574; // @[MemPrimitives.scala 82:228:@45930.4]
  assign _T_2336 = io_wPort_3_en_0 & _T_2335; // @[MemPrimitives.scala 83:102:@45931.4]
  assign _T_2338 = {_T_2318,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45933.4]
  assign _T_2340 = {_T_2324,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@45935.4]
  assign _T_2342 = {_T_2330,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@45937.4]
  assign _T_2344 = {_T_2336,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@45939.4]
  assign _T_2345 = _T_2330 ? _T_2342 : _T_2344; // @[Mux.scala 31:69:@45940.4]
  assign _T_2346 = _T_2324 ? _T_2340 : _T_2345; // @[Mux.scala 31:69:@45941.4]
  assign _T_2347 = _T_2318 ? _T_2338 : _T_2346; // @[Mux.scala 31:69:@45942.4]
  assign _T_2352 = io_wPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45949.4]
  assign _T_2355 = _T_2352 & _T_1214; // @[MemPrimitives.scala 82:228:@45951.4]
  assign _T_2356 = io_wPort_4_en_0 & _T_2355; // @[MemPrimitives.scala 83:102:@45952.4]
  assign _T_2358 = io_wPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45953.4]
  assign _T_2361 = _T_2358 & _T_1220; // @[MemPrimitives.scala 82:228:@45955.4]
  assign _T_2362 = io_wPort_5_en_0 & _T_2361; // @[MemPrimitives.scala 83:102:@45956.4]
  assign _T_2364 = io_wPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45957.4]
  assign _T_2367 = _T_2364 & _T_1226; // @[MemPrimitives.scala 82:228:@45959.4]
  assign _T_2368 = io_wPort_6_en_0 & _T_2367; // @[MemPrimitives.scala 83:102:@45960.4]
  assign _T_2370 = io_wPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45961.4]
  assign _T_2373 = _T_2370 & _T_1232; // @[MemPrimitives.scala 82:228:@45963.4]
  assign _T_2374 = io_wPort_7_en_0 & _T_2373; // @[MemPrimitives.scala 83:102:@45964.4]
  assign _T_2376 = {_T_2356,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@45966.4]
  assign _T_2378 = {_T_2362,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@45968.4]
  assign _T_2380 = {_T_2368,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@45970.4]
  assign _T_2382 = {_T_2374,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@45972.4]
  assign _T_2383 = _T_2368 ? _T_2380 : _T_2382; // @[Mux.scala 31:69:@45973.4]
  assign _T_2384 = _T_2362 ? _T_2378 : _T_2383; // @[Mux.scala 31:69:@45974.4]
  assign _T_2385 = _T_2356 ? _T_2376 : _T_2384; // @[Mux.scala 31:69:@45975.4]
  assign _T_2390 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45982.4]
  assign _T_2393 = _T_2390 & _T_1252; // @[MemPrimitives.scala 82:228:@45984.4]
  assign _T_2394 = io_wPort_0_en_0 & _T_2393; // @[MemPrimitives.scala 83:102:@45985.4]
  assign _T_2396 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45986.4]
  assign _T_2399 = _T_2396 & _T_1258; // @[MemPrimitives.scala 82:228:@45988.4]
  assign _T_2400 = io_wPort_1_en_0 & _T_2399; // @[MemPrimitives.scala 83:102:@45989.4]
  assign _T_2402 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45990.4]
  assign _T_2405 = _T_2402 & _T_1264; // @[MemPrimitives.scala 82:228:@45992.4]
  assign _T_2406 = io_wPort_2_en_0 & _T_2405; // @[MemPrimitives.scala 83:102:@45993.4]
  assign _T_2408 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@45994.4]
  assign _T_2411 = _T_2408 & _T_1270; // @[MemPrimitives.scala 82:228:@45996.4]
  assign _T_2412 = io_wPort_3_en_0 & _T_2411; // @[MemPrimitives.scala 83:102:@45997.4]
  assign _T_2414 = {_T_2394,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@45999.4]
  assign _T_2416 = {_T_2400,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@46001.4]
  assign _T_2418 = {_T_2406,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@46003.4]
  assign _T_2420 = {_T_2412,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@46005.4]
  assign _T_2421 = _T_2406 ? _T_2418 : _T_2420; // @[Mux.scala 31:69:@46006.4]
  assign _T_2422 = _T_2400 ? _T_2416 : _T_2421; // @[Mux.scala 31:69:@46007.4]
  assign _T_2423 = _T_2394 ? _T_2414 : _T_2422; // @[Mux.scala 31:69:@46008.4]
  assign _T_2431 = _T_2352 & _T_1290; // @[MemPrimitives.scala 82:228:@46017.4]
  assign _T_2432 = io_wPort_4_en_0 & _T_2431; // @[MemPrimitives.scala 83:102:@46018.4]
  assign _T_2437 = _T_2358 & _T_1296; // @[MemPrimitives.scala 82:228:@46021.4]
  assign _T_2438 = io_wPort_5_en_0 & _T_2437; // @[MemPrimitives.scala 83:102:@46022.4]
  assign _T_2443 = _T_2364 & _T_1302; // @[MemPrimitives.scala 82:228:@46025.4]
  assign _T_2444 = io_wPort_6_en_0 & _T_2443; // @[MemPrimitives.scala 83:102:@46026.4]
  assign _T_2449 = _T_2370 & _T_1308; // @[MemPrimitives.scala 82:228:@46029.4]
  assign _T_2450 = io_wPort_7_en_0 & _T_2449; // @[MemPrimitives.scala 83:102:@46030.4]
  assign _T_2452 = {_T_2432,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@46032.4]
  assign _T_2454 = {_T_2438,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@46034.4]
  assign _T_2456 = {_T_2444,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@46036.4]
  assign _T_2458 = {_T_2450,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@46038.4]
  assign _T_2459 = _T_2444 ? _T_2456 : _T_2458; // @[Mux.scala 31:69:@46039.4]
  assign _T_2460 = _T_2438 ? _T_2454 : _T_2459; // @[Mux.scala 31:69:@46040.4]
  assign _T_2461 = _T_2432 ? _T_2452 : _T_2460; // @[Mux.scala 31:69:@46041.4]
  assign _T_2469 = _T_2390 & _T_1328; // @[MemPrimitives.scala 82:228:@46050.4]
  assign _T_2470 = io_wPort_0_en_0 & _T_2469; // @[MemPrimitives.scala 83:102:@46051.4]
  assign _T_2475 = _T_2396 & _T_1334; // @[MemPrimitives.scala 82:228:@46054.4]
  assign _T_2476 = io_wPort_1_en_0 & _T_2475; // @[MemPrimitives.scala 83:102:@46055.4]
  assign _T_2481 = _T_2402 & _T_1340; // @[MemPrimitives.scala 82:228:@46058.4]
  assign _T_2482 = io_wPort_2_en_0 & _T_2481; // @[MemPrimitives.scala 83:102:@46059.4]
  assign _T_2487 = _T_2408 & _T_1346; // @[MemPrimitives.scala 82:228:@46062.4]
  assign _T_2488 = io_wPort_3_en_0 & _T_2487; // @[MemPrimitives.scala 83:102:@46063.4]
  assign _T_2490 = {_T_2470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@46065.4]
  assign _T_2492 = {_T_2476,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@46067.4]
  assign _T_2494 = {_T_2482,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@46069.4]
  assign _T_2496 = {_T_2488,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@46071.4]
  assign _T_2497 = _T_2482 ? _T_2494 : _T_2496; // @[Mux.scala 31:69:@46072.4]
  assign _T_2498 = _T_2476 ? _T_2492 : _T_2497; // @[Mux.scala 31:69:@46073.4]
  assign _T_2499 = _T_2470 ? _T_2490 : _T_2498; // @[Mux.scala 31:69:@46074.4]
  assign _T_2507 = _T_2352 & _T_1366; // @[MemPrimitives.scala 82:228:@46083.4]
  assign _T_2508 = io_wPort_4_en_0 & _T_2507; // @[MemPrimitives.scala 83:102:@46084.4]
  assign _T_2513 = _T_2358 & _T_1372; // @[MemPrimitives.scala 82:228:@46087.4]
  assign _T_2514 = io_wPort_5_en_0 & _T_2513; // @[MemPrimitives.scala 83:102:@46088.4]
  assign _T_2519 = _T_2364 & _T_1378; // @[MemPrimitives.scala 82:228:@46091.4]
  assign _T_2520 = io_wPort_6_en_0 & _T_2519; // @[MemPrimitives.scala 83:102:@46092.4]
  assign _T_2525 = _T_2370 & _T_1384; // @[MemPrimitives.scala 82:228:@46095.4]
  assign _T_2526 = io_wPort_7_en_0 & _T_2525; // @[MemPrimitives.scala 83:102:@46096.4]
  assign _T_2528 = {_T_2508,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@46098.4]
  assign _T_2530 = {_T_2514,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@46100.4]
  assign _T_2532 = {_T_2520,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@46102.4]
  assign _T_2534 = {_T_2526,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@46104.4]
  assign _T_2535 = _T_2520 ? _T_2532 : _T_2534; // @[Mux.scala 31:69:@46105.4]
  assign _T_2536 = _T_2514 ? _T_2530 : _T_2535; // @[Mux.scala 31:69:@46106.4]
  assign _T_2537 = _T_2508 ? _T_2528 : _T_2536; // @[Mux.scala 31:69:@46107.4]
  assign _T_2545 = _T_2390 & _T_1404; // @[MemPrimitives.scala 82:228:@46116.4]
  assign _T_2546 = io_wPort_0_en_0 & _T_2545; // @[MemPrimitives.scala 83:102:@46117.4]
  assign _T_2551 = _T_2396 & _T_1410; // @[MemPrimitives.scala 82:228:@46120.4]
  assign _T_2552 = io_wPort_1_en_0 & _T_2551; // @[MemPrimitives.scala 83:102:@46121.4]
  assign _T_2557 = _T_2402 & _T_1416; // @[MemPrimitives.scala 82:228:@46124.4]
  assign _T_2558 = io_wPort_2_en_0 & _T_2557; // @[MemPrimitives.scala 83:102:@46125.4]
  assign _T_2563 = _T_2408 & _T_1422; // @[MemPrimitives.scala 82:228:@46128.4]
  assign _T_2564 = io_wPort_3_en_0 & _T_2563; // @[MemPrimitives.scala 83:102:@46129.4]
  assign _T_2566 = {_T_2546,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@46131.4]
  assign _T_2568 = {_T_2552,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@46133.4]
  assign _T_2570 = {_T_2558,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@46135.4]
  assign _T_2572 = {_T_2564,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@46137.4]
  assign _T_2573 = _T_2558 ? _T_2570 : _T_2572; // @[Mux.scala 31:69:@46138.4]
  assign _T_2574 = _T_2552 ? _T_2568 : _T_2573; // @[Mux.scala 31:69:@46139.4]
  assign _T_2575 = _T_2546 ? _T_2566 : _T_2574; // @[Mux.scala 31:69:@46140.4]
  assign _T_2583 = _T_2352 & _T_1442; // @[MemPrimitives.scala 82:228:@46149.4]
  assign _T_2584 = io_wPort_4_en_0 & _T_2583; // @[MemPrimitives.scala 83:102:@46150.4]
  assign _T_2589 = _T_2358 & _T_1448; // @[MemPrimitives.scala 82:228:@46153.4]
  assign _T_2590 = io_wPort_5_en_0 & _T_2589; // @[MemPrimitives.scala 83:102:@46154.4]
  assign _T_2595 = _T_2364 & _T_1454; // @[MemPrimitives.scala 82:228:@46157.4]
  assign _T_2596 = io_wPort_6_en_0 & _T_2595; // @[MemPrimitives.scala 83:102:@46158.4]
  assign _T_2601 = _T_2370 & _T_1460; // @[MemPrimitives.scala 82:228:@46161.4]
  assign _T_2602 = io_wPort_7_en_0 & _T_2601; // @[MemPrimitives.scala 83:102:@46162.4]
  assign _T_2604 = {_T_2584,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@46164.4]
  assign _T_2606 = {_T_2590,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@46166.4]
  assign _T_2608 = {_T_2596,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@46168.4]
  assign _T_2610 = {_T_2602,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@46170.4]
  assign _T_2611 = _T_2596 ? _T_2608 : _T_2610; // @[Mux.scala 31:69:@46171.4]
  assign _T_2612 = _T_2590 ? _T_2606 : _T_2611; // @[Mux.scala 31:69:@46172.4]
  assign _T_2613 = _T_2584 ? _T_2604 : _T_2612; // @[Mux.scala 31:69:@46173.4]
  assign _T_2621 = _T_2390 & _T_1480; // @[MemPrimitives.scala 82:228:@46182.4]
  assign _T_2622 = io_wPort_0_en_0 & _T_2621; // @[MemPrimitives.scala 83:102:@46183.4]
  assign _T_2627 = _T_2396 & _T_1486; // @[MemPrimitives.scala 82:228:@46186.4]
  assign _T_2628 = io_wPort_1_en_0 & _T_2627; // @[MemPrimitives.scala 83:102:@46187.4]
  assign _T_2633 = _T_2402 & _T_1492; // @[MemPrimitives.scala 82:228:@46190.4]
  assign _T_2634 = io_wPort_2_en_0 & _T_2633; // @[MemPrimitives.scala 83:102:@46191.4]
  assign _T_2639 = _T_2408 & _T_1498; // @[MemPrimitives.scala 82:228:@46194.4]
  assign _T_2640 = io_wPort_3_en_0 & _T_2639; // @[MemPrimitives.scala 83:102:@46195.4]
  assign _T_2642 = {_T_2622,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@46197.4]
  assign _T_2644 = {_T_2628,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@46199.4]
  assign _T_2646 = {_T_2634,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@46201.4]
  assign _T_2648 = {_T_2640,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@46203.4]
  assign _T_2649 = _T_2634 ? _T_2646 : _T_2648; // @[Mux.scala 31:69:@46204.4]
  assign _T_2650 = _T_2628 ? _T_2644 : _T_2649; // @[Mux.scala 31:69:@46205.4]
  assign _T_2651 = _T_2622 ? _T_2642 : _T_2650; // @[Mux.scala 31:69:@46206.4]
  assign _T_2659 = _T_2352 & _T_1518; // @[MemPrimitives.scala 82:228:@46215.4]
  assign _T_2660 = io_wPort_4_en_0 & _T_2659; // @[MemPrimitives.scala 83:102:@46216.4]
  assign _T_2665 = _T_2358 & _T_1524; // @[MemPrimitives.scala 82:228:@46219.4]
  assign _T_2666 = io_wPort_5_en_0 & _T_2665; // @[MemPrimitives.scala 83:102:@46220.4]
  assign _T_2671 = _T_2364 & _T_1530; // @[MemPrimitives.scala 82:228:@46223.4]
  assign _T_2672 = io_wPort_6_en_0 & _T_2671; // @[MemPrimitives.scala 83:102:@46224.4]
  assign _T_2677 = _T_2370 & _T_1536; // @[MemPrimitives.scala 82:228:@46227.4]
  assign _T_2678 = io_wPort_7_en_0 & _T_2677; // @[MemPrimitives.scala 83:102:@46228.4]
  assign _T_2680 = {_T_2660,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@46230.4]
  assign _T_2682 = {_T_2666,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@46232.4]
  assign _T_2684 = {_T_2672,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@46234.4]
  assign _T_2686 = {_T_2678,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@46236.4]
  assign _T_2687 = _T_2672 ? _T_2684 : _T_2686; // @[Mux.scala 31:69:@46237.4]
  assign _T_2688 = _T_2666 ? _T_2682 : _T_2687; // @[Mux.scala 31:69:@46238.4]
  assign _T_2689 = _T_2660 ? _T_2680 : _T_2688; // @[Mux.scala 31:69:@46239.4]
  assign _T_2697 = _T_2390 & _T_1556; // @[MemPrimitives.scala 82:228:@46248.4]
  assign _T_2698 = io_wPort_0_en_0 & _T_2697; // @[MemPrimitives.scala 83:102:@46249.4]
  assign _T_2703 = _T_2396 & _T_1562; // @[MemPrimitives.scala 82:228:@46252.4]
  assign _T_2704 = io_wPort_1_en_0 & _T_2703; // @[MemPrimitives.scala 83:102:@46253.4]
  assign _T_2709 = _T_2402 & _T_1568; // @[MemPrimitives.scala 82:228:@46256.4]
  assign _T_2710 = io_wPort_2_en_0 & _T_2709; // @[MemPrimitives.scala 83:102:@46257.4]
  assign _T_2715 = _T_2408 & _T_1574; // @[MemPrimitives.scala 82:228:@46260.4]
  assign _T_2716 = io_wPort_3_en_0 & _T_2715; // @[MemPrimitives.scala 83:102:@46261.4]
  assign _T_2718 = {_T_2698,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@46263.4]
  assign _T_2720 = {_T_2704,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@46265.4]
  assign _T_2722 = {_T_2710,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@46267.4]
  assign _T_2724 = {_T_2716,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@46269.4]
  assign _T_2725 = _T_2710 ? _T_2722 : _T_2724; // @[Mux.scala 31:69:@46270.4]
  assign _T_2726 = _T_2704 ? _T_2720 : _T_2725; // @[Mux.scala 31:69:@46271.4]
  assign _T_2727 = _T_2698 ? _T_2718 : _T_2726; // @[Mux.scala 31:69:@46272.4]
  assign _T_2732 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46279.4]
  assign _T_2734 = io_rPort_0_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46280.4]
  assign _T_2735 = _T_2732 & _T_2734; // @[MemPrimitives.scala 110:228:@46281.4]
  assign _T_2738 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46283.4]
  assign _T_2740 = io_rPort_1_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46284.4]
  assign _T_2741 = _T_2738 & _T_2740; // @[MemPrimitives.scala 110:228:@46285.4]
  assign _T_2744 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46287.4]
  assign _T_2746 = io_rPort_3_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46288.4]
  assign _T_2747 = _T_2744 & _T_2746; // @[MemPrimitives.scala 110:228:@46289.4]
  assign _T_2750 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46291.4]
  assign _T_2752 = io_rPort_4_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46292.4]
  assign _T_2753 = _T_2750 & _T_2752; // @[MemPrimitives.scala 110:228:@46293.4]
  assign _T_2756 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46295.4]
  assign _T_2758 = io_rPort_5_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46296.4]
  assign _T_2759 = _T_2756 & _T_2758; // @[MemPrimitives.scala 110:228:@46297.4]
  assign _T_2762 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46299.4]
  assign _T_2764 = io_rPort_9_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46300.4]
  assign _T_2765 = _T_2762 & _T_2764; // @[MemPrimitives.scala 110:228:@46301.4]
  assign _T_2768 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46303.4]
  assign _T_2770 = io_rPort_10_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46304.4]
  assign _T_2771 = _T_2768 & _T_2770; // @[MemPrimitives.scala 110:228:@46305.4]
  assign _T_2774 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46307.4]
  assign _T_2776 = io_rPort_13_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46308.4]
  assign _T_2777 = _T_2774 & _T_2776; // @[MemPrimitives.scala 110:228:@46309.4]
  assign _T_2780 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46311.4]
  assign _T_2782 = io_rPort_15_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46312.4]
  assign _T_2783 = _T_2780 & _T_2782; // @[MemPrimitives.scala 110:228:@46313.4]
  assign _T_2786 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46315.4]
  assign _T_2788 = io_rPort_16_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46316.4]
  assign _T_2789 = _T_2786 & _T_2788; // @[MemPrimitives.scala 110:228:@46317.4]
  assign _T_2792 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46319.4]
  assign _T_2794 = io_rPort_17_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46320.4]
  assign _T_2795 = _T_2792 & _T_2794; // @[MemPrimitives.scala 110:228:@46321.4]
  assign _T_2798 = io_rPort_19_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46323.4]
  assign _T_2800 = io_rPort_19_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46324.4]
  assign _T_2801 = _T_2798 & _T_2800; // @[MemPrimitives.scala 110:228:@46325.4]
  assign _T_2804 = io_rPort_22_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46327.4]
  assign _T_2806 = io_rPort_22_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46328.4]
  assign _T_2807 = _T_2804 & _T_2806; // @[MemPrimitives.scala 110:228:@46329.4]
  assign _T_2810 = io_rPort_26_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46331.4]
  assign _T_2812 = io_rPort_26_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46332.4]
  assign _T_2813 = _T_2810 & _T_2812; // @[MemPrimitives.scala 110:228:@46333.4]
  assign _T_2816 = io_rPort_29_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46335.4]
  assign _T_2818 = io_rPort_29_banks_1 == 4'h0; // @[MemPrimitives.scala 110:210:@46336.4]
  assign _T_2819 = _T_2816 & _T_2818; // @[MemPrimitives.scala 110:228:@46337.4]
  assign _T_2821 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@46357.4]
  assign _T_2822 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@46358.4]
  assign _T_2823 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@46359.4]
  assign _T_2824 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@46360.4]
  assign _T_2825 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@46361.4]
  assign _T_2826 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@46362.4]
  assign _T_2827 = StickySelects_io_outs_6; // @[MemPrimitives.scala 123:41:@46363.4]
  assign _T_2828 = StickySelects_io_outs_7; // @[MemPrimitives.scala 123:41:@46364.4]
  assign _T_2829 = StickySelects_io_outs_8; // @[MemPrimitives.scala 123:41:@46365.4]
  assign _T_2830 = StickySelects_io_outs_9; // @[MemPrimitives.scala 123:41:@46366.4]
  assign _T_2831 = StickySelects_io_outs_10; // @[MemPrimitives.scala 123:41:@46367.4]
  assign _T_2832 = StickySelects_io_outs_11; // @[MemPrimitives.scala 123:41:@46368.4]
  assign _T_2833 = StickySelects_io_outs_12; // @[MemPrimitives.scala 123:41:@46369.4]
  assign _T_2834 = StickySelects_io_outs_13; // @[MemPrimitives.scala 123:41:@46370.4]
  assign _T_2835 = StickySelects_io_outs_14; // @[MemPrimitives.scala 123:41:@46371.4]
  assign _T_2837 = {_T_2821,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@46373.4]
  assign _T_2839 = {_T_2822,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@46375.4]
  assign _T_2841 = {_T_2823,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@46377.4]
  assign _T_2843 = {_T_2824,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@46379.4]
  assign _T_2845 = {_T_2825,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@46381.4]
  assign _T_2847 = {_T_2826,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@46383.4]
  assign _T_2849 = {_T_2827,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@46385.4]
  assign _T_2851 = {_T_2828,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@46387.4]
  assign _T_2853 = {_T_2829,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@46389.4]
  assign _T_2855 = {_T_2830,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@46391.4]
  assign _T_2857 = {_T_2831,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@46393.4]
  assign _T_2859 = {_T_2832,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@46395.4]
  assign _T_2861 = {_T_2833,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@46397.4]
  assign _T_2863 = {_T_2834,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@46399.4]
  assign _T_2865 = {_T_2835,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@46401.4]
  assign _T_2866 = _T_2834 ? _T_2863 : _T_2865; // @[Mux.scala 31:69:@46402.4]
  assign _T_2867 = _T_2833 ? _T_2861 : _T_2866; // @[Mux.scala 31:69:@46403.4]
  assign _T_2868 = _T_2832 ? _T_2859 : _T_2867; // @[Mux.scala 31:69:@46404.4]
  assign _T_2869 = _T_2831 ? _T_2857 : _T_2868; // @[Mux.scala 31:69:@46405.4]
  assign _T_2870 = _T_2830 ? _T_2855 : _T_2869; // @[Mux.scala 31:69:@46406.4]
  assign _T_2871 = _T_2829 ? _T_2853 : _T_2870; // @[Mux.scala 31:69:@46407.4]
  assign _T_2872 = _T_2828 ? _T_2851 : _T_2871; // @[Mux.scala 31:69:@46408.4]
  assign _T_2873 = _T_2827 ? _T_2849 : _T_2872; // @[Mux.scala 31:69:@46409.4]
  assign _T_2874 = _T_2826 ? _T_2847 : _T_2873; // @[Mux.scala 31:69:@46410.4]
  assign _T_2875 = _T_2825 ? _T_2845 : _T_2874; // @[Mux.scala 31:69:@46411.4]
  assign _T_2876 = _T_2824 ? _T_2843 : _T_2875; // @[Mux.scala 31:69:@46412.4]
  assign _T_2877 = _T_2823 ? _T_2841 : _T_2876; // @[Mux.scala 31:69:@46413.4]
  assign _T_2878 = _T_2822 ? _T_2839 : _T_2877; // @[Mux.scala 31:69:@46414.4]
  assign _T_2879 = _T_2821 ? _T_2837 : _T_2878; // @[Mux.scala 31:69:@46415.4]
  assign _T_2884 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46422.4]
  assign _T_2886 = io_rPort_2_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46423.4]
  assign _T_2887 = _T_2884 & _T_2886; // @[MemPrimitives.scala 110:228:@46424.4]
  assign _T_2890 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46426.4]
  assign _T_2892 = io_rPort_6_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46427.4]
  assign _T_2893 = _T_2890 & _T_2892; // @[MemPrimitives.scala 110:228:@46428.4]
  assign _T_2896 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46430.4]
  assign _T_2898 = io_rPort_7_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46431.4]
  assign _T_2899 = _T_2896 & _T_2898; // @[MemPrimitives.scala 110:228:@46432.4]
  assign _T_2902 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46434.4]
  assign _T_2904 = io_rPort_8_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46435.4]
  assign _T_2905 = _T_2902 & _T_2904; // @[MemPrimitives.scala 110:228:@46436.4]
  assign _T_2908 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46438.4]
  assign _T_2910 = io_rPort_11_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46439.4]
  assign _T_2911 = _T_2908 & _T_2910; // @[MemPrimitives.scala 110:228:@46440.4]
  assign _T_2914 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46442.4]
  assign _T_2916 = io_rPort_12_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46443.4]
  assign _T_2917 = _T_2914 & _T_2916; // @[MemPrimitives.scala 110:228:@46444.4]
  assign _T_2920 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46446.4]
  assign _T_2922 = io_rPort_14_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46447.4]
  assign _T_2923 = _T_2920 & _T_2922; // @[MemPrimitives.scala 110:228:@46448.4]
  assign _T_2926 = io_rPort_18_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46450.4]
  assign _T_2928 = io_rPort_18_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46451.4]
  assign _T_2929 = _T_2926 & _T_2928; // @[MemPrimitives.scala 110:228:@46452.4]
  assign _T_2932 = io_rPort_20_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46454.4]
  assign _T_2934 = io_rPort_20_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46455.4]
  assign _T_2935 = _T_2932 & _T_2934; // @[MemPrimitives.scala 110:228:@46456.4]
  assign _T_2938 = io_rPort_21_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46458.4]
  assign _T_2940 = io_rPort_21_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46459.4]
  assign _T_2941 = _T_2938 & _T_2940; // @[MemPrimitives.scala 110:228:@46460.4]
  assign _T_2944 = io_rPort_23_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46462.4]
  assign _T_2946 = io_rPort_23_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46463.4]
  assign _T_2947 = _T_2944 & _T_2946; // @[MemPrimitives.scala 110:228:@46464.4]
  assign _T_2950 = io_rPort_24_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46466.4]
  assign _T_2952 = io_rPort_24_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46467.4]
  assign _T_2953 = _T_2950 & _T_2952; // @[MemPrimitives.scala 110:228:@46468.4]
  assign _T_2956 = io_rPort_25_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46470.4]
  assign _T_2958 = io_rPort_25_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46471.4]
  assign _T_2959 = _T_2956 & _T_2958; // @[MemPrimitives.scala 110:228:@46472.4]
  assign _T_2962 = io_rPort_27_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46474.4]
  assign _T_2964 = io_rPort_27_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46475.4]
  assign _T_2965 = _T_2962 & _T_2964; // @[MemPrimitives.scala 110:228:@46476.4]
  assign _T_2968 = io_rPort_28_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@46478.4]
  assign _T_2970 = io_rPort_28_banks_1 == 4'h1; // @[MemPrimitives.scala 110:210:@46479.4]
  assign _T_2971 = _T_2968 & _T_2970; // @[MemPrimitives.scala 110:228:@46480.4]
  assign _T_2973 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@46500.4]
  assign _T_2974 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@46501.4]
  assign _T_2975 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@46502.4]
  assign _T_2976 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@46503.4]
  assign _T_2977 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@46504.4]
  assign _T_2978 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@46505.4]
  assign _T_2979 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 123:41:@46506.4]
  assign _T_2980 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 123:41:@46507.4]
  assign _T_2981 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 123:41:@46508.4]
  assign _T_2982 = StickySelects_1_io_outs_9; // @[MemPrimitives.scala 123:41:@46509.4]
  assign _T_2983 = StickySelects_1_io_outs_10; // @[MemPrimitives.scala 123:41:@46510.4]
  assign _T_2984 = StickySelects_1_io_outs_11; // @[MemPrimitives.scala 123:41:@46511.4]
  assign _T_2985 = StickySelects_1_io_outs_12; // @[MemPrimitives.scala 123:41:@46512.4]
  assign _T_2986 = StickySelects_1_io_outs_13; // @[MemPrimitives.scala 123:41:@46513.4]
  assign _T_2987 = StickySelects_1_io_outs_14; // @[MemPrimitives.scala 123:41:@46514.4]
  assign _T_2989 = {_T_2973,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@46516.4]
  assign _T_2991 = {_T_2974,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@46518.4]
  assign _T_2993 = {_T_2975,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@46520.4]
  assign _T_2995 = {_T_2976,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@46522.4]
  assign _T_2997 = {_T_2977,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@46524.4]
  assign _T_2999 = {_T_2978,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@46526.4]
  assign _T_3001 = {_T_2979,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@46528.4]
  assign _T_3003 = {_T_2980,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@46530.4]
  assign _T_3005 = {_T_2981,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@46532.4]
  assign _T_3007 = {_T_2982,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@46534.4]
  assign _T_3009 = {_T_2983,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@46536.4]
  assign _T_3011 = {_T_2984,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@46538.4]
  assign _T_3013 = {_T_2985,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@46540.4]
  assign _T_3015 = {_T_2986,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@46542.4]
  assign _T_3017 = {_T_2987,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@46544.4]
  assign _T_3018 = _T_2986 ? _T_3015 : _T_3017; // @[Mux.scala 31:69:@46545.4]
  assign _T_3019 = _T_2985 ? _T_3013 : _T_3018; // @[Mux.scala 31:69:@46546.4]
  assign _T_3020 = _T_2984 ? _T_3011 : _T_3019; // @[Mux.scala 31:69:@46547.4]
  assign _T_3021 = _T_2983 ? _T_3009 : _T_3020; // @[Mux.scala 31:69:@46548.4]
  assign _T_3022 = _T_2982 ? _T_3007 : _T_3021; // @[Mux.scala 31:69:@46549.4]
  assign _T_3023 = _T_2981 ? _T_3005 : _T_3022; // @[Mux.scala 31:69:@46550.4]
  assign _T_3024 = _T_2980 ? _T_3003 : _T_3023; // @[Mux.scala 31:69:@46551.4]
  assign _T_3025 = _T_2979 ? _T_3001 : _T_3024; // @[Mux.scala 31:69:@46552.4]
  assign _T_3026 = _T_2978 ? _T_2999 : _T_3025; // @[Mux.scala 31:69:@46553.4]
  assign _T_3027 = _T_2977 ? _T_2997 : _T_3026; // @[Mux.scala 31:69:@46554.4]
  assign _T_3028 = _T_2976 ? _T_2995 : _T_3027; // @[Mux.scala 31:69:@46555.4]
  assign _T_3029 = _T_2975 ? _T_2993 : _T_3028; // @[Mux.scala 31:69:@46556.4]
  assign _T_3030 = _T_2974 ? _T_2991 : _T_3029; // @[Mux.scala 31:69:@46557.4]
  assign _T_3031 = _T_2973 ? _T_2989 : _T_3030; // @[Mux.scala 31:69:@46558.4]
  assign _T_3038 = io_rPort_0_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46566.4]
  assign _T_3039 = _T_2732 & _T_3038; // @[MemPrimitives.scala 110:228:@46567.4]
  assign _T_3044 = io_rPort_1_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46570.4]
  assign _T_3045 = _T_2738 & _T_3044; // @[MemPrimitives.scala 110:228:@46571.4]
  assign _T_3050 = io_rPort_3_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46574.4]
  assign _T_3051 = _T_2744 & _T_3050; // @[MemPrimitives.scala 110:228:@46575.4]
  assign _T_3056 = io_rPort_4_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46578.4]
  assign _T_3057 = _T_2750 & _T_3056; // @[MemPrimitives.scala 110:228:@46579.4]
  assign _T_3062 = io_rPort_5_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46582.4]
  assign _T_3063 = _T_2756 & _T_3062; // @[MemPrimitives.scala 110:228:@46583.4]
  assign _T_3068 = io_rPort_9_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46586.4]
  assign _T_3069 = _T_2762 & _T_3068; // @[MemPrimitives.scala 110:228:@46587.4]
  assign _T_3074 = io_rPort_10_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46590.4]
  assign _T_3075 = _T_2768 & _T_3074; // @[MemPrimitives.scala 110:228:@46591.4]
  assign _T_3080 = io_rPort_13_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46594.4]
  assign _T_3081 = _T_2774 & _T_3080; // @[MemPrimitives.scala 110:228:@46595.4]
  assign _T_3086 = io_rPort_15_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46598.4]
  assign _T_3087 = _T_2780 & _T_3086; // @[MemPrimitives.scala 110:228:@46599.4]
  assign _T_3092 = io_rPort_16_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46602.4]
  assign _T_3093 = _T_2786 & _T_3092; // @[MemPrimitives.scala 110:228:@46603.4]
  assign _T_3098 = io_rPort_17_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46606.4]
  assign _T_3099 = _T_2792 & _T_3098; // @[MemPrimitives.scala 110:228:@46607.4]
  assign _T_3104 = io_rPort_19_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46610.4]
  assign _T_3105 = _T_2798 & _T_3104; // @[MemPrimitives.scala 110:228:@46611.4]
  assign _T_3110 = io_rPort_22_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46614.4]
  assign _T_3111 = _T_2804 & _T_3110; // @[MemPrimitives.scala 110:228:@46615.4]
  assign _T_3116 = io_rPort_26_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46618.4]
  assign _T_3117 = _T_2810 & _T_3116; // @[MemPrimitives.scala 110:228:@46619.4]
  assign _T_3122 = io_rPort_29_banks_1 == 4'h2; // @[MemPrimitives.scala 110:210:@46622.4]
  assign _T_3123 = _T_2816 & _T_3122; // @[MemPrimitives.scala 110:228:@46623.4]
  assign _T_3125 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@46643.4]
  assign _T_3126 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@46644.4]
  assign _T_3127 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@46645.4]
  assign _T_3128 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@46646.4]
  assign _T_3129 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@46647.4]
  assign _T_3130 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@46648.4]
  assign _T_3131 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@46649.4]
  assign _T_3132 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@46650.4]
  assign _T_3133 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 123:41:@46651.4]
  assign _T_3134 = StickySelects_2_io_outs_9; // @[MemPrimitives.scala 123:41:@46652.4]
  assign _T_3135 = StickySelects_2_io_outs_10; // @[MemPrimitives.scala 123:41:@46653.4]
  assign _T_3136 = StickySelects_2_io_outs_11; // @[MemPrimitives.scala 123:41:@46654.4]
  assign _T_3137 = StickySelects_2_io_outs_12; // @[MemPrimitives.scala 123:41:@46655.4]
  assign _T_3138 = StickySelects_2_io_outs_13; // @[MemPrimitives.scala 123:41:@46656.4]
  assign _T_3139 = StickySelects_2_io_outs_14; // @[MemPrimitives.scala 123:41:@46657.4]
  assign _T_3141 = {_T_3125,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@46659.4]
  assign _T_3143 = {_T_3126,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@46661.4]
  assign _T_3145 = {_T_3127,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@46663.4]
  assign _T_3147 = {_T_3128,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@46665.4]
  assign _T_3149 = {_T_3129,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@46667.4]
  assign _T_3151 = {_T_3130,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@46669.4]
  assign _T_3153 = {_T_3131,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@46671.4]
  assign _T_3155 = {_T_3132,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@46673.4]
  assign _T_3157 = {_T_3133,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@46675.4]
  assign _T_3159 = {_T_3134,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@46677.4]
  assign _T_3161 = {_T_3135,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@46679.4]
  assign _T_3163 = {_T_3136,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@46681.4]
  assign _T_3165 = {_T_3137,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@46683.4]
  assign _T_3167 = {_T_3138,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@46685.4]
  assign _T_3169 = {_T_3139,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@46687.4]
  assign _T_3170 = _T_3138 ? _T_3167 : _T_3169; // @[Mux.scala 31:69:@46688.4]
  assign _T_3171 = _T_3137 ? _T_3165 : _T_3170; // @[Mux.scala 31:69:@46689.4]
  assign _T_3172 = _T_3136 ? _T_3163 : _T_3171; // @[Mux.scala 31:69:@46690.4]
  assign _T_3173 = _T_3135 ? _T_3161 : _T_3172; // @[Mux.scala 31:69:@46691.4]
  assign _T_3174 = _T_3134 ? _T_3159 : _T_3173; // @[Mux.scala 31:69:@46692.4]
  assign _T_3175 = _T_3133 ? _T_3157 : _T_3174; // @[Mux.scala 31:69:@46693.4]
  assign _T_3176 = _T_3132 ? _T_3155 : _T_3175; // @[Mux.scala 31:69:@46694.4]
  assign _T_3177 = _T_3131 ? _T_3153 : _T_3176; // @[Mux.scala 31:69:@46695.4]
  assign _T_3178 = _T_3130 ? _T_3151 : _T_3177; // @[Mux.scala 31:69:@46696.4]
  assign _T_3179 = _T_3129 ? _T_3149 : _T_3178; // @[Mux.scala 31:69:@46697.4]
  assign _T_3180 = _T_3128 ? _T_3147 : _T_3179; // @[Mux.scala 31:69:@46698.4]
  assign _T_3181 = _T_3127 ? _T_3145 : _T_3180; // @[Mux.scala 31:69:@46699.4]
  assign _T_3182 = _T_3126 ? _T_3143 : _T_3181; // @[Mux.scala 31:69:@46700.4]
  assign _T_3183 = _T_3125 ? _T_3141 : _T_3182; // @[Mux.scala 31:69:@46701.4]
  assign _T_3190 = io_rPort_2_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46709.4]
  assign _T_3191 = _T_2884 & _T_3190; // @[MemPrimitives.scala 110:228:@46710.4]
  assign _T_3196 = io_rPort_6_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46713.4]
  assign _T_3197 = _T_2890 & _T_3196; // @[MemPrimitives.scala 110:228:@46714.4]
  assign _T_3202 = io_rPort_7_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46717.4]
  assign _T_3203 = _T_2896 & _T_3202; // @[MemPrimitives.scala 110:228:@46718.4]
  assign _T_3208 = io_rPort_8_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46721.4]
  assign _T_3209 = _T_2902 & _T_3208; // @[MemPrimitives.scala 110:228:@46722.4]
  assign _T_3214 = io_rPort_11_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46725.4]
  assign _T_3215 = _T_2908 & _T_3214; // @[MemPrimitives.scala 110:228:@46726.4]
  assign _T_3220 = io_rPort_12_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46729.4]
  assign _T_3221 = _T_2914 & _T_3220; // @[MemPrimitives.scala 110:228:@46730.4]
  assign _T_3226 = io_rPort_14_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46733.4]
  assign _T_3227 = _T_2920 & _T_3226; // @[MemPrimitives.scala 110:228:@46734.4]
  assign _T_3232 = io_rPort_18_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46737.4]
  assign _T_3233 = _T_2926 & _T_3232; // @[MemPrimitives.scala 110:228:@46738.4]
  assign _T_3238 = io_rPort_20_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46741.4]
  assign _T_3239 = _T_2932 & _T_3238; // @[MemPrimitives.scala 110:228:@46742.4]
  assign _T_3244 = io_rPort_21_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46745.4]
  assign _T_3245 = _T_2938 & _T_3244; // @[MemPrimitives.scala 110:228:@46746.4]
  assign _T_3250 = io_rPort_23_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46749.4]
  assign _T_3251 = _T_2944 & _T_3250; // @[MemPrimitives.scala 110:228:@46750.4]
  assign _T_3256 = io_rPort_24_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46753.4]
  assign _T_3257 = _T_2950 & _T_3256; // @[MemPrimitives.scala 110:228:@46754.4]
  assign _T_3262 = io_rPort_25_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46757.4]
  assign _T_3263 = _T_2956 & _T_3262; // @[MemPrimitives.scala 110:228:@46758.4]
  assign _T_3268 = io_rPort_27_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46761.4]
  assign _T_3269 = _T_2962 & _T_3268; // @[MemPrimitives.scala 110:228:@46762.4]
  assign _T_3274 = io_rPort_28_banks_1 == 4'h3; // @[MemPrimitives.scala 110:210:@46765.4]
  assign _T_3275 = _T_2968 & _T_3274; // @[MemPrimitives.scala 110:228:@46766.4]
  assign _T_3277 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@46786.4]
  assign _T_3278 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@46787.4]
  assign _T_3279 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@46788.4]
  assign _T_3280 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@46789.4]
  assign _T_3281 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@46790.4]
  assign _T_3282 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@46791.4]
  assign _T_3283 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@46792.4]
  assign _T_3284 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@46793.4]
  assign _T_3285 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 123:41:@46794.4]
  assign _T_3286 = StickySelects_3_io_outs_9; // @[MemPrimitives.scala 123:41:@46795.4]
  assign _T_3287 = StickySelects_3_io_outs_10; // @[MemPrimitives.scala 123:41:@46796.4]
  assign _T_3288 = StickySelects_3_io_outs_11; // @[MemPrimitives.scala 123:41:@46797.4]
  assign _T_3289 = StickySelects_3_io_outs_12; // @[MemPrimitives.scala 123:41:@46798.4]
  assign _T_3290 = StickySelects_3_io_outs_13; // @[MemPrimitives.scala 123:41:@46799.4]
  assign _T_3291 = StickySelects_3_io_outs_14; // @[MemPrimitives.scala 123:41:@46800.4]
  assign _T_3293 = {_T_3277,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@46802.4]
  assign _T_3295 = {_T_3278,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@46804.4]
  assign _T_3297 = {_T_3279,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@46806.4]
  assign _T_3299 = {_T_3280,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@46808.4]
  assign _T_3301 = {_T_3281,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@46810.4]
  assign _T_3303 = {_T_3282,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@46812.4]
  assign _T_3305 = {_T_3283,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@46814.4]
  assign _T_3307 = {_T_3284,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@46816.4]
  assign _T_3309 = {_T_3285,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@46818.4]
  assign _T_3311 = {_T_3286,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@46820.4]
  assign _T_3313 = {_T_3287,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@46822.4]
  assign _T_3315 = {_T_3288,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@46824.4]
  assign _T_3317 = {_T_3289,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@46826.4]
  assign _T_3319 = {_T_3290,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@46828.4]
  assign _T_3321 = {_T_3291,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@46830.4]
  assign _T_3322 = _T_3290 ? _T_3319 : _T_3321; // @[Mux.scala 31:69:@46831.4]
  assign _T_3323 = _T_3289 ? _T_3317 : _T_3322; // @[Mux.scala 31:69:@46832.4]
  assign _T_3324 = _T_3288 ? _T_3315 : _T_3323; // @[Mux.scala 31:69:@46833.4]
  assign _T_3325 = _T_3287 ? _T_3313 : _T_3324; // @[Mux.scala 31:69:@46834.4]
  assign _T_3326 = _T_3286 ? _T_3311 : _T_3325; // @[Mux.scala 31:69:@46835.4]
  assign _T_3327 = _T_3285 ? _T_3309 : _T_3326; // @[Mux.scala 31:69:@46836.4]
  assign _T_3328 = _T_3284 ? _T_3307 : _T_3327; // @[Mux.scala 31:69:@46837.4]
  assign _T_3329 = _T_3283 ? _T_3305 : _T_3328; // @[Mux.scala 31:69:@46838.4]
  assign _T_3330 = _T_3282 ? _T_3303 : _T_3329; // @[Mux.scala 31:69:@46839.4]
  assign _T_3331 = _T_3281 ? _T_3301 : _T_3330; // @[Mux.scala 31:69:@46840.4]
  assign _T_3332 = _T_3280 ? _T_3299 : _T_3331; // @[Mux.scala 31:69:@46841.4]
  assign _T_3333 = _T_3279 ? _T_3297 : _T_3332; // @[Mux.scala 31:69:@46842.4]
  assign _T_3334 = _T_3278 ? _T_3295 : _T_3333; // @[Mux.scala 31:69:@46843.4]
  assign _T_3335 = _T_3277 ? _T_3293 : _T_3334; // @[Mux.scala 31:69:@46844.4]
  assign _T_3342 = io_rPort_0_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46852.4]
  assign _T_3343 = _T_2732 & _T_3342; // @[MemPrimitives.scala 110:228:@46853.4]
  assign _T_3348 = io_rPort_1_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46856.4]
  assign _T_3349 = _T_2738 & _T_3348; // @[MemPrimitives.scala 110:228:@46857.4]
  assign _T_3354 = io_rPort_3_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46860.4]
  assign _T_3355 = _T_2744 & _T_3354; // @[MemPrimitives.scala 110:228:@46861.4]
  assign _T_3360 = io_rPort_4_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46864.4]
  assign _T_3361 = _T_2750 & _T_3360; // @[MemPrimitives.scala 110:228:@46865.4]
  assign _T_3366 = io_rPort_5_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46868.4]
  assign _T_3367 = _T_2756 & _T_3366; // @[MemPrimitives.scala 110:228:@46869.4]
  assign _T_3372 = io_rPort_9_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46872.4]
  assign _T_3373 = _T_2762 & _T_3372; // @[MemPrimitives.scala 110:228:@46873.4]
  assign _T_3378 = io_rPort_10_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46876.4]
  assign _T_3379 = _T_2768 & _T_3378; // @[MemPrimitives.scala 110:228:@46877.4]
  assign _T_3384 = io_rPort_13_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46880.4]
  assign _T_3385 = _T_2774 & _T_3384; // @[MemPrimitives.scala 110:228:@46881.4]
  assign _T_3390 = io_rPort_15_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46884.4]
  assign _T_3391 = _T_2780 & _T_3390; // @[MemPrimitives.scala 110:228:@46885.4]
  assign _T_3396 = io_rPort_16_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46888.4]
  assign _T_3397 = _T_2786 & _T_3396; // @[MemPrimitives.scala 110:228:@46889.4]
  assign _T_3402 = io_rPort_17_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46892.4]
  assign _T_3403 = _T_2792 & _T_3402; // @[MemPrimitives.scala 110:228:@46893.4]
  assign _T_3408 = io_rPort_19_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46896.4]
  assign _T_3409 = _T_2798 & _T_3408; // @[MemPrimitives.scala 110:228:@46897.4]
  assign _T_3414 = io_rPort_22_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46900.4]
  assign _T_3415 = _T_2804 & _T_3414; // @[MemPrimitives.scala 110:228:@46901.4]
  assign _T_3420 = io_rPort_26_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46904.4]
  assign _T_3421 = _T_2810 & _T_3420; // @[MemPrimitives.scala 110:228:@46905.4]
  assign _T_3426 = io_rPort_29_banks_1 == 4'h4; // @[MemPrimitives.scala 110:210:@46908.4]
  assign _T_3427 = _T_2816 & _T_3426; // @[MemPrimitives.scala 110:228:@46909.4]
  assign _T_3429 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@46929.4]
  assign _T_3430 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@46930.4]
  assign _T_3431 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@46931.4]
  assign _T_3432 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@46932.4]
  assign _T_3433 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@46933.4]
  assign _T_3434 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@46934.4]
  assign _T_3435 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 123:41:@46935.4]
  assign _T_3436 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 123:41:@46936.4]
  assign _T_3437 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 123:41:@46937.4]
  assign _T_3438 = StickySelects_4_io_outs_9; // @[MemPrimitives.scala 123:41:@46938.4]
  assign _T_3439 = StickySelects_4_io_outs_10; // @[MemPrimitives.scala 123:41:@46939.4]
  assign _T_3440 = StickySelects_4_io_outs_11; // @[MemPrimitives.scala 123:41:@46940.4]
  assign _T_3441 = StickySelects_4_io_outs_12; // @[MemPrimitives.scala 123:41:@46941.4]
  assign _T_3442 = StickySelects_4_io_outs_13; // @[MemPrimitives.scala 123:41:@46942.4]
  assign _T_3443 = StickySelects_4_io_outs_14; // @[MemPrimitives.scala 123:41:@46943.4]
  assign _T_3445 = {_T_3429,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@46945.4]
  assign _T_3447 = {_T_3430,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@46947.4]
  assign _T_3449 = {_T_3431,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@46949.4]
  assign _T_3451 = {_T_3432,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@46951.4]
  assign _T_3453 = {_T_3433,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@46953.4]
  assign _T_3455 = {_T_3434,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@46955.4]
  assign _T_3457 = {_T_3435,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@46957.4]
  assign _T_3459 = {_T_3436,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@46959.4]
  assign _T_3461 = {_T_3437,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@46961.4]
  assign _T_3463 = {_T_3438,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@46963.4]
  assign _T_3465 = {_T_3439,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@46965.4]
  assign _T_3467 = {_T_3440,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@46967.4]
  assign _T_3469 = {_T_3441,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@46969.4]
  assign _T_3471 = {_T_3442,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@46971.4]
  assign _T_3473 = {_T_3443,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@46973.4]
  assign _T_3474 = _T_3442 ? _T_3471 : _T_3473; // @[Mux.scala 31:69:@46974.4]
  assign _T_3475 = _T_3441 ? _T_3469 : _T_3474; // @[Mux.scala 31:69:@46975.4]
  assign _T_3476 = _T_3440 ? _T_3467 : _T_3475; // @[Mux.scala 31:69:@46976.4]
  assign _T_3477 = _T_3439 ? _T_3465 : _T_3476; // @[Mux.scala 31:69:@46977.4]
  assign _T_3478 = _T_3438 ? _T_3463 : _T_3477; // @[Mux.scala 31:69:@46978.4]
  assign _T_3479 = _T_3437 ? _T_3461 : _T_3478; // @[Mux.scala 31:69:@46979.4]
  assign _T_3480 = _T_3436 ? _T_3459 : _T_3479; // @[Mux.scala 31:69:@46980.4]
  assign _T_3481 = _T_3435 ? _T_3457 : _T_3480; // @[Mux.scala 31:69:@46981.4]
  assign _T_3482 = _T_3434 ? _T_3455 : _T_3481; // @[Mux.scala 31:69:@46982.4]
  assign _T_3483 = _T_3433 ? _T_3453 : _T_3482; // @[Mux.scala 31:69:@46983.4]
  assign _T_3484 = _T_3432 ? _T_3451 : _T_3483; // @[Mux.scala 31:69:@46984.4]
  assign _T_3485 = _T_3431 ? _T_3449 : _T_3484; // @[Mux.scala 31:69:@46985.4]
  assign _T_3486 = _T_3430 ? _T_3447 : _T_3485; // @[Mux.scala 31:69:@46986.4]
  assign _T_3487 = _T_3429 ? _T_3445 : _T_3486; // @[Mux.scala 31:69:@46987.4]
  assign _T_3494 = io_rPort_2_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@46995.4]
  assign _T_3495 = _T_2884 & _T_3494; // @[MemPrimitives.scala 110:228:@46996.4]
  assign _T_3500 = io_rPort_6_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@46999.4]
  assign _T_3501 = _T_2890 & _T_3500; // @[MemPrimitives.scala 110:228:@47000.4]
  assign _T_3506 = io_rPort_7_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47003.4]
  assign _T_3507 = _T_2896 & _T_3506; // @[MemPrimitives.scala 110:228:@47004.4]
  assign _T_3512 = io_rPort_8_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47007.4]
  assign _T_3513 = _T_2902 & _T_3512; // @[MemPrimitives.scala 110:228:@47008.4]
  assign _T_3518 = io_rPort_11_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47011.4]
  assign _T_3519 = _T_2908 & _T_3518; // @[MemPrimitives.scala 110:228:@47012.4]
  assign _T_3524 = io_rPort_12_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47015.4]
  assign _T_3525 = _T_2914 & _T_3524; // @[MemPrimitives.scala 110:228:@47016.4]
  assign _T_3530 = io_rPort_14_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47019.4]
  assign _T_3531 = _T_2920 & _T_3530; // @[MemPrimitives.scala 110:228:@47020.4]
  assign _T_3536 = io_rPort_18_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47023.4]
  assign _T_3537 = _T_2926 & _T_3536; // @[MemPrimitives.scala 110:228:@47024.4]
  assign _T_3542 = io_rPort_20_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47027.4]
  assign _T_3543 = _T_2932 & _T_3542; // @[MemPrimitives.scala 110:228:@47028.4]
  assign _T_3548 = io_rPort_21_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47031.4]
  assign _T_3549 = _T_2938 & _T_3548; // @[MemPrimitives.scala 110:228:@47032.4]
  assign _T_3554 = io_rPort_23_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47035.4]
  assign _T_3555 = _T_2944 & _T_3554; // @[MemPrimitives.scala 110:228:@47036.4]
  assign _T_3560 = io_rPort_24_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47039.4]
  assign _T_3561 = _T_2950 & _T_3560; // @[MemPrimitives.scala 110:228:@47040.4]
  assign _T_3566 = io_rPort_25_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47043.4]
  assign _T_3567 = _T_2956 & _T_3566; // @[MemPrimitives.scala 110:228:@47044.4]
  assign _T_3572 = io_rPort_27_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47047.4]
  assign _T_3573 = _T_2962 & _T_3572; // @[MemPrimitives.scala 110:228:@47048.4]
  assign _T_3578 = io_rPort_28_banks_1 == 4'h5; // @[MemPrimitives.scala 110:210:@47051.4]
  assign _T_3579 = _T_2968 & _T_3578; // @[MemPrimitives.scala 110:228:@47052.4]
  assign _T_3581 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@47072.4]
  assign _T_3582 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@47073.4]
  assign _T_3583 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@47074.4]
  assign _T_3584 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@47075.4]
  assign _T_3585 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@47076.4]
  assign _T_3586 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@47077.4]
  assign _T_3587 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 123:41:@47078.4]
  assign _T_3588 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 123:41:@47079.4]
  assign _T_3589 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 123:41:@47080.4]
  assign _T_3590 = StickySelects_5_io_outs_9; // @[MemPrimitives.scala 123:41:@47081.4]
  assign _T_3591 = StickySelects_5_io_outs_10; // @[MemPrimitives.scala 123:41:@47082.4]
  assign _T_3592 = StickySelects_5_io_outs_11; // @[MemPrimitives.scala 123:41:@47083.4]
  assign _T_3593 = StickySelects_5_io_outs_12; // @[MemPrimitives.scala 123:41:@47084.4]
  assign _T_3594 = StickySelects_5_io_outs_13; // @[MemPrimitives.scala 123:41:@47085.4]
  assign _T_3595 = StickySelects_5_io_outs_14; // @[MemPrimitives.scala 123:41:@47086.4]
  assign _T_3597 = {_T_3581,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@47088.4]
  assign _T_3599 = {_T_3582,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@47090.4]
  assign _T_3601 = {_T_3583,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@47092.4]
  assign _T_3603 = {_T_3584,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@47094.4]
  assign _T_3605 = {_T_3585,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@47096.4]
  assign _T_3607 = {_T_3586,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@47098.4]
  assign _T_3609 = {_T_3587,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@47100.4]
  assign _T_3611 = {_T_3588,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@47102.4]
  assign _T_3613 = {_T_3589,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@47104.4]
  assign _T_3615 = {_T_3590,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@47106.4]
  assign _T_3617 = {_T_3591,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@47108.4]
  assign _T_3619 = {_T_3592,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@47110.4]
  assign _T_3621 = {_T_3593,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@47112.4]
  assign _T_3623 = {_T_3594,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@47114.4]
  assign _T_3625 = {_T_3595,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@47116.4]
  assign _T_3626 = _T_3594 ? _T_3623 : _T_3625; // @[Mux.scala 31:69:@47117.4]
  assign _T_3627 = _T_3593 ? _T_3621 : _T_3626; // @[Mux.scala 31:69:@47118.4]
  assign _T_3628 = _T_3592 ? _T_3619 : _T_3627; // @[Mux.scala 31:69:@47119.4]
  assign _T_3629 = _T_3591 ? _T_3617 : _T_3628; // @[Mux.scala 31:69:@47120.4]
  assign _T_3630 = _T_3590 ? _T_3615 : _T_3629; // @[Mux.scala 31:69:@47121.4]
  assign _T_3631 = _T_3589 ? _T_3613 : _T_3630; // @[Mux.scala 31:69:@47122.4]
  assign _T_3632 = _T_3588 ? _T_3611 : _T_3631; // @[Mux.scala 31:69:@47123.4]
  assign _T_3633 = _T_3587 ? _T_3609 : _T_3632; // @[Mux.scala 31:69:@47124.4]
  assign _T_3634 = _T_3586 ? _T_3607 : _T_3633; // @[Mux.scala 31:69:@47125.4]
  assign _T_3635 = _T_3585 ? _T_3605 : _T_3634; // @[Mux.scala 31:69:@47126.4]
  assign _T_3636 = _T_3584 ? _T_3603 : _T_3635; // @[Mux.scala 31:69:@47127.4]
  assign _T_3637 = _T_3583 ? _T_3601 : _T_3636; // @[Mux.scala 31:69:@47128.4]
  assign _T_3638 = _T_3582 ? _T_3599 : _T_3637; // @[Mux.scala 31:69:@47129.4]
  assign _T_3639 = _T_3581 ? _T_3597 : _T_3638; // @[Mux.scala 31:69:@47130.4]
  assign _T_3646 = io_rPort_0_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47138.4]
  assign _T_3647 = _T_2732 & _T_3646; // @[MemPrimitives.scala 110:228:@47139.4]
  assign _T_3652 = io_rPort_1_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47142.4]
  assign _T_3653 = _T_2738 & _T_3652; // @[MemPrimitives.scala 110:228:@47143.4]
  assign _T_3658 = io_rPort_3_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47146.4]
  assign _T_3659 = _T_2744 & _T_3658; // @[MemPrimitives.scala 110:228:@47147.4]
  assign _T_3664 = io_rPort_4_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47150.4]
  assign _T_3665 = _T_2750 & _T_3664; // @[MemPrimitives.scala 110:228:@47151.4]
  assign _T_3670 = io_rPort_5_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47154.4]
  assign _T_3671 = _T_2756 & _T_3670; // @[MemPrimitives.scala 110:228:@47155.4]
  assign _T_3676 = io_rPort_9_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47158.4]
  assign _T_3677 = _T_2762 & _T_3676; // @[MemPrimitives.scala 110:228:@47159.4]
  assign _T_3682 = io_rPort_10_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47162.4]
  assign _T_3683 = _T_2768 & _T_3682; // @[MemPrimitives.scala 110:228:@47163.4]
  assign _T_3688 = io_rPort_13_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47166.4]
  assign _T_3689 = _T_2774 & _T_3688; // @[MemPrimitives.scala 110:228:@47167.4]
  assign _T_3694 = io_rPort_15_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47170.4]
  assign _T_3695 = _T_2780 & _T_3694; // @[MemPrimitives.scala 110:228:@47171.4]
  assign _T_3700 = io_rPort_16_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47174.4]
  assign _T_3701 = _T_2786 & _T_3700; // @[MemPrimitives.scala 110:228:@47175.4]
  assign _T_3706 = io_rPort_17_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47178.4]
  assign _T_3707 = _T_2792 & _T_3706; // @[MemPrimitives.scala 110:228:@47179.4]
  assign _T_3712 = io_rPort_19_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47182.4]
  assign _T_3713 = _T_2798 & _T_3712; // @[MemPrimitives.scala 110:228:@47183.4]
  assign _T_3718 = io_rPort_22_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47186.4]
  assign _T_3719 = _T_2804 & _T_3718; // @[MemPrimitives.scala 110:228:@47187.4]
  assign _T_3724 = io_rPort_26_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47190.4]
  assign _T_3725 = _T_2810 & _T_3724; // @[MemPrimitives.scala 110:228:@47191.4]
  assign _T_3730 = io_rPort_29_banks_1 == 4'h6; // @[MemPrimitives.scala 110:210:@47194.4]
  assign _T_3731 = _T_2816 & _T_3730; // @[MemPrimitives.scala 110:228:@47195.4]
  assign _T_3733 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@47215.4]
  assign _T_3734 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@47216.4]
  assign _T_3735 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@47217.4]
  assign _T_3736 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@47218.4]
  assign _T_3737 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@47219.4]
  assign _T_3738 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@47220.4]
  assign _T_3739 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@47221.4]
  assign _T_3740 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@47222.4]
  assign _T_3741 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 123:41:@47223.4]
  assign _T_3742 = StickySelects_6_io_outs_9; // @[MemPrimitives.scala 123:41:@47224.4]
  assign _T_3743 = StickySelects_6_io_outs_10; // @[MemPrimitives.scala 123:41:@47225.4]
  assign _T_3744 = StickySelects_6_io_outs_11; // @[MemPrimitives.scala 123:41:@47226.4]
  assign _T_3745 = StickySelects_6_io_outs_12; // @[MemPrimitives.scala 123:41:@47227.4]
  assign _T_3746 = StickySelects_6_io_outs_13; // @[MemPrimitives.scala 123:41:@47228.4]
  assign _T_3747 = StickySelects_6_io_outs_14; // @[MemPrimitives.scala 123:41:@47229.4]
  assign _T_3749 = {_T_3733,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@47231.4]
  assign _T_3751 = {_T_3734,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@47233.4]
  assign _T_3753 = {_T_3735,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@47235.4]
  assign _T_3755 = {_T_3736,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@47237.4]
  assign _T_3757 = {_T_3737,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@47239.4]
  assign _T_3759 = {_T_3738,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@47241.4]
  assign _T_3761 = {_T_3739,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@47243.4]
  assign _T_3763 = {_T_3740,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@47245.4]
  assign _T_3765 = {_T_3741,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@47247.4]
  assign _T_3767 = {_T_3742,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@47249.4]
  assign _T_3769 = {_T_3743,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@47251.4]
  assign _T_3771 = {_T_3744,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@47253.4]
  assign _T_3773 = {_T_3745,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@47255.4]
  assign _T_3775 = {_T_3746,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@47257.4]
  assign _T_3777 = {_T_3747,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@47259.4]
  assign _T_3778 = _T_3746 ? _T_3775 : _T_3777; // @[Mux.scala 31:69:@47260.4]
  assign _T_3779 = _T_3745 ? _T_3773 : _T_3778; // @[Mux.scala 31:69:@47261.4]
  assign _T_3780 = _T_3744 ? _T_3771 : _T_3779; // @[Mux.scala 31:69:@47262.4]
  assign _T_3781 = _T_3743 ? _T_3769 : _T_3780; // @[Mux.scala 31:69:@47263.4]
  assign _T_3782 = _T_3742 ? _T_3767 : _T_3781; // @[Mux.scala 31:69:@47264.4]
  assign _T_3783 = _T_3741 ? _T_3765 : _T_3782; // @[Mux.scala 31:69:@47265.4]
  assign _T_3784 = _T_3740 ? _T_3763 : _T_3783; // @[Mux.scala 31:69:@47266.4]
  assign _T_3785 = _T_3739 ? _T_3761 : _T_3784; // @[Mux.scala 31:69:@47267.4]
  assign _T_3786 = _T_3738 ? _T_3759 : _T_3785; // @[Mux.scala 31:69:@47268.4]
  assign _T_3787 = _T_3737 ? _T_3757 : _T_3786; // @[Mux.scala 31:69:@47269.4]
  assign _T_3788 = _T_3736 ? _T_3755 : _T_3787; // @[Mux.scala 31:69:@47270.4]
  assign _T_3789 = _T_3735 ? _T_3753 : _T_3788; // @[Mux.scala 31:69:@47271.4]
  assign _T_3790 = _T_3734 ? _T_3751 : _T_3789; // @[Mux.scala 31:69:@47272.4]
  assign _T_3791 = _T_3733 ? _T_3749 : _T_3790; // @[Mux.scala 31:69:@47273.4]
  assign _T_3798 = io_rPort_2_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47281.4]
  assign _T_3799 = _T_2884 & _T_3798; // @[MemPrimitives.scala 110:228:@47282.4]
  assign _T_3804 = io_rPort_6_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47285.4]
  assign _T_3805 = _T_2890 & _T_3804; // @[MemPrimitives.scala 110:228:@47286.4]
  assign _T_3810 = io_rPort_7_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47289.4]
  assign _T_3811 = _T_2896 & _T_3810; // @[MemPrimitives.scala 110:228:@47290.4]
  assign _T_3816 = io_rPort_8_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47293.4]
  assign _T_3817 = _T_2902 & _T_3816; // @[MemPrimitives.scala 110:228:@47294.4]
  assign _T_3822 = io_rPort_11_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47297.4]
  assign _T_3823 = _T_2908 & _T_3822; // @[MemPrimitives.scala 110:228:@47298.4]
  assign _T_3828 = io_rPort_12_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47301.4]
  assign _T_3829 = _T_2914 & _T_3828; // @[MemPrimitives.scala 110:228:@47302.4]
  assign _T_3834 = io_rPort_14_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47305.4]
  assign _T_3835 = _T_2920 & _T_3834; // @[MemPrimitives.scala 110:228:@47306.4]
  assign _T_3840 = io_rPort_18_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47309.4]
  assign _T_3841 = _T_2926 & _T_3840; // @[MemPrimitives.scala 110:228:@47310.4]
  assign _T_3846 = io_rPort_20_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47313.4]
  assign _T_3847 = _T_2932 & _T_3846; // @[MemPrimitives.scala 110:228:@47314.4]
  assign _T_3852 = io_rPort_21_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47317.4]
  assign _T_3853 = _T_2938 & _T_3852; // @[MemPrimitives.scala 110:228:@47318.4]
  assign _T_3858 = io_rPort_23_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47321.4]
  assign _T_3859 = _T_2944 & _T_3858; // @[MemPrimitives.scala 110:228:@47322.4]
  assign _T_3864 = io_rPort_24_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47325.4]
  assign _T_3865 = _T_2950 & _T_3864; // @[MemPrimitives.scala 110:228:@47326.4]
  assign _T_3870 = io_rPort_25_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47329.4]
  assign _T_3871 = _T_2956 & _T_3870; // @[MemPrimitives.scala 110:228:@47330.4]
  assign _T_3876 = io_rPort_27_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47333.4]
  assign _T_3877 = _T_2962 & _T_3876; // @[MemPrimitives.scala 110:228:@47334.4]
  assign _T_3882 = io_rPort_28_banks_1 == 4'h7; // @[MemPrimitives.scala 110:210:@47337.4]
  assign _T_3883 = _T_2968 & _T_3882; // @[MemPrimitives.scala 110:228:@47338.4]
  assign _T_3885 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@47358.4]
  assign _T_3886 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@47359.4]
  assign _T_3887 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@47360.4]
  assign _T_3888 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@47361.4]
  assign _T_3889 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@47362.4]
  assign _T_3890 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@47363.4]
  assign _T_3891 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@47364.4]
  assign _T_3892 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@47365.4]
  assign _T_3893 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 123:41:@47366.4]
  assign _T_3894 = StickySelects_7_io_outs_9; // @[MemPrimitives.scala 123:41:@47367.4]
  assign _T_3895 = StickySelects_7_io_outs_10; // @[MemPrimitives.scala 123:41:@47368.4]
  assign _T_3896 = StickySelects_7_io_outs_11; // @[MemPrimitives.scala 123:41:@47369.4]
  assign _T_3897 = StickySelects_7_io_outs_12; // @[MemPrimitives.scala 123:41:@47370.4]
  assign _T_3898 = StickySelects_7_io_outs_13; // @[MemPrimitives.scala 123:41:@47371.4]
  assign _T_3899 = StickySelects_7_io_outs_14; // @[MemPrimitives.scala 123:41:@47372.4]
  assign _T_3901 = {_T_3885,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@47374.4]
  assign _T_3903 = {_T_3886,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@47376.4]
  assign _T_3905 = {_T_3887,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@47378.4]
  assign _T_3907 = {_T_3888,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@47380.4]
  assign _T_3909 = {_T_3889,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@47382.4]
  assign _T_3911 = {_T_3890,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@47384.4]
  assign _T_3913 = {_T_3891,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@47386.4]
  assign _T_3915 = {_T_3892,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@47388.4]
  assign _T_3917 = {_T_3893,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@47390.4]
  assign _T_3919 = {_T_3894,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@47392.4]
  assign _T_3921 = {_T_3895,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@47394.4]
  assign _T_3923 = {_T_3896,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@47396.4]
  assign _T_3925 = {_T_3897,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@47398.4]
  assign _T_3927 = {_T_3898,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@47400.4]
  assign _T_3929 = {_T_3899,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@47402.4]
  assign _T_3930 = _T_3898 ? _T_3927 : _T_3929; // @[Mux.scala 31:69:@47403.4]
  assign _T_3931 = _T_3897 ? _T_3925 : _T_3930; // @[Mux.scala 31:69:@47404.4]
  assign _T_3932 = _T_3896 ? _T_3923 : _T_3931; // @[Mux.scala 31:69:@47405.4]
  assign _T_3933 = _T_3895 ? _T_3921 : _T_3932; // @[Mux.scala 31:69:@47406.4]
  assign _T_3934 = _T_3894 ? _T_3919 : _T_3933; // @[Mux.scala 31:69:@47407.4]
  assign _T_3935 = _T_3893 ? _T_3917 : _T_3934; // @[Mux.scala 31:69:@47408.4]
  assign _T_3936 = _T_3892 ? _T_3915 : _T_3935; // @[Mux.scala 31:69:@47409.4]
  assign _T_3937 = _T_3891 ? _T_3913 : _T_3936; // @[Mux.scala 31:69:@47410.4]
  assign _T_3938 = _T_3890 ? _T_3911 : _T_3937; // @[Mux.scala 31:69:@47411.4]
  assign _T_3939 = _T_3889 ? _T_3909 : _T_3938; // @[Mux.scala 31:69:@47412.4]
  assign _T_3940 = _T_3888 ? _T_3907 : _T_3939; // @[Mux.scala 31:69:@47413.4]
  assign _T_3941 = _T_3887 ? _T_3905 : _T_3940; // @[Mux.scala 31:69:@47414.4]
  assign _T_3942 = _T_3886 ? _T_3903 : _T_3941; // @[Mux.scala 31:69:@47415.4]
  assign _T_3943 = _T_3885 ? _T_3901 : _T_3942; // @[Mux.scala 31:69:@47416.4]
  assign _T_3950 = io_rPort_0_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47424.4]
  assign _T_3951 = _T_2732 & _T_3950; // @[MemPrimitives.scala 110:228:@47425.4]
  assign _T_3956 = io_rPort_1_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47428.4]
  assign _T_3957 = _T_2738 & _T_3956; // @[MemPrimitives.scala 110:228:@47429.4]
  assign _T_3962 = io_rPort_3_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47432.4]
  assign _T_3963 = _T_2744 & _T_3962; // @[MemPrimitives.scala 110:228:@47433.4]
  assign _T_3968 = io_rPort_4_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47436.4]
  assign _T_3969 = _T_2750 & _T_3968; // @[MemPrimitives.scala 110:228:@47437.4]
  assign _T_3974 = io_rPort_5_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47440.4]
  assign _T_3975 = _T_2756 & _T_3974; // @[MemPrimitives.scala 110:228:@47441.4]
  assign _T_3980 = io_rPort_9_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47444.4]
  assign _T_3981 = _T_2762 & _T_3980; // @[MemPrimitives.scala 110:228:@47445.4]
  assign _T_3986 = io_rPort_10_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47448.4]
  assign _T_3987 = _T_2768 & _T_3986; // @[MemPrimitives.scala 110:228:@47449.4]
  assign _T_3992 = io_rPort_13_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47452.4]
  assign _T_3993 = _T_2774 & _T_3992; // @[MemPrimitives.scala 110:228:@47453.4]
  assign _T_3998 = io_rPort_15_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47456.4]
  assign _T_3999 = _T_2780 & _T_3998; // @[MemPrimitives.scala 110:228:@47457.4]
  assign _T_4004 = io_rPort_16_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47460.4]
  assign _T_4005 = _T_2786 & _T_4004; // @[MemPrimitives.scala 110:228:@47461.4]
  assign _T_4010 = io_rPort_17_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47464.4]
  assign _T_4011 = _T_2792 & _T_4010; // @[MemPrimitives.scala 110:228:@47465.4]
  assign _T_4016 = io_rPort_19_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47468.4]
  assign _T_4017 = _T_2798 & _T_4016; // @[MemPrimitives.scala 110:228:@47469.4]
  assign _T_4022 = io_rPort_22_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47472.4]
  assign _T_4023 = _T_2804 & _T_4022; // @[MemPrimitives.scala 110:228:@47473.4]
  assign _T_4028 = io_rPort_26_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47476.4]
  assign _T_4029 = _T_2810 & _T_4028; // @[MemPrimitives.scala 110:228:@47477.4]
  assign _T_4034 = io_rPort_29_banks_1 == 4'h8; // @[MemPrimitives.scala 110:210:@47480.4]
  assign _T_4035 = _T_2816 & _T_4034; // @[MemPrimitives.scala 110:228:@47481.4]
  assign _T_4037 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@47501.4]
  assign _T_4038 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@47502.4]
  assign _T_4039 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@47503.4]
  assign _T_4040 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@47504.4]
  assign _T_4041 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@47505.4]
  assign _T_4042 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@47506.4]
  assign _T_4043 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 123:41:@47507.4]
  assign _T_4044 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 123:41:@47508.4]
  assign _T_4045 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 123:41:@47509.4]
  assign _T_4046 = StickySelects_8_io_outs_9; // @[MemPrimitives.scala 123:41:@47510.4]
  assign _T_4047 = StickySelects_8_io_outs_10; // @[MemPrimitives.scala 123:41:@47511.4]
  assign _T_4048 = StickySelects_8_io_outs_11; // @[MemPrimitives.scala 123:41:@47512.4]
  assign _T_4049 = StickySelects_8_io_outs_12; // @[MemPrimitives.scala 123:41:@47513.4]
  assign _T_4050 = StickySelects_8_io_outs_13; // @[MemPrimitives.scala 123:41:@47514.4]
  assign _T_4051 = StickySelects_8_io_outs_14; // @[MemPrimitives.scala 123:41:@47515.4]
  assign _T_4053 = {_T_4037,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@47517.4]
  assign _T_4055 = {_T_4038,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@47519.4]
  assign _T_4057 = {_T_4039,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@47521.4]
  assign _T_4059 = {_T_4040,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@47523.4]
  assign _T_4061 = {_T_4041,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@47525.4]
  assign _T_4063 = {_T_4042,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@47527.4]
  assign _T_4065 = {_T_4043,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@47529.4]
  assign _T_4067 = {_T_4044,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@47531.4]
  assign _T_4069 = {_T_4045,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@47533.4]
  assign _T_4071 = {_T_4046,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@47535.4]
  assign _T_4073 = {_T_4047,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@47537.4]
  assign _T_4075 = {_T_4048,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@47539.4]
  assign _T_4077 = {_T_4049,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@47541.4]
  assign _T_4079 = {_T_4050,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@47543.4]
  assign _T_4081 = {_T_4051,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@47545.4]
  assign _T_4082 = _T_4050 ? _T_4079 : _T_4081; // @[Mux.scala 31:69:@47546.4]
  assign _T_4083 = _T_4049 ? _T_4077 : _T_4082; // @[Mux.scala 31:69:@47547.4]
  assign _T_4084 = _T_4048 ? _T_4075 : _T_4083; // @[Mux.scala 31:69:@47548.4]
  assign _T_4085 = _T_4047 ? _T_4073 : _T_4084; // @[Mux.scala 31:69:@47549.4]
  assign _T_4086 = _T_4046 ? _T_4071 : _T_4085; // @[Mux.scala 31:69:@47550.4]
  assign _T_4087 = _T_4045 ? _T_4069 : _T_4086; // @[Mux.scala 31:69:@47551.4]
  assign _T_4088 = _T_4044 ? _T_4067 : _T_4087; // @[Mux.scala 31:69:@47552.4]
  assign _T_4089 = _T_4043 ? _T_4065 : _T_4088; // @[Mux.scala 31:69:@47553.4]
  assign _T_4090 = _T_4042 ? _T_4063 : _T_4089; // @[Mux.scala 31:69:@47554.4]
  assign _T_4091 = _T_4041 ? _T_4061 : _T_4090; // @[Mux.scala 31:69:@47555.4]
  assign _T_4092 = _T_4040 ? _T_4059 : _T_4091; // @[Mux.scala 31:69:@47556.4]
  assign _T_4093 = _T_4039 ? _T_4057 : _T_4092; // @[Mux.scala 31:69:@47557.4]
  assign _T_4094 = _T_4038 ? _T_4055 : _T_4093; // @[Mux.scala 31:69:@47558.4]
  assign _T_4095 = _T_4037 ? _T_4053 : _T_4094; // @[Mux.scala 31:69:@47559.4]
  assign _T_4102 = io_rPort_2_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47567.4]
  assign _T_4103 = _T_2884 & _T_4102; // @[MemPrimitives.scala 110:228:@47568.4]
  assign _T_4108 = io_rPort_6_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47571.4]
  assign _T_4109 = _T_2890 & _T_4108; // @[MemPrimitives.scala 110:228:@47572.4]
  assign _T_4114 = io_rPort_7_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47575.4]
  assign _T_4115 = _T_2896 & _T_4114; // @[MemPrimitives.scala 110:228:@47576.4]
  assign _T_4120 = io_rPort_8_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47579.4]
  assign _T_4121 = _T_2902 & _T_4120; // @[MemPrimitives.scala 110:228:@47580.4]
  assign _T_4126 = io_rPort_11_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47583.4]
  assign _T_4127 = _T_2908 & _T_4126; // @[MemPrimitives.scala 110:228:@47584.4]
  assign _T_4132 = io_rPort_12_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47587.4]
  assign _T_4133 = _T_2914 & _T_4132; // @[MemPrimitives.scala 110:228:@47588.4]
  assign _T_4138 = io_rPort_14_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47591.4]
  assign _T_4139 = _T_2920 & _T_4138; // @[MemPrimitives.scala 110:228:@47592.4]
  assign _T_4144 = io_rPort_18_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47595.4]
  assign _T_4145 = _T_2926 & _T_4144; // @[MemPrimitives.scala 110:228:@47596.4]
  assign _T_4150 = io_rPort_20_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47599.4]
  assign _T_4151 = _T_2932 & _T_4150; // @[MemPrimitives.scala 110:228:@47600.4]
  assign _T_4156 = io_rPort_21_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47603.4]
  assign _T_4157 = _T_2938 & _T_4156; // @[MemPrimitives.scala 110:228:@47604.4]
  assign _T_4162 = io_rPort_23_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47607.4]
  assign _T_4163 = _T_2944 & _T_4162; // @[MemPrimitives.scala 110:228:@47608.4]
  assign _T_4168 = io_rPort_24_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47611.4]
  assign _T_4169 = _T_2950 & _T_4168; // @[MemPrimitives.scala 110:228:@47612.4]
  assign _T_4174 = io_rPort_25_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47615.4]
  assign _T_4175 = _T_2956 & _T_4174; // @[MemPrimitives.scala 110:228:@47616.4]
  assign _T_4180 = io_rPort_27_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47619.4]
  assign _T_4181 = _T_2962 & _T_4180; // @[MemPrimitives.scala 110:228:@47620.4]
  assign _T_4186 = io_rPort_28_banks_1 == 4'h9; // @[MemPrimitives.scala 110:210:@47623.4]
  assign _T_4187 = _T_2968 & _T_4186; // @[MemPrimitives.scala 110:228:@47624.4]
  assign _T_4189 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@47644.4]
  assign _T_4190 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@47645.4]
  assign _T_4191 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@47646.4]
  assign _T_4192 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@47647.4]
  assign _T_4193 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@47648.4]
  assign _T_4194 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@47649.4]
  assign _T_4195 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 123:41:@47650.4]
  assign _T_4196 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 123:41:@47651.4]
  assign _T_4197 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 123:41:@47652.4]
  assign _T_4198 = StickySelects_9_io_outs_9; // @[MemPrimitives.scala 123:41:@47653.4]
  assign _T_4199 = StickySelects_9_io_outs_10; // @[MemPrimitives.scala 123:41:@47654.4]
  assign _T_4200 = StickySelects_9_io_outs_11; // @[MemPrimitives.scala 123:41:@47655.4]
  assign _T_4201 = StickySelects_9_io_outs_12; // @[MemPrimitives.scala 123:41:@47656.4]
  assign _T_4202 = StickySelects_9_io_outs_13; // @[MemPrimitives.scala 123:41:@47657.4]
  assign _T_4203 = StickySelects_9_io_outs_14; // @[MemPrimitives.scala 123:41:@47658.4]
  assign _T_4205 = {_T_4189,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@47660.4]
  assign _T_4207 = {_T_4190,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@47662.4]
  assign _T_4209 = {_T_4191,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@47664.4]
  assign _T_4211 = {_T_4192,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@47666.4]
  assign _T_4213 = {_T_4193,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@47668.4]
  assign _T_4215 = {_T_4194,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@47670.4]
  assign _T_4217 = {_T_4195,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@47672.4]
  assign _T_4219 = {_T_4196,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@47674.4]
  assign _T_4221 = {_T_4197,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@47676.4]
  assign _T_4223 = {_T_4198,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@47678.4]
  assign _T_4225 = {_T_4199,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@47680.4]
  assign _T_4227 = {_T_4200,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@47682.4]
  assign _T_4229 = {_T_4201,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@47684.4]
  assign _T_4231 = {_T_4202,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@47686.4]
  assign _T_4233 = {_T_4203,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@47688.4]
  assign _T_4234 = _T_4202 ? _T_4231 : _T_4233; // @[Mux.scala 31:69:@47689.4]
  assign _T_4235 = _T_4201 ? _T_4229 : _T_4234; // @[Mux.scala 31:69:@47690.4]
  assign _T_4236 = _T_4200 ? _T_4227 : _T_4235; // @[Mux.scala 31:69:@47691.4]
  assign _T_4237 = _T_4199 ? _T_4225 : _T_4236; // @[Mux.scala 31:69:@47692.4]
  assign _T_4238 = _T_4198 ? _T_4223 : _T_4237; // @[Mux.scala 31:69:@47693.4]
  assign _T_4239 = _T_4197 ? _T_4221 : _T_4238; // @[Mux.scala 31:69:@47694.4]
  assign _T_4240 = _T_4196 ? _T_4219 : _T_4239; // @[Mux.scala 31:69:@47695.4]
  assign _T_4241 = _T_4195 ? _T_4217 : _T_4240; // @[Mux.scala 31:69:@47696.4]
  assign _T_4242 = _T_4194 ? _T_4215 : _T_4241; // @[Mux.scala 31:69:@47697.4]
  assign _T_4243 = _T_4193 ? _T_4213 : _T_4242; // @[Mux.scala 31:69:@47698.4]
  assign _T_4244 = _T_4192 ? _T_4211 : _T_4243; // @[Mux.scala 31:69:@47699.4]
  assign _T_4245 = _T_4191 ? _T_4209 : _T_4244; // @[Mux.scala 31:69:@47700.4]
  assign _T_4246 = _T_4190 ? _T_4207 : _T_4245; // @[Mux.scala 31:69:@47701.4]
  assign _T_4247 = _T_4189 ? _T_4205 : _T_4246; // @[Mux.scala 31:69:@47702.4]
  assign _T_4252 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47709.4]
  assign _T_4255 = _T_4252 & _T_2734; // @[MemPrimitives.scala 110:228:@47711.4]
  assign _T_4258 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47713.4]
  assign _T_4261 = _T_4258 & _T_2740; // @[MemPrimitives.scala 110:228:@47715.4]
  assign _T_4264 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47717.4]
  assign _T_4267 = _T_4264 & _T_2746; // @[MemPrimitives.scala 110:228:@47719.4]
  assign _T_4270 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47721.4]
  assign _T_4273 = _T_4270 & _T_2752; // @[MemPrimitives.scala 110:228:@47723.4]
  assign _T_4276 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47725.4]
  assign _T_4279 = _T_4276 & _T_2758; // @[MemPrimitives.scala 110:228:@47727.4]
  assign _T_4282 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47729.4]
  assign _T_4285 = _T_4282 & _T_2764; // @[MemPrimitives.scala 110:228:@47731.4]
  assign _T_4288 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47733.4]
  assign _T_4291 = _T_4288 & _T_2770; // @[MemPrimitives.scala 110:228:@47735.4]
  assign _T_4294 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47737.4]
  assign _T_4297 = _T_4294 & _T_2776; // @[MemPrimitives.scala 110:228:@47739.4]
  assign _T_4300 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47741.4]
  assign _T_4303 = _T_4300 & _T_2782; // @[MemPrimitives.scala 110:228:@47743.4]
  assign _T_4306 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47745.4]
  assign _T_4309 = _T_4306 & _T_2788; // @[MemPrimitives.scala 110:228:@47747.4]
  assign _T_4312 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47749.4]
  assign _T_4315 = _T_4312 & _T_2794; // @[MemPrimitives.scala 110:228:@47751.4]
  assign _T_4318 = io_rPort_19_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47753.4]
  assign _T_4321 = _T_4318 & _T_2800; // @[MemPrimitives.scala 110:228:@47755.4]
  assign _T_4324 = io_rPort_22_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47757.4]
  assign _T_4327 = _T_4324 & _T_2806; // @[MemPrimitives.scala 110:228:@47759.4]
  assign _T_4330 = io_rPort_26_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47761.4]
  assign _T_4333 = _T_4330 & _T_2812; // @[MemPrimitives.scala 110:228:@47763.4]
  assign _T_4336 = io_rPort_29_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47765.4]
  assign _T_4339 = _T_4336 & _T_2818; // @[MemPrimitives.scala 110:228:@47767.4]
  assign _T_4341 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@47787.4]
  assign _T_4342 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@47788.4]
  assign _T_4343 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@47789.4]
  assign _T_4344 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@47790.4]
  assign _T_4345 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@47791.4]
  assign _T_4346 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@47792.4]
  assign _T_4347 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@47793.4]
  assign _T_4348 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@47794.4]
  assign _T_4349 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 123:41:@47795.4]
  assign _T_4350 = StickySelects_10_io_outs_9; // @[MemPrimitives.scala 123:41:@47796.4]
  assign _T_4351 = StickySelects_10_io_outs_10; // @[MemPrimitives.scala 123:41:@47797.4]
  assign _T_4352 = StickySelects_10_io_outs_11; // @[MemPrimitives.scala 123:41:@47798.4]
  assign _T_4353 = StickySelects_10_io_outs_12; // @[MemPrimitives.scala 123:41:@47799.4]
  assign _T_4354 = StickySelects_10_io_outs_13; // @[MemPrimitives.scala 123:41:@47800.4]
  assign _T_4355 = StickySelects_10_io_outs_14; // @[MemPrimitives.scala 123:41:@47801.4]
  assign _T_4357 = {_T_4341,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@47803.4]
  assign _T_4359 = {_T_4342,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@47805.4]
  assign _T_4361 = {_T_4343,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@47807.4]
  assign _T_4363 = {_T_4344,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@47809.4]
  assign _T_4365 = {_T_4345,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@47811.4]
  assign _T_4367 = {_T_4346,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@47813.4]
  assign _T_4369 = {_T_4347,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@47815.4]
  assign _T_4371 = {_T_4348,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@47817.4]
  assign _T_4373 = {_T_4349,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@47819.4]
  assign _T_4375 = {_T_4350,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@47821.4]
  assign _T_4377 = {_T_4351,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@47823.4]
  assign _T_4379 = {_T_4352,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@47825.4]
  assign _T_4381 = {_T_4353,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@47827.4]
  assign _T_4383 = {_T_4354,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@47829.4]
  assign _T_4385 = {_T_4355,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@47831.4]
  assign _T_4386 = _T_4354 ? _T_4383 : _T_4385; // @[Mux.scala 31:69:@47832.4]
  assign _T_4387 = _T_4353 ? _T_4381 : _T_4386; // @[Mux.scala 31:69:@47833.4]
  assign _T_4388 = _T_4352 ? _T_4379 : _T_4387; // @[Mux.scala 31:69:@47834.4]
  assign _T_4389 = _T_4351 ? _T_4377 : _T_4388; // @[Mux.scala 31:69:@47835.4]
  assign _T_4390 = _T_4350 ? _T_4375 : _T_4389; // @[Mux.scala 31:69:@47836.4]
  assign _T_4391 = _T_4349 ? _T_4373 : _T_4390; // @[Mux.scala 31:69:@47837.4]
  assign _T_4392 = _T_4348 ? _T_4371 : _T_4391; // @[Mux.scala 31:69:@47838.4]
  assign _T_4393 = _T_4347 ? _T_4369 : _T_4392; // @[Mux.scala 31:69:@47839.4]
  assign _T_4394 = _T_4346 ? _T_4367 : _T_4393; // @[Mux.scala 31:69:@47840.4]
  assign _T_4395 = _T_4345 ? _T_4365 : _T_4394; // @[Mux.scala 31:69:@47841.4]
  assign _T_4396 = _T_4344 ? _T_4363 : _T_4395; // @[Mux.scala 31:69:@47842.4]
  assign _T_4397 = _T_4343 ? _T_4361 : _T_4396; // @[Mux.scala 31:69:@47843.4]
  assign _T_4398 = _T_4342 ? _T_4359 : _T_4397; // @[Mux.scala 31:69:@47844.4]
  assign _T_4399 = _T_4341 ? _T_4357 : _T_4398; // @[Mux.scala 31:69:@47845.4]
  assign _T_4404 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47852.4]
  assign _T_4407 = _T_4404 & _T_2886; // @[MemPrimitives.scala 110:228:@47854.4]
  assign _T_4410 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47856.4]
  assign _T_4413 = _T_4410 & _T_2892; // @[MemPrimitives.scala 110:228:@47858.4]
  assign _T_4416 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47860.4]
  assign _T_4419 = _T_4416 & _T_2898; // @[MemPrimitives.scala 110:228:@47862.4]
  assign _T_4422 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47864.4]
  assign _T_4425 = _T_4422 & _T_2904; // @[MemPrimitives.scala 110:228:@47866.4]
  assign _T_4428 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47868.4]
  assign _T_4431 = _T_4428 & _T_2910; // @[MemPrimitives.scala 110:228:@47870.4]
  assign _T_4434 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47872.4]
  assign _T_4437 = _T_4434 & _T_2916; // @[MemPrimitives.scala 110:228:@47874.4]
  assign _T_4440 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47876.4]
  assign _T_4443 = _T_4440 & _T_2922; // @[MemPrimitives.scala 110:228:@47878.4]
  assign _T_4446 = io_rPort_18_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47880.4]
  assign _T_4449 = _T_4446 & _T_2928; // @[MemPrimitives.scala 110:228:@47882.4]
  assign _T_4452 = io_rPort_20_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47884.4]
  assign _T_4455 = _T_4452 & _T_2934; // @[MemPrimitives.scala 110:228:@47886.4]
  assign _T_4458 = io_rPort_21_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47888.4]
  assign _T_4461 = _T_4458 & _T_2940; // @[MemPrimitives.scala 110:228:@47890.4]
  assign _T_4464 = io_rPort_23_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47892.4]
  assign _T_4467 = _T_4464 & _T_2946; // @[MemPrimitives.scala 110:228:@47894.4]
  assign _T_4470 = io_rPort_24_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47896.4]
  assign _T_4473 = _T_4470 & _T_2952; // @[MemPrimitives.scala 110:228:@47898.4]
  assign _T_4476 = io_rPort_25_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47900.4]
  assign _T_4479 = _T_4476 & _T_2958; // @[MemPrimitives.scala 110:228:@47902.4]
  assign _T_4482 = io_rPort_27_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47904.4]
  assign _T_4485 = _T_4482 & _T_2964; // @[MemPrimitives.scala 110:228:@47906.4]
  assign _T_4488 = io_rPort_28_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@47908.4]
  assign _T_4491 = _T_4488 & _T_2970; // @[MemPrimitives.scala 110:228:@47910.4]
  assign _T_4493 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@47930.4]
  assign _T_4494 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@47931.4]
  assign _T_4495 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@47932.4]
  assign _T_4496 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@47933.4]
  assign _T_4497 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@47934.4]
  assign _T_4498 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@47935.4]
  assign _T_4499 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@47936.4]
  assign _T_4500 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@47937.4]
  assign _T_4501 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 123:41:@47938.4]
  assign _T_4502 = StickySelects_11_io_outs_9; // @[MemPrimitives.scala 123:41:@47939.4]
  assign _T_4503 = StickySelects_11_io_outs_10; // @[MemPrimitives.scala 123:41:@47940.4]
  assign _T_4504 = StickySelects_11_io_outs_11; // @[MemPrimitives.scala 123:41:@47941.4]
  assign _T_4505 = StickySelects_11_io_outs_12; // @[MemPrimitives.scala 123:41:@47942.4]
  assign _T_4506 = StickySelects_11_io_outs_13; // @[MemPrimitives.scala 123:41:@47943.4]
  assign _T_4507 = StickySelects_11_io_outs_14; // @[MemPrimitives.scala 123:41:@47944.4]
  assign _T_4509 = {_T_4493,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@47946.4]
  assign _T_4511 = {_T_4494,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@47948.4]
  assign _T_4513 = {_T_4495,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@47950.4]
  assign _T_4515 = {_T_4496,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@47952.4]
  assign _T_4517 = {_T_4497,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@47954.4]
  assign _T_4519 = {_T_4498,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@47956.4]
  assign _T_4521 = {_T_4499,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@47958.4]
  assign _T_4523 = {_T_4500,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@47960.4]
  assign _T_4525 = {_T_4501,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@47962.4]
  assign _T_4527 = {_T_4502,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@47964.4]
  assign _T_4529 = {_T_4503,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@47966.4]
  assign _T_4531 = {_T_4504,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@47968.4]
  assign _T_4533 = {_T_4505,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@47970.4]
  assign _T_4535 = {_T_4506,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@47972.4]
  assign _T_4537 = {_T_4507,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@47974.4]
  assign _T_4538 = _T_4506 ? _T_4535 : _T_4537; // @[Mux.scala 31:69:@47975.4]
  assign _T_4539 = _T_4505 ? _T_4533 : _T_4538; // @[Mux.scala 31:69:@47976.4]
  assign _T_4540 = _T_4504 ? _T_4531 : _T_4539; // @[Mux.scala 31:69:@47977.4]
  assign _T_4541 = _T_4503 ? _T_4529 : _T_4540; // @[Mux.scala 31:69:@47978.4]
  assign _T_4542 = _T_4502 ? _T_4527 : _T_4541; // @[Mux.scala 31:69:@47979.4]
  assign _T_4543 = _T_4501 ? _T_4525 : _T_4542; // @[Mux.scala 31:69:@47980.4]
  assign _T_4544 = _T_4500 ? _T_4523 : _T_4543; // @[Mux.scala 31:69:@47981.4]
  assign _T_4545 = _T_4499 ? _T_4521 : _T_4544; // @[Mux.scala 31:69:@47982.4]
  assign _T_4546 = _T_4498 ? _T_4519 : _T_4545; // @[Mux.scala 31:69:@47983.4]
  assign _T_4547 = _T_4497 ? _T_4517 : _T_4546; // @[Mux.scala 31:69:@47984.4]
  assign _T_4548 = _T_4496 ? _T_4515 : _T_4547; // @[Mux.scala 31:69:@47985.4]
  assign _T_4549 = _T_4495 ? _T_4513 : _T_4548; // @[Mux.scala 31:69:@47986.4]
  assign _T_4550 = _T_4494 ? _T_4511 : _T_4549; // @[Mux.scala 31:69:@47987.4]
  assign _T_4551 = _T_4493 ? _T_4509 : _T_4550; // @[Mux.scala 31:69:@47988.4]
  assign _T_4559 = _T_4252 & _T_3038; // @[MemPrimitives.scala 110:228:@47997.4]
  assign _T_4565 = _T_4258 & _T_3044; // @[MemPrimitives.scala 110:228:@48001.4]
  assign _T_4571 = _T_4264 & _T_3050; // @[MemPrimitives.scala 110:228:@48005.4]
  assign _T_4577 = _T_4270 & _T_3056; // @[MemPrimitives.scala 110:228:@48009.4]
  assign _T_4583 = _T_4276 & _T_3062; // @[MemPrimitives.scala 110:228:@48013.4]
  assign _T_4589 = _T_4282 & _T_3068; // @[MemPrimitives.scala 110:228:@48017.4]
  assign _T_4595 = _T_4288 & _T_3074; // @[MemPrimitives.scala 110:228:@48021.4]
  assign _T_4601 = _T_4294 & _T_3080; // @[MemPrimitives.scala 110:228:@48025.4]
  assign _T_4607 = _T_4300 & _T_3086; // @[MemPrimitives.scala 110:228:@48029.4]
  assign _T_4613 = _T_4306 & _T_3092; // @[MemPrimitives.scala 110:228:@48033.4]
  assign _T_4619 = _T_4312 & _T_3098; // @[MemPrimitives.scala 110:228:@48037.4]
  assign _T_4625 = _T_4318 & _T_3104; // @[MemPrimitives.scala 110:228:@48041.4]
  assign _T_4631 = _T_4324 & _T_3110; // @[MemPrimitives.scala 110:228:@48045.4]
  assign _T_4637 = _T_4330 & _T_3116; // @[MemPrimitives.scala 110:228:@48049.4]
  assign _T_4643 = _T_4336 & _T_3122; // @[MemPrimitives.scala 110:228:@48053.4]
  assign _T_4645 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@48073.4]
  assign _T_4646 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@48074.4]
  assign _T_4647 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@48075.4]
  assign _T_4648 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@48076.4]
  assign _T_4649 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@48077.4]
  assign _T_4650 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@48078.4]
  assign _T_4651 = StickySelects_12_io_outs_6; // @[MemPrimitives.scala 123:41:@48079.4]
  assign _T_4652 = StickySelects_12_io_outs_7; // @[MemPrimitives.scala 123:41:@48080.4]
  assign _T_4653 = StickySelects_12_io_outs_8; // @[MemPrimitives.scala 123:41:@48081.4]
  assign _T_4654 = StickySelects_12_io_outs_9; // @[MemPrimitives.scala 123:41:@48082.4]
  assign _T_4655 = StickySelects_12_io_outs_10; // @[MemPrimitives.scala 123:41:@48083.4]
  assign _T_4656 = StickySelects_12_io_outs_11; // @[MemPrimitives.scala 123:41:@48084.4]
  assign _T_4657 = StickySelects_12_io_outs_12; // @[MemPrimitives.scala 123:41:@48085.4]
  assign _T_4658 = StickySelects_12_io_outs_13; // @[MemPrimitives.scala 123:41:@48086.4]
  assign _T_4659 = StickySelects_12_io_outs_14; // @[MemPrimitives.scala 123:41:@48087.4]
  assign _T_4661 = {_T_4645,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@48089.4]
  assign _T_4663 = {_T_4646,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@48091.4]
  assign _T_4665 = {_T_4647,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@48093.4]
  assign _T_4667 = {_T_4648,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@48095.4]
  assign _T_4669 = {_T_4649,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@48097.4]
  assign _T_4671 = {_T_4650,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@48099.4]
  assign _T_4673 = {_T_4651,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@48101.4]
  assign _T_4675 = {_T_4652,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@48103.4]
  assign _T_4677 = {_T_4653,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@48105.4]
  assign _T_4679 = {_T_4654,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@48107.4]
  assign _T_4681 = {_T_4655,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@48109.4]
  assign _T_4683 = {_T_4656,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@48111.4]
  assign _T_4685 = {_T_4657,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@48113.4]
  assign _T_4687 = {_T_4658,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@48115.4]
  assign _T_4689 = {_T_4659,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@48117.4]
  assign _T_4690 = _T_4658 ? _T_4687 : _T_4689; // @[Mux.scala 31:69:@48118.4]
  assign _T_4691 = _T_4657 ? _T_4685 : _T_4690; // @[Mux.scala 31:69:@48119.4]
  assign _T_4692 = _T_4656 ? _T_4683 : _T_4691; // @[Mux.scala 31:69:@48120.4]
  assign _T_4693 = _T_4655 ? _T_4681 : _T_4692; // @[Mux.scala 31:69:@48121.4]
  assign _T_4694 = _T_4654 ? _T_4679 : _T_4693; // @[Mux.scala 31:69:@48122.4]
  assign _T_4695 = _T_4653 ? _T_4677 : _T_4694; // @[Mux.scala 31:69:@48123.4]
  assign _T_4696 = _T_4652 ? _T_4675 : _T_4695; // @[Mux.scala 31:69:@48124.4]
  assign _T_4697 = _T_4651 ? _T_4673 : _T_4696; // @[Mux.scala 31:69:@48125.4]
  assign _T_4698 = _T_4650 ? _T_4671 : _T_4697; // @[Mux.scala 31:69:@48126.4]
  assign _T_4699 = _T_4649 ? _T_4669 : _T_4698; // @[Mux.scala 31:69:@48127.4]
  assign _T_4700 = _T_4648 ? _T_4667 : _T_4699; // @[Mux.scala 31:69:@48128.4]
  assign _T_4701 = _T_4647 ? _T_4665 : _T_4700; // @[Mux.scala 31:69:@48129.4]
  assign _T_4702 = _T_4646 ? _T_4663 : _T_4701; // @[Mux.scala 31:69:@48130.4]
  assign _T_4703 = _T_4645 ? _T_4661 : _T_4702; // @[Mux.scala 31:69:@48131.4]
  assign _T_4711 = _T_4404 & _T_3190; // @[MemPrimitives.scala 110:228:@48140.4]
  assign _T_4717 = _T_4410 & _T_3196; // @[MemPrimitives.scala 110:228:@48144.4]
  assign _T_4723 = _T_4416 & _T_3202; // @[MemPrimitives.scala 110:228:@48148.4]
  assign _T_4729 = _T_4422 & _T_3208; // @[MemPrimitives.scala 110:228:@48152.4]
  assign _T_4735 = _T_4428 & _T_3214; // @[MemPrimitives.scala 110:228:@48156.4]
  assign _T_4741 = _T_4434 & _T_3220; // @[MemPrimitives.scala 110:228:@48160.4]
  assign _T_4747 = _T_4440 & _T_3226; // @[MemPrimitives.scala 110:228:@48164.4]
  assign _T_4753 = _T_4446 & _T_3232; // @[MemPrimitives.scala 110:228:@48168.4]
  assign _T_4759 = _T_4452 & _T_3238; // @[MemPrimitives.scala 110:228:@48172.4]
  assign _T_4765 = _T_4458 & _T_3244; // @[MemPrimitives.scala 110:228:@48176.4]
  assign _T_4771 = _T_4464 & _T_3250; // @[MemPrimitives.scala 110:228:@48180.4]
  assign _T_4777 = _T_4470 & _T_3256; // @[MemPrimitives.scala 110:228:@48184.4]
  assign _T_4783 = _T_4476 & _T_3262; // @[MemPrimitives.scala 110:228:@48188.4]
  assign _T_4789 = _T_4482 & _T_3268; // @[MemPrimitives.scala 110:228:@48192.4]
  assign _T_4795 = _T_4488 & _T_3274; // @[MemPrimitives.scala 110:228:@48196.4]
  assign _T_4797 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@48216.4]
  assign _T_4798 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@48217.4]
  assign _T_4799 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@48218.4]
  assign _T_4800 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@48219.4]
  assign _T_4801 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@48220.4]
  assign _T_4802 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@48221.4]
  assign _T_4803 = StickySelects_13_io_outs_6; // @[MemPrimitives.scala 123:41:@48222.4]
  assign _T_4804 = StickySelects_13_io_outs_7; // @[MemPrimitives.scala 123:41:@48223.4]
  assign _T_4805 = StickySelects_13_io_outs_8; // @[MemPrimitives.scala 123:41:@48224.4]
  assign _T_4806 = StickySelects_13_io_outs_9; // @[MemPrimitives.scala 123:41:@48225.4]
  assign _T_4807 = StickySelects_13_io_outs_10; // @[MemPrimitives.scala 123:41:@48226.4]
  assign _T_4808 = StickySelects_13_io_outs_11; // @[MemPrimitives.scala 123:41:@48227.4]
  assign _T_4809 = StickySelects_13_io_outs_12; // @[MemPrimitives.scala 123:41:@48228.4]
  assign _T_4810 = StickySelects_13_io_outs_13; // @[MemPrimitives.scala 123:41:@48229.4]
  assign _T_4811 = StickySelects_13_io_outs_14; // @[MemPrimitives.scala 123:41:@48230.4]
  assign _T_4813 = {_T_4797,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@48232.4]
  assign _T_4815 = {_T_4798,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@48234.4]
  assign _T_4817 = {_T_4799,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@48236.4]
  assign _T_4819 = {_T_4800,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@48238.4]
  assign _T_4821 = {_T_4801,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@48240.4]
  assign _T_4823 = {_T_4802,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@48242.4]
  assign _T_4825 = {_T_4803,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@48244.4]
  assign _T_4827 = {_T_4804,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@48246.4]
  assign _T_4829 = {_T_4805,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@48248.4]
  assign _T_4831 = {_T_4806,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@48250.4]
  assign _T_4833 = {_T_4807,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@48252.4]
  assign _T_4835 = {_T_4808,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@48254.4]
  assign _T_4837 = {_T_4809,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@48256.4]
  assign _T_4839 = {_T_4810,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@48258.4]
  assign _T_4841 = {_T_4811,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@48260.4]
  assign _T_4842 = _T_4810 ? _T_4839 : _T_4841; // @[Mux.scala 31:69:@48261.4]
  assign _T_4843 = _T_4809 ? _T_4837 : _T_4842; // @[Mux.scala 31:69:@48262.4]
  assign _T_4844 = _T_4808 ? _T_4835 : _T_4843; // @[Mux.scala 31:69:@48263.4]
  assign _T_4845 = _T_4807 ? _T_4833 : _T_4844; // @[Mux.scala 31:69:@48264.4]
  assign _T_4846 = _T_4806 ? _T_4831 : _T_4845; // @[Mux.scala 31:69:@48265.4]
  assign _T_4847 = _T_4805 ? _T_4829 : _T_4846; // @[Mux.scala 31:69:@48266.4]
  assign _T_4848 = _T_4804 ? _T_4827 : _T_4847; // @[Mux.scala 31:69:@48267.4]
  assign _T_4849 = _T_4803 ? _T_4825 : _T_4848; // @[Mux.scala 31:69:@48268.4]
  assign _T_4850 = _T_4802 ? _T_4823 : _T_4849; // @[Mux.scala 31:69:@48269.4]
  assign _T_4851 = _T_4801 ? _T_4821 : _T_4850; // @[Mux.scala 31:69:@48270.4]
  assign _T_4852 = _T_4800 ? _T_4819 : _T_4851; // @[Mux.scala 31:69:@48271.4]
  assign _T_4853 = _T_4799 ? _T_4817 : _T_4852; // @[Mux.scala 31:69:@48272.4]
  assign _T_4854 = _T_4798 ? _T_4815 : _T_4853; // @[Mux.scala 31:69:@48273.4]
  assign _T_4855 = _T_4797 ? _T_4813 : _T_4854; // @[Mux.scala 31:69:@48274.4]
  assign _T_4863 = _T_4252 & _T_3342; // @[MemPrimitives.scala 110:228:@48283.4]
  assign _T_4869 = _T_4258 & _T_3348; // @[MemPrimitives.scala 110:228:@48287.4]
  assign _T_4875 = _T_4264 & _T_3354; // @[MemPrimitives.scala 110:228:@48291.4]
  assign _T_4881 = _T_4270 & _T_3360; // @[MemPrimitives.scala 110:228:@48295.4]
  assign _T_4887 = _T_4276 & _T_3366; // @[MemPrimitives.scala 110:228:@48299.4]
  assign _T_4893 = _T_4282 & _T_3372; // @[MemPrimitives.scala 110:228:@48303.4]
  assign _T_4899 = _T_4288 & _T_3378; // @[MemPrimitives.scala 110:228:@48307.4]
  assign _T_4905 = _T_4294 & _T_3384; // @[MemPrimitives.scala 110:228:@48311.4]
  assign _T_4911 = _T_4300 & _T_3390; // @[MemPrimitives.scala 110:228:@48315.4]
  assign _T_4917 = _T_4306 & _T_3396; // @[MemPrimitives.scala 110:228:@48319.4]
  assign _T_4923 = _T_4312 & _T_3402; // @[MemPrimitives.scala 110:228:@48323.4]
  assign _T_4929 = _T_4318 & _T_3408; // @[MemPrimitives.scala 110:228:@48327.4]
  assign _T_4935 = _T_4324 & _T_3414; // @[MemPrimitives.scala 110:228:@48331.4]
  assign _T_4941 = _T_4330 & _T_3420; // @[MemPrimitives.scala 110:228:@48335.4]
  assign _T_4947 = _T_4336 & _T_3426; // @[MemPrimitives.scala 110:228:@48339.4]
  assign _T_4949 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@48359.4]
  assign _T_4950 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@48360.4]
  assign _T_4951 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@48361.4]
  assign _T_4952 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@48362.4]
  assign _T_4953 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@48363.4]
  assign _T_4954 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@48364.4]
  assign _T_4955 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 123:41:@48365.4]
  assign _T_4956 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 123:41:@48366.4]
  assign _T_4957 = StickySelects_14_io_outs_8; // @[MemPrimitives.scala 123:41:@48367.4]
  assign _T_4958 = StickySelects_14_io_outs_9; // @[MemPrimitives.scala 123:41:@48368.4]
  assign _T_4959 = StickySelects_14_io_outs_10; // @[MemPrimitives.scala 123:41:@48369.4]
  assign _T_4960 = StickySelects_14_io_outs_11; // @[MemPrimitives.scala 123:41:@48370.4]
  assign _T_4961 = StickySelects_14_io_outs_12; // @[MemPrimitives.scala 123:41:@48371.4]
  assign _T_4962 = StickySelects_14_io_outs_13; // @[MemPrimitives.scala 123:41:@48372.4]
  assign _T_4963 = StickySelects_14_io_outs_14; // @[MemPrimitives.scala 123:41:@48373.4]
  assign _T_4965 = {_T_4949,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@48375.4]
  assign _T_4967 = {_T_4950,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@48377.4]
  assign _T_4969 = {_T_4951,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@48379.4]
  assign _T_4971 = {_T_4952,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@48381.4]
  assign _T_4973 = {_T_4953,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@48383.4]
  assign _T_4975 = {_T_4954,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@48385.4]
  assign _T_4977 = {_T_4955,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@48387.4]
  assign _T_4979 = {_T_4956,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@48389.4]
  assign _T_4981 = {_T_4957,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@48391.4]
  assign _T_4983 = {_T_4958,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@48393.4]
  assign _T_4985 = {_T_4959,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@48395.4]
  assign _T_4987 = {_T_4960,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@48397.4]
  assign _T_4989 = {_T_4961,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@48399.4]
  assign _T_4991 = {_T_4962,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@48401.4]
  assign _T_4993 = {_T_4963,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@48403.4]
  assign _T_4994 = _T_4962 ? _T_4991 : _T_4993; // @[Mux.scala 31:69:@48404.4]
  assign _T_4995 = _T_4961 ? _T_4989 : _T_4994; // @[Mux.scala 31:69:@48405.4]
  assign _T_4996 = _T_4960 ? _T_4987 : _T_4995; // @[Mux.scala 31:69:@48406.4]
  assign _T_4997 = _T_4959 ? _T_4985 : _T_4996; // @[Mux.scala 31:69:@48407.4]
  assign _T_4998 = _T_4958 ? _T_4983 : _T_4997; // @[Mux.scala 31:69:@48408.4]
  assign _T_4999 = _T_4957 ? _T_4981 : _T_4998; // @[Mux.scala 31:69:@48409.4]
  assign _T_5000 = _T_4956 ? _T_4979 : _T_4999; // @[Mux.scala 31:69:@48410.4]
  assign _T_5001 = _T_4955 ? _T_4977 : _T_5000; // @[Mux.scala 31:69:@48411.4]
  assign _T_5002 = _T_4954 ? _T_4975 : _T_5001; // @[Mux.scala 31:69:@48412.4]
  assign _T_5003 = _T_4953 ? _T_4973 : _T_5002; // @[Mux.scala 31:69:@48413.4]
  assign _T_5004 = _T_4952 ? _T_4971 : _T_5003; // @[Mux.scala 31:69:@48414.4]
  assign _T_5005 = _T_4951 ? _T_4969 : _T_5004; // @[Mux.scala 31:69:@48415.4]
  assign _T_5006 = _T_4950 ? _T_4967 : _T_5005; // @[Mux.scala 31:69:@48416.4]
  assign _T_5007 = _T_4949 ? _T_4965 : _T_5006; // @[Mux.scala 31:69:@48417.4]
  assign _T_5015 = _T_4404 & _T_3494; // @[MemPrimitives.scala 110:228:@48426.4]
  assign _T_5021 = _T_4410 & _T_3500; // @[MemPrimitives.scala 110:228:@48430.4]
  assign _T_5027 = _T_4416 & _T_3506; // @[MemPrimitives.scala 110:228:@48434.4]
  assign _T_5033 = _T_4422 & _T_3512; // @[MemPrimitives.scala 110:228:@48438.4]
  assign _T_5039 = _T_4428 & _T_3518; // @[MemPrimitives.scala 110:228:@48442.4]
  assign _T_5045 = _T_4434 & _T_3524; // @[MemPrimitives.scala 110:228:@48446.4]
  assign _T_5051 = _T_4440 & _T_3530; // @[MemPrimitives.scala 110:228:@48450.4]
  assign _T_5057 = _T_4446 & _T_3536; // @[MemPrimitives.scala 110:228:@48454.4]
  assign _T_5063 = _T_4452 & _T_3542; // @[MemPrimitives.scala 110:228:@48458.4]
  assign _T_5069 = _T_4458 & _T_3548; // @[MemPrimitives.scala 110:228:@48462.4]
  assign _T_5075 = _T_4464 & _T_3554; // @[MemPrimitives.scala 110:228:@48466.4]
  assign _T_5081 = _T_4470 & _T_3560; // @[MemPrimitives.scala 110:228:@48470.4]
  assign _T_5087 = _T_4476 & _T_3566; // @[MemPrimitives.scala 110:228:@48474.4]
  assign _T_5093 = _T_4482 & _T_3572; // @[MemPrimitives.scala 110:228:@48478.4]
  assign _T_5099 = _T_4488 & _T_3578; // @[MemPrimitives.scala 110:228:@48482.4]
  assign _T_5101 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@48502.4]
  assign _T_5102 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@48503.4]
  assign _T_5103 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@48504.4]
  assign _T_5104 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@48505.4]
  assign _T_5105 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@48506.4]
  assign _T_5106 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@48507.4]
  assign _T_5107 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 123:41:@48508.4]
  assign _T_5108 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 123:41:@48509.4]
  assign _T_5109 = StickySelects_15_io_outs_8; // @[MemPrimitives.scala 123:41:@48510.4]
  assign _T_5110 = StickySelects_15_io_outs_9; // @[MemPrimitives.scala 123:41:@48511.4]
  assign _T_5111 = StickySelects_15_io_outs_10; // @[MemPrimitives.scala 123:41:@48512.4]
  assign _T_5112 = StickySelects_15_io_outs_11; // @[MemPrimitives.scala 123:41:@48513.4]
  assign _T_5113 = StickySelects_15_io_outs_12; // @[MemPrimitives.scala 123:41:@48514.4]
  assign _T_5114 = StickySelects_15_io_outs_13; // @[MemPrimitives.scala 123:41:@48515.4]
  assign _T_5115 = StickySelects_15_io_outs_14; // @[MemPrimitives.scala 123:41:@48516.4]
  assign _T_5117 = {_T_5101,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@48518.4]
  assign _T_5119 = {_T_5102,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@48520.4]
  assign _T_5121 = {_T_5103,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@48522.4]
  assign _T_5123 = {_T_5104,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@48524.4]
  assign _T_5125 = {_T_5105,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@48526.4]
  assign _T_5127 = {_T_5106,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@48528.4]
  assign _T_5129 = {_T_5107,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@48530.4]
  assign _T_5131 = {_T_5108,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@48532.4]
  assign _T_5133 = {_T_5109,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@48534.4]
  assign _T_5135 = {_T_5110,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@48536.4]
  assign _T_5137 = {_T_5111,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@48538.4]
  assign _T_5139 = {_T_5112,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@48540.4]
  assign _T_5141 = {_T_5113,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@48542.4]
  assign _T_5143 = {_T_5114,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@48544.4]
  assign _T_5145 = {_T_5115,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@48546.4]
  assign _T_5146 = _T_5114 ? _T_5143 : _T_5145; // @[Mux.scala 31:69:@48547.4]
  assign _T_5147 = _T_5113 ? _T_5141 : _T_5146; // @[Mux.scala 31:69:@48548.4]
  assign _T_5148 = _T_5112 ? _T_5139 : _T_5147; // @[Mux.scala 31:69:@48549.4]
  assign _T_5149 = _T_5111 ? _T_5137 : _T_5148; // @[Mux.scala 31:69:@48550.4]
  assign _T_5150 = _T_5110 ? _T_5135 : _T_5149; // @[Mux.scala 31:69:@48551.4]
  assign _T_5151 = _T_5109 ? _T_5133 : _T_5150; // @[Mux.scala 31:69:@48552.4]
  assign _T_5152 = _T_5108 ? _T_5131 : _T_5151; // @[Mux.scala 31:69:@48553.4]
  assign _T_5153 = _T_5107 ? _T_5129 : _T_5152; // @[Mux.scala 31:69:@48554.4]
  assign _T_5154 = _T_5106 ? _T_5127 : _T_5153; // @[Mux.scala 31:69:@48555.4]
  assign _T_5155 = _T_5105 ? _T_5125 : _T_5154; // @[Mux.scala 31:69:@48556.4]
  assign _T_5156 = _T_5104 ? _T_5123 : _T_5155; // @[Mux.scala 31:69:@48557.4]
  assign _T_5157 = _T_5103 ? _T_5121 : _T_5156; // @[Mux.scala 31:69:@48558.4]
  assign _T_5158 = _T_5102 ? _T_5119 : _T_5157; // @[Mux.scala 31:69:@48559.4]
  assign _T_5159 = _T_5101 ? _T_5117 : _T_5158; // @[Mux.scala 31:69:@48560.4]
  assign _T_5167 = _T_4252 & _T_3646; // @[MemPrimitives.scala 110:228:@48569.4]
  assign _T_5173 = _T_4258 & _T_3652; // @[MemPrimitives.scala 110:228:@48573.4]
  assign _T_5179 = _T_4264 & _T_3658; // @[MemPrimitives.scala 110:228:@48577.4]
  assign _T_5185 = _T_4270 & _T_3664; // @[MemPrimitives.scala 110:228:@48581.4]
  assign _T_5191 = _T_4276 & _T_3670; // @[MemPrimitives.scala 110:228:@48585.4]
  assign _T_5197 = _T_4282 & _T_3676; // @[MemPrimitives.scala 110:228:@48589.4]
  assign _T_5203 = _T_4288 & _T_3682; // @[MemPrimitives.scala 110:228:@48593.4]
  assign _T_5209 = _T_4294 & _T_3688; // @[MemPrimitives.scala 110:228:@48597.4]
  assign _T_5215 = _T_4300 & _T_3694; // @[MemPrimitives.scala 110:228:@48601.4]
  assign _T_5221 = _T_4306 & _T_3700; // @[MemPrimitives.scala 110:228:@48605.4]
  assign _T_5227 = _T_4312 & _T_3706; // @[MemPrimitives.scala 110:228:@48609.4]
  assign _T_5233 = _T_4318 & _T_3712; // @[MemPrimitives.scala 110:228:@48613.4]
  assign _T_5239 = _T_4324 & _T_3718; // @[MemPrimitives.scala 110:228:@48617.4]
  assign _T_5245 = _T_4330 & _T_3724; // @[MemPrimitives.scala 110:228:@48621.4]
  assign _T_5251 = _T_4336 & _T_3730; // @[MemPrimitives.scala 110:228:@48625.4]
  assign _T_5253 = StickySelects_16_io_outs_0; // @[MemPrimitives.scala 123:41:@48645.4]
  assign _T_5254 = StickySelects_16_io_outs_1; // @[MemPrimitives.scala 123:41:@48646.4]
  assign _T_5255 = StickySelects_16_io_outs_2; // @[MemPrimitives.scala 123:41:@48647.4]
  assign _T_5256 = StickySelects_16_io_outs_3; // @[MemPrimitives.scala 123:41:@48648.4]
  assign _T_5257 = StickySelects_16_io_outs_4; // @[MemPrimitives.scala 123:41:@48649.4]
  assign _T_5258 = StickySelects_16_io_outs_5; // @[MemPrimitives.scala 123:41:@48650.4]
  assign _T_5259 = StickySelects_16_io_outs_6; // @[MemPrimitives.scala 123:41:@48651.4]
  assign _T_5260 = StickySelects_16_io_outs_7; // @[MemPrimitives.scala 123:41:@48652.4]
  assign _T_5261 = StickySelects_16_io_outs_8; // @[MemPrimitives.scala 123:41:@48653.4]
  assign _T_5262 = StickySelects_16_io_outs_9; // @[MemPrimitives.scala 123:41:@48654.4]
  assign _T_5263 = StickySelects_16_io_outs_10; // @[MemPrimitives.scala 123:41:@48655.4]
  assign _T_5264 = StickySelects_16_io_outs_11; // @[MemPrimitives.scala 123:41:@48656.4]
  assign _T_5265 = StickySelects_16_io_outs_12; // @[MemPrimitives.scala 123:41:@48657.4]
  assign _T_5266 = StickySelects_16_io_outs_13; // @[MemPrimitives.scala 123:41:@48658.4]
  assign _T_5267 = StickySelects_16_io_outs_14; // @[MemPrimitives.scala 123:41:@48659.4]
  assign _T_5269 = {_T_5253,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@48661.4]
  assign _T_5271 = {_T_5254,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@48663.4]
  assign _T_5273 = {_T_5255,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@48665.4]
  assign _T_5275 = {_T_5256,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@48667.4]
  assign _T_5277 = {_T_5257,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@48669.4]
  assign _T_5279 = {_T_5258,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@48671.4]
  assign _T_5281 = {_T_5259,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@48673.4]
  assign _T_5283 = {_T_5260,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@48675.4]
  assign _T_5285 = {_T_5261,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@48677.4]
  assign _T_5287 = {_T_5262,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@48679.4]
  assign _T_5289 = {_T_5263,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@48681.4]
  assign _T_5291 = {_T_5264,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@48683.4]
  assign _T_5293 = {_T_5265,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@48685.4]
  assign _T_5295 = {_T_5266,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@48687.4]
  assign _T_5297 = {_T_5267,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@48689.4]
  assign _T_5298 = _T_5266 ? _T_5295 : _T_5297; // @[Mux.scala 31:69:@48690.4]
  assign _T_5299 = _T_5265 ? _T_5293 : _T_5298; // @[Mux.scala 31:69:@48691.4]
  assign _T_5300 = _T_5264 ? _T_5291 : _T_5299; // @[Mux.scala 31:69:@48692.4]
  assign _T_5301 = _T_5263 ? _T_5289 : _T_5300; // @[Mux.scala 31:69:@48693.4]
  assign _T_5302 = _T_5262 ? _T_5287 : _T_5301; // @[Mux.scala 31:69:@48694.4]
  assign _T_5303 = _T_5261 ? _T_5285 : _T_5302; // @[Mux.scala 31:69:@48695.4]
  assign _T_5304 = _T_5260 ? _T_5283 : _T_5303; // @[Mux.scala 31:69:@48696.4]
  assign _T_5305 = _T_5259 ? _T_5281 : _T_5304; // @[Mux.scala 31:69:@48697.4]
  assign _T_5306 = _T_5258 ? _T_5279 : _T_5305; // @[Mux.scala 31:69:@48698.4]
  assign _T_5307 = _T_5257 ? _T_5277 : _T_5306; // @[Mux.scala 31:69:@48699.4]
  assign _T_5308 = _T_5256 ? _T_5275 : _T_5307; // @[Mux.scala 31:69:@48700.4]
  assign _T_5309 = _T_5255 ? _T_5273 : _T_5308; // @[Mux.scala 31:69:@48701.4]
  assign _T_5310 = _T_5254 ? _T_5271 : _T_5309; // @[Mux.scala 31:69:@48702.4]
  assign _T_5311 = _T_5253 ? _T_5269 : _T_5310; // @[Mux.scala 31:69:@48703.4]
  assign _T_5319 = _T_4404 & _T_3798; // @[MemPrimitives.scala 110:228:@48712.4]
  assign _T_5325 = _T_4410 & _T_3804; // @[MemPrimitives.scala 110:228:@48716.4]
  assign _T_5331 = _T_4416 & _T_3810; // @[MemPrimitives.scala 110:228:@48720.4]
  assign _T_5337 = _T_4422 & _T_3816; // @[MemPrimitives.scala 110:228:@48724.4]
  assign _T_5343 = _T_4428 & _T_3822; // @[MemPrimitives.scala 110:228:@48728.4]
  assign _T_5349 = _T_4434 & _T_3828; // @[MemPrimitives.scala 110:228:@48732.4]
  assign _T_5355 = _T_4440 & _T_3834; // @[MemPrimitives.scala 110:228:@48736.4]
  assign _T_5361 = _T_4446 & _T_3840; // @[MemPrimitives.scala 110:228:@48740.4]
  assign _T_5367 = _T_4452 & _T_3846; // @[MemPrimitives.scala 110:228:@48744.4]
  assign _T_5373 = _T_4458 & _T_3852; // @[MemPrimitives.scala 110:228:@48748.4]
  assign _T_5379 = _T_4464 & _T_3858; // @[MemPrimitives.scala 110:228:@48752.4]
  assign _T_5385 = _T_4470 & _T_3864; // @[MemPrimitives.scala 110:228:@48756.4]
  assign _T_5391 = _T_4476 & _T_3870; // @[MemPrimitives.scala 110:228:@48760.4]
  assign _T_5397 = _T_4482 & _T_3876; // @[MemPrimitives.scala 110:228:@48764.4]
  assign _T_5403 = _T_4488 & _T_3882; // @[MemPrimitives.scala 110:228:@48768.4]
  assign _T_5405 = StickySelects_17_io_outs_0; // @[MemPrimitives.scala 123:41:@48788.4]
  assign _T_5406 = StickySelects_17_io_outs_1; // @[MemPrimitives.scala 123:41:@48789.4]
  assign _T_5407 = StickySelects_17_io_outs_2; // @[MemPrimitives.scala 123:41:@48790.4]
  assign _T_5408 = StickySelects_17_io_outs_3; // @[MemPrimitives.scala 123:41:@48791.4]
  assign _T_5409 = StickySelects_17_io_outs_4; // @[MemPrimitives.scala 123:41:@48792.4]
  assign _T_5410 = StickySelects_17_io_outs_5; // @[MemPrimitives.scala 123:41:@48793.4]
  assign _T_5411 = StickySelects_17_io_outs_6; // @[MemPrimitives.scala 123:41:@48794.4]
  assign _T_5412 = StickySelects_17_io_outs_7; // @[MemPrimitives.scala 123:41:@48795.4]
  assign _T_5413 = StickySelects_17_io_outs_8; // @[MemPrimitives.scala 123:41:@48796.4]
  assign _T_5414 = StickySelects_17_io_outs_9; // @[MemPrimitives.scala 123:41:@48797.4]
  assign _T_5415 = StickySelects_17_io_outs_10; // @[MemPrimitives.scala 123:41:@48798.4]
  assign _T_5416 = StickySelects_17_io_outs_11; // @[MemPrimitives.scala 123:41:@48799.4]
  assign _T_5417 = StickySelects_17_io_outs_12; // @[MemPrimitives.scala 123:41:@48800.4]
  assign _T_5418 = StickySelects_17_io_outs_13; // @[MemPrimitives.scala 123:41:@48801.4]
  assign _T_5419 = StickySelects_17_io_outs_14; // @[MemPrimitives.scala 123:41:@48802.4]
  assign _T_5421 = {_T_5405,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@48804.4]
  assign _T_5423 = {_T_5406,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@48806.4]
  assign _T_5425 = {_T_5407,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@48808.4]
  assign _T_5427 = {_T_5408,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@48810.4]
  assign _T_5429 = {_T_5409,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@48812.4]
  assign _T_5431 = {_T_5410,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@48814.4]
  assign _T_5433 = {_T_5411,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@48816.4]
  assign _T_5435 = {_T_5412,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@48818.4]
  assign _T_5437 = {_T_5413,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@48820.4]
  assign _T_5439 = {_T_5414,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@48822.4]
  assign _T_5441 = {_T_5415,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@48824.4]
  assign _T_5443 = {_T_5416,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@48826.4]
  assign _T_5445 = {_T_5417,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@48828.4]
  assign _T_5447 = {_T_5418,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@48830.4]
  assign _T_5449 = {_T_5419,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@48832.4]
  assign _T_5450 = _T_5418 ? _T_5447 : _T_5449; // @[Mux.scala 31:69:@48833.4]
  assign _T_5451 = _T_5417 ? _T_5445 : _T_5450; // @[Mux.scala 31:69:@48834.4]
  assign _T_5452 = _T_5416 ? _T_5443 : _T_5451; // @[Mux.scala 31:69:@48835.4]
  assign _T_5453 = _T_5415 ? _T_5441 : _T_5452; // @[Mux.scala 31:69:@48836.4]
  assign _T_5454 = _T_5414 ? _T_5439 : _T_5453; // @[Mux.scala 31:69:@48837.4]
  assign _T_5455 = _T_5413 ? _T_5437 : _T_5454; // @[Mux.scala 31:69:@48838.4]
  assign _T_5456 = _T_5412 ? _T_5435 : _T_5455; // @[Mux.scala 31:69:@48839.4]
  assign _T_5457 = _T_5411 ? _T_5433 : _T_5456; // @[Mux.scala 31:69:@48840.4]
  assign _T_5458 = _T_5410 ? _T_5431 : _T_5457; // @[Mux.scala 31:69:@48841.4]
  assign _T_5459 = _T_5409 ? _T_5429 : _T_5458; // @[Mux.scala 31:69:@48842.4]
  assign _T_5460 = _T_5408 ? _T_5427 : _T_5459; // @[Mux.scala 31:69:@48843.4]
  assign _T_5461 = _T_5407 ? _T_5425 : _T_5460; // @[Mux.scala 31:69:@48844.4]
  assign _T_5462 = _T_5406 ? _T_5423 : _T_5461; // @[Mux.scala 31:69:@48845.4]
  assign _T_5463 = _T_5405 ? _T_5421 : _T_5462; // @[Mux.scala 31:69:@48846.4]
  assign _T_5471 = _T_4252 & _T_3950; // @[MemPrimitives.scala 110:228:@48855.4]
  assign _T_5477 = _T_4258 & _T_3956; // @[MemPrimitives.scala 110:228:@48859.4]
  assign _T_5483 = _T_4264 & _T_3962; // @[MemPrimitives.scala 110:228:@48863.4]
  assign _T_5489 = _T_4270 & _T_3968; // @[MemPrimitives.scala 110:228:@48867.4]
  assign _T_5495 = _T_4276 & _T_3974; // @[MemPrimitives.scala 110:228:@48871.4]
  assign _T_5501 = _T_4282 & _T_3980; // @[MemPrimitives.scala 110:228:@48875.4]
  assign _T_5507 = _T_4288 & _T_3986; // @[MemPrimitives.scala 110:228:@48879.4]
  assign _T_5513 = _T_4294 & _T_3992; // @[MemPrimitives.scala 110:228:@48883.4]
  assign _T_5519 = _T_4300 & _T_3998; // @[MemPrimitives.scala 110:228:@48887.4]
  assign _T_5525 = _T_4306 & _T_4004; // @[MemPrimitives.scala 110:228:@48891.4]
  assign _T_5531 = _T_4312 & _T_4010; // @[MemPrimitives.scala 110:228:@48895.4]
  assign _T_5537 = _T_4318 & _T_4016; // @[MemPrimitives.scala 110:228:@48899.4]
  assign _T_5543 = _T_4324 & _T_4022; // @[MemPrimitives.scala 110:228:@48903.4]
  assign _T_5549 = _T_4330 & _T_4028; // @[MemPrimitives.scala 110:228:@48907.4]
  assign _T_5555 = _T_4336 & _T_4034; // @[MemPrimitives.scala 110:228:@48911.4]
  assign _T_5557 = StickySelects_18_io_outs_0; // @[MemPrimitives.scala 123:41:@48931.4]
  assign _T_5558 = StickySelects_18_io_outs_1; // @[MemPrimitives.scala 123:41:@48932.4]
  assign _T_5559 = StickySelects_18_io_outs_2; // @[MemPrimitives.scala 123:41:@48933.4]
  assign _T_5560 = StickySelects_18_io_outs_3; // @[MemPrimitives.scala 123:41:@48934.4]
  assign _T_5561 = StickySelects_18_io_outs_4; // @[MemPrimitives.scala 123:41:@48935.4]
  assign _T_5562 = StickySelects_18_io_outs_5; // @[MemPrimitives.scala 123:41:@48936.4]
  assign _T_5563 = StickySelects_18_io_outs_6; // @[MemPrimitives.scala 123:41:@48937.4]
  assign _T_5564 = StickySelects_18_io_outs_7; // @[MemPrimitives.scala 123:41:@48938.4]
  assign _T_5565 = StickySelects_18_io_outs_8; // @[MemPrimitives.scala 123:41:@48939.4]
  assign _T_5566 = StickySelects_18_io_outs_9; // @[MemPrimitives.scala 123:41:@48940.4]
  assign _T_5567 = StickySelects_18_io_outs_10; // @[MemPrimitives.scala 123:41:@48941.4]
  assign _T_5568 = StickySelects_18_io_outs_11; // @[MemPrimitives.scala 123:41:@48942.4]
  assign _T_5569 = StickySelects_18_io_outs_12; // @[MemPrimitives.scala 123:41:@48943.4]
  assign _T_5570 = StickySelects_18_io_outs_13; // @[MemPrimitives.scala 123:41:@48944.4]
  assign _T_5571 = StickySelects_18_io_outs_14; // @[MemPrimitives.scala 123:41:@48945.4]
  assign _T_5573 = {_T_5557,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@48947.4]
  assign _T_5575 = {_T_5558,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@48949.4]
  assign _T_5577 = {_T_5559,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@48951.4]
  assign _T_5579 = {_T_5560,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@48953.4]
  assign _T_5581 = {_T_5561,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@48955.4]
  assign _T_5583 = {_T_5562,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@48957.4]
  assign _T_5585 = {_T_5563,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@48959.4]
  assign _T_5587 = {_T_5564,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@48961.4]
  assign _T_5589 = {_T_5565,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@48963.4]
  assign _T_5591 = {_T_5566,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@48965.4]
  assign _T_5593 = {_T_5567,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@48967.4]
  assign _T_5595 = {_T_5568,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@48969.4]
  assign _T_5597 = {_T_5569,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@48971.4]
  assign _T_5599 = {_T_5570,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@48973.4]
  assign _T_5601 = {_T_5571,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@48975.4]
  assign _T_5602 = _T_5570 ? _T_5599 : _T_5601; // @[Mux.scala 31:69:@48976.4]
  assign _T_5603 = _T_5569 ? _T_5597 : _T_5602; // @[Mux.scala 31:69:@48977.4]
  assign _T_5604 = _T_5568 ? _T_5595 : _T_5603; // @[Mux.scala 31:69:@48978.4]
  assign _T_5605 = _T_5567 ? _T_5593 : _T_5604; // @[Mux.scala 31:69:@48979.4]
  assign _T_5606 = _T_5566 ? _T_5591 : _T_5605; // @[Mux.scala 31:69:@48980.4]
  assign _T_5607 = _T_5565 ? _T_5589 : _T_5606; // @[Mux.scala 31:69:@48981.4]
  assign _T_5608 = _T_5564 ? _T_5587 : _T_5607; // @[Mux.scala 31:69:@48982.4]
  assign _T_5609 = _T_5563 ? _T_5585 : _T_5608; // @[Mux.scala 31:69:@48983.4]
  assign _T_5610 = _T_5562 ? _T_5583 : _T_5609; // @[Mux.scala 31:69:@48984.4]
  assign _T_5611 = _T_5561 ? _T_5581 : _T_5610; // @[Mux.scala 31:69:@48985.4]
  assign _T_5612 = _T_5560 ? _T_5579 : _T_5611; // @[Mux.scala 31:69:@48986.4]
  assign _T_5613 = _T_5559 ? _T_5577 : _T_5612; // @[Mux.scala 31:69:@48987.4]
  assign _T_5614 = _T_5558 ? _T_5575 : _T_5613; // @[Mux.scala 31:69:@48988.4]
  assign _T_5615 = _T_5557 ? _T_5573 : _T_5614; // @[Mux.scala 31:69:@48989.4]
  assign _T_5623 = _T_4404 & _T_4102; // @[MemPrimitives.scala 110:228:@48998.4]
  assign _T_5629 = _T_4410 & _T_4108; // @[MemPrimitives.scala 110:228:@49002.4]
  assign _T_5635 = _T_4416 & _T_4114; // @[MemPrimitives.scala 110:228:@49006.4]
  assign _T_5641 = _T_4422 & _T_4120; // @[MemPrimitives.scala 110:228:@49010.4]
  assign _T_5647 = _T_4428 & _T_4126; // @[MemPrimitives.scala 110:228:@49014.4]
  assign _T_5653 = _T_4434 & _T_4132; // @[MemPrimitives.scala 110:228:@49018.4]
  assign _T_5659 = _T_4440 & _T_4138; // @[MemPrimitives.scala 110:228:@49022.4]
  assign _T_5665 = _T_4446 & _T_4144; // @[MemPrimitives.scala 110:228:@49026.4]
  assign _T_5671 = _T_4452 & _T_4150; // @[MemPrimitives.scala 110:228:@49030.4]
  assign _T_5677 = _T_4458 & _T_4156; // @[MemPrimitives.scala 110:228:@49034.4]
  assign _T_5683 = _T_4464 & _T_4162; // @[MemPrimitives.scala 110:228:@49038.4]
  assign _T_5689 = _T_4470 & _T_4168; // @[MemPrimitives.scala 110:228:@49042.4]
  assign _T_5695 = _T_4476 & _T_4174; // @[MemPrimitives.scala 110:228:@49046.4]
  assign _T_5701 = _T_4482 & _T_4180; // @[MemPrimitives.scala 110:228:@49050.4]
  assign _T_5707 = _T_4488 & _T_4186; // @[MemPrimitives.scala 110:228:@49054.4]
  assign _T_5709 = StickySelects_19_io_outs_0; // @[MemPrimitives.scala 123:41:@49074.4]
  assign _T_5710 = StickySelects_19_io_outs_1; // @[MemPrimitives.scala 123:41:@49075.4]
  assign _T_5711 = StickySelects_19_io_outs_2; // @[MemPrimitives.scala 123:41:@49076.4]
  assign _T_5712 = StickySelects_19_io_outs_3; // @[MemPrimitives.scala 123:41:@49077.4]
  assign _T_5713 = StickySelects_19_io_outs_4; // @[MemPrimitives.scala 123:41:@49078.4]
  assign _T_5714 = StickySelects_19_io_outs_5; // @[MemPrimitives.scala 123:41:@49079.4]
  assign _T_5715 = StickySelects_19_io_outs_6; // @[MemPrimitives.scala 123:41:@49080.4]
  assign _T_5716 = StickySelects_19_io_outs_7; // @[MemPrimitives.scala 123:41:@49081.4]
  assign _T_5717 = StickySelects_19_io_outs_8; // @[MemPrimitives.scala 123:41:@49082.4]
  assign _T_5718 = StickySelects_19_io_outs_9; // @[MemPrimitives.scala 123:41:@49083.4]
  assign _T_5719 = StickySelects_19_io_outs_10; // @[MemPrimitives.scala 123:41:@49084.4]
  assign _T_5720 = StickySelects_19_io_outs_11; // @[MemPrimitives.scala 123:41:@49085.4]
  assign _T_5721 = StickySelects_19_io_outs_12; // @[MemPrimitives.scala 123:41:@49086.4]
  assign _T_5722 = StickySelects_19_io_outs_13; // @[MemPrimitives.scala 123:41:@49087.4]
  assign _T_5723 = StickySelects_19_io_outs_14; // @[MemPrimitives.scala 123:41:@49088.4]
  assign _T_5725 = {_T_5709,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@49090.4]
  assign _T_5727 = {_T_5710,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@49092.4]
  assign _T_5729 = {_T_5711,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@49094.4]
  assign _T_5731 = {_T_5712,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@49096.4]
  assign _T_5733 = {_T_5713,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@49098.4]
  assign _T_5735 = {_T_5714,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@49100.4]
  assign _T_5737 = {_T_5715,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@49102.4]
  assign _T_5739 = {_T_5716,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@49104.4]
  assign _T_5741 = {_T_5717,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@49106.4]
  assign _T_5743 = {_T_5718,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@49108.4]
  assign _T_5745 = {_T_5719,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@49110.4]
  assign _T_5747 = {_T_5720,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@49112.4]
  assign _T_5749 = {_T_5721,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@49114.4]
  assign _T_5751 = {_T_5722,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@49116.4]
  assign _T_5753 = {_T_5723,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@49118.4]
  assign _T_5754 = _T_5722 ? _T_5751 : _T_5753; // @[Mux.scala 31:69:@49119.4]
  assign _T_5755 = _T_5721 ? _T_5749 : _T_5754; // @[Mux.scala 31:69:@49120.4]
  assign _T_5756 = _T_5720 ? _T_5747 : _T_5755; // @[Mux.scala 31:69:@49121.4]
  assign _T_5757 = _T_5719 ? _T_5745 : _T_5756; // @[Mux.scala 31:69:@49122.4]
  assign _T_5758 = _T_5718 ? _T_5743 : _T_5757; // @[Mux.scala 31:69:@49123.4]
  assign _T_5759 = _T_5717 ? _T_5741 : _T_5758; // @[Mux.scala 31:69:@49124.4]
  assign _T_5760 = _T_5716 ? _T_5739 : _T_5759; // @[Mux.scala 31:69:@49125.4]
  assign _T_5761 = _T_5715 ? _T_5737 : _T_5760; // @[Mux.scala 31:69:@49126.4]
  assign _T_5762 = _T_5714 ? _T_5735 : _T_5761; // @[Mux.scala 31:69:@49127.4]
  assign _T_5763 = _T_5713 ? _T_5733 : _T_5762; // @[Mux.scala 31:69:@49128.4]
  assign _T_5764 = _T_5712 ? _T_5731 : _T_5763; // @[Mux.scala 31:69:@49129.4]
  assign _T_5765 = _T_5711 ? _T_5729 : _T_5764; // @[Mux.scala 31:69:@49130.4]
  assign _T_5766 = _T_5710 ? _T_5727 : _T_5765; // @[Mux.scala 31:69:@49131.4]
  assign _T_5767 = _T_5709 ? _T_5725 : _T_5766; // @[Mux.scala 31:69:@49132.4]
  assign _T_5772 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49139.4]
  assign _T_5775 = _T_5772 & _T_2734; // @[MemPrimitives.scala 110:228:@49141.4]
  assign _T_5778 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49143.4]
  assign _T_5781 = _T_5778 & _T_2740; // @[MemPrimitives.scala 110:228:@49145.4]
  assign _T_5784 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49147.4]
  assign _T_5787 = _T_5784 & _T_2746; // @[MemPrimitives.scala 110:228:@49149.4]
  assign _T_5790 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49151.4]
  assign _T_5793 = _T_5790 & _T_2752; // @[MemPrimitives.scala 110:228:@49153.4]
  assign _T_5796 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49155.4]
  assign _T_5799 = _T_5796 & _T_2758; // @[MemPrimitives.scala 110:228:@49157.4]
  assign _T_5802 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49159.4]
  assign _T_5805 = _T_5802 & _T_2764; // @[MemPrimitives.scala 110:228:@49161.4]
  assign _T_5808 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49163.4]
  assign _T_5811 = _T_5808 & _T_2770; // @[MemPrimitives.scala 110:228:@49165.4]
  assign _T_5814 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49167.4]
  assign _T_5817 = _T_5814 & _T_2776; // @[MemPrimitives.scala 110:228:@49169.4]
  assign _T_5820 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49171.4]
  assign _T_5823 = _T_5820 & _T_2782; // @[MemPrimitives.scala 110:228:@49173.4]
  assign _T_5826 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49175.4]
  assign _T_5829 = _T_5826 & _T_2788; // @[MemPrimitives.scala 110:228:@49177.4]
  assign _T_5832 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49179.4]
  assign _T_5835 = _T_5832 & _T_2794; // @[MemPrimitives.scala 110:228:@49181.4]
  assign _T_5838 = io_rPort_19_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49183.4]
  assign _T_5841 = _T_5838 & _T_2800; // @[MemPrimitives.scala 110:228:@49185.4]
  assign _T_5844 = io_rPort_22_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49187.4]
  assign _T_5847 = _T_5844 & _T_2806; // @[MemPrimitives.scala 110:228:@49189.4]
  assign _T_5850 = io_rPort_26_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49191.4]
  assign _T_5853 = _T_5850 & _T_2812; // @[MemPrimitives.scala 110:228:@49193.4]
  assign _T_5856 = io_rPort_29_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49195.4]
  assign _T_5859 = _T_5856 & _T_2818; // @[MemPrimitives.scala 110:228:@49197.4]
  assign _T_5861 = StickySelects_20_io_outs_0; // @[MemPrimitives.scala 123:41:@49217.4]
  assign _T_5862 = StickySelects_20_io_outs_1; // @[MemPrimitives.scala 123:41:@49218.4]
  assign _T_5863 = StickySelects_20_io_outs_2; // @[MemPrimitives.scala 123:41:@49219.4]
  assign _T_5864 = StickySelects_20_io_outs_3; // @[MemPrimitives.scala 123:41:@49220.4]
  assign _T_5865 = StickySelects_20_io_outs_4; // @[MemPrimitives.scala 123:41:@49221.4]
  assign _T_5866 = StickySelects_20_io_outs_5; // @[MemPrimitives.scala 123:41:@49222.4]
  assign _T_5867 = StickySelects_20_io_outs_6; // @[MemPrimitives.scala 123:41:@49223.4]
  assign _T_5868 = StickySelects_20_io_outs_7; // @[MemPrimitives.scala 123:41:@49224.4]
  assign _T_5869 = StickySelects_20_io_outs_8; // @[MemPrimitives.scala 123:41:@49225.4]
  assign _T_5870 = StickySelects_20_io_outs_9; // @[MemPrimitives.scala 123:41:@49226.4]
  assign _T_5871 = StickySelects_20_io_outs_10; // @[MemPrimitives.scala 123:41:@49227.4]
  assign _T_5872 = StickySelects_20_io_outs_11; // @[MemPrimitives.scala 123:41:@49228.4]
  assign _T_5873 = StickySelects_20_io_outs_12; // @[MemPrimitives.scala 123:41:@49229.4]
  assign _T_5874 = StickySelects_20_io_outs_13; // @[MemPrimitives.scala 123:41:@49230.4]
  assign _T_5875 = StickySelects_20_io_outs_14; // @[MemPrimitives.scala 123:41:@49231.4]
  assign _T_5877 = {_T_5861,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@49233.4]
  assign _T_5879 = {_T_5862,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@49235.4]
  assign _T_5881 = {_T_5863,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@49237.4]
  assign _T_5883 = {_T_5864,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@49239.4]
  assign _T_5885 = {_T_5865,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@49241.4]
  assign _T_5887 = {_T_5866,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@49243.4]
  assign _T_5889 = {_T_5867,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@49245.4]
  assign _T_5891 = {_T_5868,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@49247.4]
  assign _T_5893 = {_T_5869,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@49249.4]
  assign _T_5895 = {_T_5870,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@49251.4]
  assign _T_5897 = {_T_5871,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@49253.4]
  assign _T_5899 = {_T_5872,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@49255.4]
  assign _T_5901 = {_T_5873,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@49257.4]
  assign _T_5903 = {_T_5874,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@49259.4]
  assign _T_5905 = {_T_5875,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@49261.4]
  assign _T_5906 = _T_5874 ? _T_5903 : _T_5905; // @[Mux.scala 31:69:@49262.4]
  assign _T_5907 = _T_5873 ? _T_5901 : _T_5906; // @[Mux.scala 31:69:@49263.4]
  assign _T_5908 = _T_5872 ? _T_5899 : _T_5907; // @[Mux.scala 31:69:@49264.4]
  assign _T_5909 = _T_5871 ? _T_5897 : _T_5908; // @[Mux.scala 31:69:@49265.4]
  assign _T_5910 = _T_5870 ? _T_5895 : _T_5909; // @[Mux.scala 31:69:@49266.4]
  assign _T_5911 = _T_5869 ? _T_5893 : _T_5910; // @[Mux.scala 31:69:@49267.4]
  assign _T_5912 = _T_5868 ? _T_5891 : _T_5911; // @[Mux.scala 31:69:@49268.4]
  assign _T_5913 = _T_5867 ? _T_5889 : _T_5912; // @[Mux.scala 31:69:@49269.4]
  assign _T_5914 = _T_5866 ? _T_5887 : _T_5913; // @[Mux.scala 31:69:@49270.4]
  assign _T_5915 = _T_5865 ? _T_5885 : _T_5914; // @[Mux.scala 31:69:@49271.4]
  assign _T_5916 = _T_5864 ? _T_5883 : _T_5915; // @[Mux.scala 31:69:@49272.4]
  assign _T_5917 = _T_5863 ? _T_5881 : _T_5916; // @[Mux.scala 31:69:@49273.4]
  assign _T_5918 = _T_5862 ? _T_5879 : _T_5917; // @[Mux.scala 31:69:@49274.4]
  assign _T_5919 = _T_5861 ? _T_5877 : _T_5918; // @[Mux.scala 31:69:@49275.4]
  assign _T_5924 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49282.4]
  assign _T_5927 = _T_5924 & _T_2886; // @[MemPrimitives.scala 110:228:@49284.4]
  assign _T_5930 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49286.4]
  assign _T_5933 = _T_5930 & _T_2892; // @[MemPrimitives.scala 110:228:@49288.4]
  assign _T_5936 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49290.4]
  assign _T_5939 = _T_5936 & _T_2898; // @[MemPrimitives.scala 110:228:@49292.4]
  assign _T_5942 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49294.4]
  assign _T_5945 = _T_5942 & _T_2904; // @[MemPrimitives.scala 110:228:@49296.4]
  assign _T_5948 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49298.4]
  assign _T_5951 = _T_5948 & _T_2910; // @[MemPrimitives.scala 110:228:@49300.4]
  assign _T_5954 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49302.4]
  assign _T_5957 = _T_5954 & _T_2916; // @[MemPrimitives.scala 110:228:@49304.4]
  assign _T_5960 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49306.4]
  assign _T_5963 = _T_5960 & _T_2922; // @[MemPrimitives.scala 110:228:@49308.4]
  assign _T_5966 = io_rPort_18_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49310.4]
  assign _T_5969 = _T_5966 & _T_2928; // @[MemPrimitives.scala 110:228:@49312.4]
  assign _T_5972 = io_rPort_20_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49314.4]
  assign _T_5975 = _T_5972 & _T_2934; // @[MemPrimitives.scala 110:228:@49316.4]
  assign _T_5978 = io_rPort_21_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49318.4]
  assign _T_5981 = _T_5978 & _T_2940; // @[MemPrimitives.scala 110:228:@49320.4]
  assign _T_5984 = io_rPort_23_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49322.4]
  assign _T_5987 = _T_5984 & _T_2946; // @[MemPrimitives.scala 110:228:@49324.4]
  assign _T_5990 = io_rPort_24_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49326.4]
  assign _T_5993 = _T_5990 & _T_2952; // @[MemPrimitives.scala 110:228:@49328.4]
  assign _T_5996 = io_rPort_25_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49330.4]
  assign _T_5999 = _T_5996 & _T_2958; // @[MemPrimitives.scala 110:228:@49332.4]
  assign _T_6002 = io_rPort_27_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49334.4]
  assign _T_6005 = _T_6002 & _T_2964; // @[MemPrimitives.scala 110:228:@49336.4]
  assign _T_6008 = io_rPort_28_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@49338.4]
  assign _T_6011 = _T_6008 & _T_2970; // @[MemPrimitives.scala 110:228:@49340.4]
  assign _T_6013 = StickySelects_21_io_outs_0; // @[MemPrimitives.scala 123:41:@49360.4]
  assign _T_6014 = StickySelects_21_io_outs_1; // @[MemPrimitives.scala 123:41:@49361.4]
  assign _T_6015 = StickySelects_21_io_outs_2; // @[MemPrimitives.scala 123:41:@49362.4]
  assign _T_6016 = StickySelects_21_io_outs_3; // @[MemPrimitives.scala 123:41:@49363.4]
  assign _T_6017 = StickySelects_21_io_outs_4; // @[MemPrimitives.scala 123:41:@49364.4]
  assign _T_6018 = StickySelects_21_io_outs_5; // @[MemPrimitives.scala 123:41:@49365.4]
  assign _T_6019 = StickySelects_21_io_outs_6; // @[MemPrimitives.scala 123:41:@49366.4]
  assign _T_6020 = StickySelects_21_io_outs_7; // @[MemPrimitives.scala 123:41:@49367.4]
  assign _T_6021 = StickySelects_21_io_outs_8; // @[MemPrimitives.scala 123:41:@49368.4]
  assign _T_6022 = StickySelects_21_io_outs_9; // @[MemPrimitives.scala 123:41:@49369.4]
  assign _T_6023 = StickySelects_21_io_outs_10; // @[MemPrimitives.scala 123:41:@49370.4]
  assign _T_6024 = StickySelects_21_io_outs_11; // @[MemPrimitives.scala 123:41:@49371.4]
  assign _T_6025 = StickySelects_21_io_outs_12; // @[MemPrimitives.scala 123:41:@49372.4]
  assign _T_6026 = StickySelects_21_io_outs_13; // @[MemPrimitives.scala 123:41:@49373.4]
  assign _T_6027 = StickySelects_21_io_outs_14; // @[MemPrimitives.scala 123:41:@49374.4]
  assign _T_6029 = {_T_6013,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@49376.4]
  assign _T_6031 = {_T_6014,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@49378.4]
  assign _T_6033 = {_T_6015,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@49380.4]
  assign _T_6035 = {_T_6016,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@49382.4]
  assign _T_6037 = {_T_6017,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@49384.4]
  assign _T_6039 = {_T_6018,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@49386.4]
  assign _T_6041 = {_T_6019,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@49388.4]
  assign _T_6043 = {_T_6020,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@49390.4]
  assign _T_6045 = {_T_6021,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@49392.4]
  assign _T_6047 = {_T_6022,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@49394.4]
  assign _T_6049 = {_T_6023,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@49396.4]
  assign _T_6051 = {_T_6024,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@49398.4]
  assign _T_6053 = {_T_6025,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@49400.4]
  assign _T_6055 = {_T_6026,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@49402.4]
  assign _T_6057 = {_T_6027,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@49404.4]
  assign _T_6058 = _T_6026 ? _T_6055 : _T_6057; // @[Mux.scala 31:69:@49405.4]
  assign _T_6059 = _T_6025 ? _T_6053 : _T_6058; // @[Mux.scala 31:69:@49406.4]
  assign _T_6060 = _T_6024 ? _T_6051 : _T_6059; // @[Mux.scala 31:69:@49407.4]
  assign _T_6061 = _T_6023 ? _T_6049 : _T_6060; // @[Mux.scala 31:69:@49408.4]
  assign _T_6062 = _T_6022 ? _T_6047 : _T_6061; // @[Mux.scala 31:69:@49409.4]
  assign _T_6063 = _T_6021 ? _T_6045 : _T_6062; // @[Mux.scala 31:69:@49410.4]
  assign _T_6064 = _T_6020 ? _T_6043 : _T_6063; // @[Mux.scala 31:69:@49411.4]
  assign _T_6065 = _T_6019 ? _T_6041 : _T_6064; // @[Mux.scala 31:69:@49412.4]
  assign _T_6066 = _T_6018 ? _T_6039 : _T_6065; // @[Mux.scala 31:69:@49413.4]
  assign _T_6067 = _T_6017 ? _T_6037 : _T_6066; // @[Mux.scala 31:69:@49414.4]
  assign _T_6068 = _T_6016 ? _T_6035 : _T_6067; // @[Mux.scala 31:69:@49415.4]
  assign _T_6069 = _T_6015 ? _T_6033 : _T_6068; // @[Mux.scala 31:69:@49416.4]
  assign _T_6070 = _T_6014 ? _T_6031 : _T_6069; // @[Mux.scala 31:69:@49417.4]
  assign _T_6071 = _T_6013 ? _T_6029 : _T_6070; // @[Mux.scala 31:69:@49418.4]
  assign _T_6079 = _T_5772 & _T_3038; // @[MemPrimitives.scala 110:228:@49427.4]
  assign _T_6085 = _T_5778 & _T_3044; // @[MemPrimitives.scala 110:228:@49431.4]
  assign _T_6091 = _T_5784 & _T_3050; // @[MemPrimitives.scala 110:228:@49435.4]
  assign _T_6097 = _T_5790 & _T_3056; // @[MemPrimitives.scala 110:228:@49439.4]
  assign _T_6103 = _T_5796 & _T_3062; // @[MemPrimitives.scala 110:228:@49443.4]
  assign _T_6109 = _T_5802 & _T_3068; // @[MemPrimitives.scala 110:228:@49447.4]
  assign _T_6115 = _T_5808 & _T_3074; // @[MemPrimitives.scala 110:228:@49451.4]
  assign _T_6121 = _T_5814 & _T_3080; // @[MemPrimitives.scala 110:228:@49455.4]
  assign _T_6127 = _T_5820 & _T_3086; // @[MemPrimitives.scala 110:228:@49459.4]
  assign _T_6133 = _T_5826 & _T_3092; // @[MemPrimitives.scala 110:228:@49463.4]
  assign _T_6139 = _T_5832 & _T_3098; // @[MemPrimitives.scala 110:228:@49467.4]
  assign _T_6145 = _T_5838 & _T_3104; // @[MemPrimitives.scala 110:228:@49471.4]
  assign _T_6151 = _T_5844 & _T_3110; // @[MemPrimitives.scala 110:228:@49475.4]
  assign _T_6157 = _T_5850 & _T_3116; // @[MemPrimitives.scala 110:228:@49479.4]
  assign _T_6163 = _T_5856 & _T_3122; // @[MemPrimitives.scala 110:228:@49483.4]
  assign _T_6165 = StickySelects_22_io_outs_0; // @[MemPrimitives.scala 123:41:@49503.4]
  assign _T_6166 = StickySelects_22_io_outs_1; // @[MemPrimitives.scala 123:41:@49504.4]
  assign _T_6167 = StickySelects_22_io_outs_2; // @[MemPrimitives.scala 123:41:@49505.4]
  assign _T_6168 = StickySelects_22_io_outs_3; // @[MemPrimitives.scala 123:41:@49506.4]
  assign _T_6169 = StickySelects_22_io_outs_4; // @[MemPrimitives.scala 123:41:@49507.4]
  assign _T_6170 = StickySelects_22_io_outs_5; // @[MemPrimitives.scala 123:41:@49508.4]
  assign _T_6171 = StickySelects_22_io_outs_6; // @[MemPrimitives.scala 123:41:@49509.4]
  assign _T_6172 = StickySelects_22_io_outs_7; // @[MemPrimitives.scala 123:41:@49510.4]
  assign _T_6173 = StickySelects_22_io_outs_8; // @[MemPrimitives.scala 123:41:@49511.4]
  assign _T_6174 = StickySelects_22_io_outs_9; // @[MemPrimitives.scala 123:41:@49512.4]
  assign _T_6175 = StickySelects_22_io_outs_10; // @[MemPrimitives.scala 123:41:@49513.4]
  assign _T_6176 = StickySelects_22_io_outs_11; // @[MemPrimitives.scala 123:41:@49514.4]
  assign _T_6177 = StickySelects_22_io_outs_12; // @[MemPrimitives.scala 123:41:@49515.4]
  assign _T_6178 = StickySelects_22_io_outs_13; // @[MemPrimitives.scala 123:41:@49516.4]
  assign _T_6179 = StickySelects_22_io_outs_14; // @[MemPrimitives.scala 123:41:@49517.4]
  assign _T_6181 = {_T_6165,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@49519.4]
  assign _T_6183 = {_T_6166,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@49521.4]
  assign _T_6185 = {_T_6167,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@49523.4]
  assign _T_6187 = {_T_6168,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@49525.4]
  assign _T_6189 = {_T_6169,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@49527.4]
  assign _T_6191 = {_T_6170,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@49529.4]
  assign _T_6193 = {_T_6171,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@49531.4]
  assign _T_6195 = {_T_6172,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@49533.4]
  assign _T_6197 = {_T_6173,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@49535.4]
  assign _T_6199 = {_T_6174,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@49537.4]
  assign _T_6201 = {_T_6175,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@49539.4]
  assign _T_6203 = {_T_6176,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@49541.4]
  assign _T_6205 = {_T_6177,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@49543.4]
  assign _T_6207 = {_T_6178,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@49545.4]
  assign _T_6209 = {_T_6179,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@49547.4]
  assign _T_6210 = _T_6178 ? _T_6207 : _T_6209; // @[Mux.scala 31:69:@49548.4]
  assign _T_6211 = _T_6177 ? _T_6205 : _T_6210; // @[Mux.scala 31:69:@49549.4]
  assign _T_6212 = _T_6176 ? _T_6203 : _T_6211; // @[Mux.scala 31:69:@49550.4]
  assign _T_6213 = _T_6175 ? _T_6201 : _T_6212; // @[Mux.scala 31:69:@49551.4]
  assign _T_6214 = _T_6174 ? _T_6199 : _T_6213; // @[Mux.scala 31:69:@49552.4]
  assign _T_6215 = _T_6173 ? _T_6197 : _T_6214; // @[Mux.scala 31:69:@49553.4]
  assign _T_6216 = _T_6172 ? _T_6195 : _T_6215; // @[Mux.scala 31:69:@49554.4]
  assign _T_6217 = _T_6171 ? _T_6193 : _T_6216; // @[Mux.scala 31:69:@49555.4]
  assign _T_6218 = _T_6170 ? _T_6191 : _T_6217; // @[Mux.scala 31:69:@49556.4]
  assign _T_6219 = _T_6169 ? _T_6189 : _T_6218; // @[Mux.scala 31:69:@49557.4]
  assign _T_6220 = _T_6168 ? _T_6187 : _T_6219; // @[Mux.scala 31:69:@49558.4]
  assign _T_6221 = _T_6167 ? _T_6185 : _T_6220; // @[Mux.scala 31:69:@49559.4]
  assign _T_6222 = _T_6166 ? _T_6183 : _T_6221; // @[Mux.scala 31:69:@49560.4]
  assign _T_6223 = _T_6165 ? _T_6181 : _T_6222; // @[Mux.scala 31:69:@49561.4]
  assign _T_6231 = _T_5924 & _T_3190; // @[MemPrimitives.scala 110:228:@49570.4]
  assign _T_6237 = _T_5930 & _T_3196; // @[MemPrimitives.scala 110:228:@49574.4]
  assign _T_6243 = _T_5936 & _T_3202; // @[MemPrimitives.scala 110:228:@49578.4]
  assign _T_6249 = _T_5942 & _T_3208; // @[MemPrimitives.scala 110:228:@49582.4]
  assign _T_6255 = _T_5948 & _T_3214; // @[MemPrimitives.scala 110:228:@49586.4]
  assign _T_6261 = _T_5954 & _T_3220; // @[MemPrimitives.scala 110:228:@49590.4]
  assign _T_6267 = _T_5960 & _T_3226; // @[MemPrimitives.scala 110:228:@49594.4]
  assign _T_6273 = _T_5966 & _T_3232; // @[MemPrimitives.scala 110:228:@49598.4]
  assign _T_6279 = _T_5972 & _T_3238; // @[MemPrimitives.scala 110:228:@49602.4]
  assign _T_6285 = _T_5978 & _T_3244; // @[MemPrimitives.scala 110:228:@49606.4]
  assign _T_6291 = _T_5984 & _T_3250; // @[MemPrimitives.scala 110:228:@49610.4]
  assign _T_6297 = _T_5990 & _T_3256; // @[MemPrimitives.scala 110:228:@49614.4]
  assign _T_6303 = _T_5996 & _T_3262; // @[MemPrimitives.scala 110:228:@49618.4]
  assign _T_6309 = _T_6002 & _T_3268; // @[MemPrimitives.scala 110:228:@49622.4]
  assign _T_6315 = _T_6008 & _T_3274; // @[MemPrimitives.scala 110:228:@49626.4]
  assign _T_6317 = StickySelects_23_io_outs_0; // @[MemPrimitives.scala 123:41:@49646.4]
  assign _T_6318 = StickySelects_23_io_outs_1; // @[MemPrimitives.scala 123:41:@49647.4]
  assign _T_6319 = StickySelects_23_io_outs_2; // @[MemPrimitives.scala 123:41:@49648.4]
  assign _T_6320 = StickySelects_23_io_outs_3; // @[MemPrimitives.scala 123:41:@49649.4]
  assign _T_6321 = StickySelects_23_io_outs_4; // @[MemPrimitives.scala 123:41:@49650.4]
  assign _T_6322 = StickySelects_23_io_outs_5; // @[MemPrimitives.scala 123:41:@49651.4]
  assign _T_6323 = StickySelects_23_io_outs_6; // @[MemPrimitives.scala 123:41:@49652.4]
  assign _T_6324 = StickySelects_23_io_outs_7; // @[MemPrimitives.scala 123:41:@49653.4]
  assign _T_6325 = StickySelects_23_io_outs_8; // @[MemPrimitives.scala 123:41:@49654.4]
  assign _T_6326 = StickySelects_23_io_outs_9; // @[MemPrimitives.scala 123:41:@49655.4]
  assign _T_6327 = StickySelects_23_io_outs_10; // @[MemPrimitives.scala 123:41:@49656.4]
  assign _T_6328 = StickySelects_23_io_outs_11; // @[MemPrimitives.scala 123:41:@49657.4]
  assign _T_6329 = StickySelects_23_io_outs_12; // @[MemPrimitives.scala 123:41:@49658.4]
  assign _T_6330 = StickySelects_23_io_outs_13; // @[MemPrimitives.scala 123:41:@49659.4]
  assign _T_6331 = StickySelects_23_io_outs_14; // @[MemPrimitives.scala 123:41:@49660.4]
  assign _T_6333 = {_T_6317,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@49662.4]
  assign _T_6335 = {_T_6318,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@49664.4]
  assign _T_6337 = {_T_6319,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@49666.4]
  assign _T_6339 = {_T_6320,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@49668.4]
  assign _T_6341 = {_T_6321,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@49670.4]
  assign _T_6343 = {_T_6322,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@49672.4]
  assign _T_6345 = {_T_6323,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@49674.4]
  assign _T_6347 = {_T_6324,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@49676.4]
  assign _T_6349 = {_T_6325,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@49678.4]
  assign _T_6351 = {_T_6326,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@49680.4]
  assign _T_6353 = {_T_6327,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@49682.4]
  assign _T_6355 = {_T_6328,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@49684.4]
  assign _T_6357 = {_T_6329,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@49686.4]
  assign _T_6359 = {_T_6330,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@49688.4]
  assign _T_6361 = {_T_6331,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@49690.4]
  assign _T_6362 = _T_6330 ? _T_6359 : _T_6361; // @[Mux.scala 31:69:@49691.4]
  assign _T_6363 = _T_6329 ? _T_6357 : _T_6362; // @[Mux.scala 31:69:@49692.4]
  assign _T_6364 = _T_6328 ? _T_6355 : _T_6363; // @[Mux.scala 31:69:@49693.4]
  assign _T_6365 = _T_6327 ? _T_6353 : _T_6364; // @[Mux.scala 31:69:@49694.4]
  assign _T_6366 = _T_6326 ? _T_6351 : _T_6365; // @[Mux.scala 31:69:@49695.4]
  assign _T_6367 = _T_6325 ? _T_6349 : _T_6366; // @[Mux.scala 31:69:@49696.4]
  assign _T_6368 = _T_6324 ? _T_6347 : _T_6367; // @[Mux.scala 31:69:@49697.4]
  assign _T_6369 = _T_6323 ? _T_6345 : _T_6368; // @[Mux.scala 31:69:@49698.4]
  assign _T_6370 = _T_6322 ? _T_6343 : _T_6369; // @[Mux.scala 31:69:@49699.4]
  assign _T_6371 = _T_6321 ? _T_6341 : _T_6370; // @[Mux.scala 31:69:@49700.4]
  assign _T_6372 = _T_6320 ? _T_6339 : _T_6371; // @[Mux.scala 31:69:@49701.4]
  assign _T_6373 = _T_6319 ? _T_6337 : _T_6372; // @[Mux.scala 31:69:@49702.4]
  assign _T_6374 = _T_6318 ? _T_6335 : _T_6373; // @[Mux.scala 31:69:@49703.4]
  assign _T_6375 = _T_6317 ? _T_6333 : _T_6374; // @[Mux.scala 31:69:@49704.4]
  assign _T_6383 = _T_5772 & _T_3342; // @[MemPrimitives.scala 110:228:@49713.4]
  assign _T_6389 = _T_5778 & _T_3348; // @[MemPrimitives.scala 110:228:@49717.4]
  assign _T_6395 = _T_5784 & _T_3354; // @[MemPrimitives.scala 110:228:@49721.4]
  assign _T_6401 = _T_5790 & _T_3360; // @[MemPrimitives.scala 110:228:@49725.4]
  assign _T_6407 = _T_5796 & _T_3366; // @[MemPrimitives.scala 110:228:@49729.4]
  assign _T_6413 = _T_5802 & _T_3372; // @[MemPrimitives.scala 110:228:@49733.4]
  assign _T_6419 = _T_5808 & _T_3378; // @[MemPrimitives.scala 110:228:@49737.4]
  assign _T_6425 = _T_5814 & _T_3384; // @[MemPrimitives.scala 110:228:@49741.4]
  assign _T_6431 = _T_5820 & _T_3390; // @[MemPrimitives.scala 110:228:@49745.4]
  assign _T_6437 = _T_5826 & _T_3396; // @[MemPrimitives.scala 110:228:@49749.4]
  assign _T_6443 = _T_5832 & _T_3402; // @[MemPrimitives.scala 110:228:@49753.4]
  assign _T_6449 = _T_5838 & _T_3408; // @[MemPrimitives.scala 110:228:@49757.4]
  assign _T_6455 = _T_5844 & _T_3414; // @[MemPrimitives.scala 110:228:@49761.4]
  assign _T_6461 = _T_5850 & _T_3420; // @[MemPrimitives.scala 110:228:@49765.4]
  assign _T_6467 = _T_5856 & _T_3426; // @[MemPrimitives.scala 110:228:@49769.4]
  assign _T_6469 = StickySelects_24_io_outs_0; // @[MemPrimitives.scala 123:41:@49789.4]
  assign _T_6470 = StickySelects_24_io_outs_1; // @[MemPrimitives.scala 123:41:@49790.4]
  assign _T_6471 = StickySelects_24_io_outs_2; // @[MemPrimitives.scala 123:41:@49791.4]
  assign _T_6472 = StickySelects_24_io_outs_3; // @[MemPrimitives.scala 123:41:@49792.4]
  assign _T_6473 = StickySelects_24_io_outs_4; // @[MemPrimitives.scala 123:41:@49793.4]
  assign _T_6474 = StickySelects_24_io_outs_5; // @[MemPrimitives.scala 123:41:@49794.4]
  assign _T_6475 = StickySelects_24_io_outs_6; // @[MemPrimitives.scala 123:41:@49795.4]
  assign _T_6476 = StickySelects_24_io_outs_7; // @[MemPrimitives.scala 123:41:@49796.4]
  assign _T_6477 = StickySelects_24_io_outs_8; // @[MemPrimitives.scala 123:41:@49797.4]
  assign _T_6478 = StickySelects_24_io_outs_9; // @[MemPrimitives.scala 123:41:@49798.4]
  assign _T_6479 = StickySelects_24_io_outs_10; // @[MemPrimitives.scala 123:41:@49799.4]
  assign _T_6480 = StickySelects_24_io_outs_11; // @[MemPrimitives.scala 123:41:@49800.4]
  assign _T_6481 = StickySelects_24_io_outs_12; // @[MemPrimitives.scala 123:41:@49801.4]
  assign _T_6482 = StickySelects_24_io_outs_13; // @[MemPrimitives.scala 123:41:@49802.4]
  assign _T_6483 = StickySelects_24_io_outs_14; // @[MemPrimitives.scala 123:41:@49803.4]
  assign _T_6485 = {_T_6469,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@49805.4]
  assign _T_6487 = {_T_6470,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@49807.4]
  assign _T_6489 = {_T_6471,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@49809.4]
  assign _T_6491 = {_T_6472,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@49811.4]
  assign _T_6493 = {_T_6473,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@49813.4]
  assign _T_6495 = {_T_6474,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@49815.4]
  assign _T_6497 = {_T_6475,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@49817.4]
  assign _T_6499 = {_T_6476,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@49819.4]
  assign _T_6501 = {_T_6477,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@49821.4]
  assign _T_6503 = {_T_6478,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@49823.4]
  assign _T_6505 = {_T_6479,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@49825.4]
  assign _T_6507 = {_T_6480,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@49827.4]
  assign _T_6509 = {_T_6481,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@49829.4]
  assign _T_6511 = {_T_6482,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@49831.4]
  assign _T_6513 = {_T_6483,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@49833.4]
  assign _T_6514 = _T_6482 ? _T_6511 : _T_6513; // @[Mux.scala 31:69:@49834.4]
  assign _T_6515 = _T_6481 ? _T_6509 : _T_6514; // @[Mux.scala 31:69:@49835.4]
  assign _T_6516 = _T_6480 ? _T_6507 : _T_6515; // @[Mux.scala 31:69:@49836.4]
  assign _T_6517 = _T_6479 ? _T_6505 : _T_6516; // @[Mux.scala 31:69:@49837.4]
  assign _T_6518 = _T_6478 ? _T_6503 : _T_6517; // @[Mux.scala 31:69:@49838.4]
  assign _T_6519 = _T_6477 ? _T_6501 : _T_6518; // @[Mux.scala 31:69:@49839.4]
  assign _T_6520 = _T_6476 ? _T_6499 : _T_6519; // @[Mux.scala 31:69:@49840.4]
  assign _T_6521 = _T_6475 ? _T_6497 : _T_6520; // @[Mux.scala 31:69:@49841.4]
  assign _T_6522 = _T_6474 ? _T_6495 : _T_6521; // @[Mux.scala 31:69:@49842.4]
  assign _T_6523 = _T_6473 ? _T_6493 : _T_6522; // @[Mux.scala 31:69:@49843.4]
  assign _T_6524 = _T_6472 ? _T_6491 : _T_6523; // @[Mux.scala 31:69:@49844.4]
  assign _T_6525 = _T_6471 ? _T_6489 : _T_6524; // @[Mux.scala 31:69:@49845.4]
  assign _T_6526 = _T_6470 ? _T_6487 : _T_6525; // @[Mux.scala 31:69:@49846.4]
  assign _T_6527 = _T_6469 ? _T_6485 : _T_6526; // @[Mux.scala 31:69:@49847.4]
  assign _T_6535 = _T_5924 & _T_3494; // @[MemPrimitives.scala 110:228:@49856.4]
  assign _T_6541 = _T_5930 & _T_3500; // @[MemPrimitives.scala 110:228:@49860.4]
  assign _T_6547 = _T_5936 & _T_3506; // @[MemPrimitives.scala 110:228:@49864.4]
  assign _T_6553 = _T_5942 & _T_3512; // @[MemPrimitives.scala 110:228:@49868.4]
  assign _T_6559 = _T_5948 & _T_3518; // @[MemPrimitives.scala 110:228:@49872.4]
  assign _T_6565 = _T_5954 & _T_3524; // @[MemPrimitives.scala 110:228:@49876.4]
  assign _T_6571 = _T_5960 & _T_3530; // @[MemPrimitives.scala 110:228:@49880.4]
  assign _T_6577 = _T_5966 & _T_3536; // @[MemPrimitives.scala 110:228:@49884.4]
  assign _T_6583 = _T_5972 & _T_3542; // @[MemPrimitives.scala 110:228:@49888.4]
  assign _T_6589 = _T_5978 & _T_3548; // @[MemPrimitives.scala 110:228:@49892.4]
  assign _T_6595 = _T_5984 & _T_3554; // @[MemPrimitives.scala 110:228:@49896.4]
  assign _T_6601 = _T_5990 & _T_3560; // @[MemPrimitives.scala 110:228:@49900.4]
  assign _T_6607 = _T_5996 & _T_3566; // @[MemPrimitives.scala 110:228:@49904.4]
  assign _T_6613 = _T_6002 & _T_3572; // @[MemPrimitives.scala 110:228:@49908.4]
  assign _T_6619 = _T_6008 & _T_3578; // @[MemPrimitives.scala 110:228:@49912.4]
  assign _T_6621 = StickySelects_25_io_outs_0; // @[MemPrimitives.scala 123:41:@49932.4]
  assign _T_6622 = StickySelects_25_io_outs_1; // @[MemPrimitives.scala 123:41:@49933.4]
  assign _T_6623 = StickySelects_25_io_outs_2; // @[MemPrimitives.scala 123:41:@49934.4]
  assign _T_6624 = StickySelects_25_io_outs_3; // @[MemPrimitives.scala 123:41:@49935.4]
  assign _T_6625 = StickySelects_25_io_outs_4; // @[MemPrimitives.scala 123:41:@49936.4]
  assign _T_6626 = StickySelects_25_io_outs_5; // @[MemPrimitives.scala 123:41:@49937.4]
  assign _T_6627 = StickySelects_25_io_outs_6; // @[MemPrimitives.scala 123:41:@49938.4]
  assign _T_6628 = StickySelects_25_io_outs_7; // @[MemPrimitives.scala 123:41:@49939.4]
  assign _T_6629 = StickySelects_25_io_outs_8; // @[MemPrimitives.scala 123:41:@49940.4]
  assign _T_6630 = StickySelects_25_io_outs_9; // @[MemPrimitives.scala 123:41:@49941.4]
  assign _T_6631 = StickySelects_25_io_outs_10; // @[MemPrimitives.scala 123:41:@49942.4]
  assign _T_6632 = StickySelects_25_io_outs_11; // @[MemPrimitives.scala 123:41:@49943.4]
  assign _T_6633 = StickySelects_25_io_outs_12; // @[MemPrimitives.scala 123:41:@49944.4]
  assign _T_6634 = StickySelects_25_io_outs_13; // @[MemPrimitives.scala 123:41:@49945.4]
  assign _T_6635 = StickySelects_25_io_outs_14; // @[MemPrimitives.scala 123:41:@49946.4]
  assign _T_6637 = {_T_6621,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@49948.4]
  assign _T_6639 = {_T_6622,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@49950.4]
  assign _T_6641 = {_T_6623,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@49952.4]
  assign _T_6643 = {_T_6624,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@49954.4]
  assign _T_6645 = {_T_6625,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@49956.4]
  assign _T_6647 = {_T_6626,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@49958.4]
  assign _T_6649 = {_T_6627,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@49960.4]
  assign _T_6651 = {_T_6628,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@49962.4]
  assign _T_6653 = {_T_6629,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@49964.4]
  assign _T_6655 = {_T_6630,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@49966.4]
  assign _T_6657 = {_T_6631,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@49968.4]
  assign _T_6659 = {_T_6632,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@49970.4]
  assign _T_6661 = {_T_6633,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@49972.4]
  assign _T_6663 = {_T_6634,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@49974.4]
  assign _T_6665 = {_T_6635,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@49976.4]
  assign _T_6666 = _T_6634 ? _T_6663 : _T_6665; // @[Mux.scala 31:69:@49977.4]
  assign _T_6667 = _T_6633 ? _T_6661 : _T_6666; // @[Mux.scala 31:69:@49978.4]
  assign _T_6668 = _T_6632 ? _T_6659 : _T_6667; // @[Mux.scala 31:69:@49979.4]
  assign _T_6669 = _T_6631 ? _T_6657 : _T_6668; // @[Mux.scala 31:69:@49980.4]
  assign _T_6670 = _T_6630 ? _T_6655 : _T_6669; // @[Mux.scala 31:69:@49981.4]
  assign _T_6671 = _T_6629 ? _T_6653 : _T_6670; // @[Mux.scala 31:69:@49982.4]
  assign _T_6672 = _T_6628 ? _T_6651 : _T_6671; // @[Mux.scala 31:69:@49983.4]
  assign _T_6673 = _T_6627 ? _T_6649 : _T_6672; // @[Mux.scala 31:69:@49984.4]
  assign _T_6674 = _T_6626 ? _T_6647 : _T_6673; // @[Mux.scala 31:69:@49985.4]
  assign _T_6675 = _T_6625 ? _T_6645 : _T_6674; // @[Mux.scala 31:69:@49986.4]
  assign _T_6676 = _T_6624 ? _T_6643 : _T_6675; // @[Mux.scala 31:69:@49987.4]
  assign _T_6677 = _T_6623 ? _T_6641 : _T_6676; // @[Mux.scala 31:69:@49988.4]
  assign _T_6678 = _T_6622 ? _T_6639 : _T_6677; // @[Mux.scala 31:69:@49989.4]
  assign _T_6679 = _T_6621 ? _T_6637 : _T_6678; // @[Mux.scala 31:69:@49990.4]
  assign _T_6687 = _T_5772 & _T_3646; // @[MemPrimitives.scala 110:228:@49999.4]
  assign _T_6693 = _T_5778 & _T_3652; // @[MemPrimitives.scala 110:228:@50003.4]
  assign _T_6699 = _T_5784 & _T_3658; // @[MemPrimitives.scala 110:228:@50007.4]
  assign _T_6705 = _T_5790 & _T_3664; // @[MemPrimitives.scala 110:228:@50011.4]
  assign _T_6711 = _T_5796 & _T_3670; // @[MemPrimitives.scala 110:228:@50015.4]
  assign _T_6717 = _T_5802 & _T_3676; // @[MemPrimitives.scala 110:228:@50019.4]
  assign _T_6723 = _T_5808 & _T_3682; // @[MemPrimitives.scala 110:228:@50023.4]
  assign _T_6729 = _T_5814 & _T_3688; // @[MemPrimitives.scala 110:228:@50027.4]
  assign _T_6735 = _T_5820 & _T_3694; // @[MemPrimitives.scala 110:228:@50031.4]
  assign _T_6741 = _T_5826 & _T_3700; // @[MemPrimitives.scala 110:228:@50035.4]
  assign _T_6747 = _T_5832 & _T_3706; // @[MemPrimitives.scala 110:228:@50039.4]
  assign _T_6753 = _T_5838 & _T_3712; // @[MemPrimitives.scala 110:228:@50043.4]
  assign _T_6759 = _T_5844 & _T_3718; // @[MemPrimitives.scala 110:228:@50047.4]
  assign _T_6765 = _T_5850 & _T_3724; // @[MemPrimitives.scala 110:228:@50051.4]
  assign _T_6771 = _T_5856 & _T_3730; // @[MemPrimitives.scala 110:228:@50055.4]
  assign _T_6773 = StickySelects_26_io_outs_0; // @[MemPrimitives.scala 123:41:@50075.4]
  assign _T_6774 = StickySelects_26_io_outs_1; // @[MemPrimitives.scala 123:41:@50076.4]
  assign _T_6775 = StickySelects_26_io_outs_2; // @[MemPrimitives.scala 123:41:@50077.4]
  assign _T_6776 = StickySelects_26_io_outs_3; // @[MemPrimitives.scala 123:41:@50078.4]
  assign _T_6777 = StickySelects_26_io_outs_4; // @[MemPrimitives.scala 123:41:@50079.4]
  assign _T_6778 = StickySelects_26_io_outs_5; // @[MemPrimitives.scala 123:41:@50080.4]
  assign _T_6779 = StickySelects_26_io_outs_6; // @[MemPrimitives.scala 123:41:@50081.4]
  assign _T_6780 = StickySelects_26_io_outs_7; // @[MemPrimitives.scala 123:41:@50082.4]
  assign _T_6781 = StickySelects_26_io_outs_8; // @[MemPrimitives.scala 123:41:@50083.4]
  assign _T_6782 = StickySelects_26_io_outs_9; // @[MemPrimitives.scala 123:41:@50084.4]
  assign _T_6783 = StickySelects_26_io_outs_10; // @[MemPrimitives.scala 123:41:@50085.4]
  assign _T_6784 = StickySelects_26_io_outs_11; // @[MemPrimitives.scala 123:41:@50086.4]
  assign _T_6785 = StickySelects_26_io_outs_12; // @[MemPrimitives.scala 123:41:@50087.4]
  assign _T_6786 = StickySelects_26_io_outs_13; // @[MemPrimitives.scala 123:41:@50088.4]
  assign _T_6787 = StickySelects_26_io_outs_14; // @[MemPrimitives.scala 123:41:@50089.4]
  assign _T_6789 = {_T_6773,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@50091.4]
  assign _T_6791 = {_T_6774,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@50093.4]
  assign _T_6793 = {_T_6775,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@50095.4]
  assign _T_6795 = {_T_6776,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@50097.4]
  assign _T_6797 = {_T_6777,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@50099.4]
  assign _T_6799 = {_T_6778,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@50101.4]
  assign _T_6801 = {_T_6779,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@50103.4]
  assign _T_6803 = {_T_6780,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@50105.4]
  assign _T_6805 = {_T_6781,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@50107.4]
  assign _T_6807 = {_T_6782,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@50109.4]
  assign _T_6809 = {_T_6783,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@50111.4]
  assign _T_6811 = {_T_6784,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@50113.4]
  assign _T_6813 = {_T_6785,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@50115.4]
  assign _T_6815 = {_T_6786,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@50117.4]
  assign _T_6817 = {_T_6787,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@50119.4]
  assign _T_6818 = _T_6786 ? _T_6815 : _T_6817; // @[Mux.scala 31:69:@50120.4]
  assign _T_6819 = _T_6785 ? _T_6813 : _T_6818; // @[Mux.scala 31:69:@50121.4]
  assign _T_6820 = _T_6784 ? _T_6811 : _T_6819; // @[Mux.scala 31:69:@50122.4]
  assign _T_6821 = _T_6783 ? _T_6809 : _T_6820; // @[Mux.scala 31:69:@50123.4]
  assign _T_6822 = _T_6782 ? _T_6807 : _T_6821; // @[Mux.scala 31:69:@50124.4]
  assign _T_6823 = _T_6781 ? _T_6805 : _T_6822; // @[Mux.scala 31:69:@50125.4]
  assign _T_6824 = _T_6780 ? _T_6803 : _T_6823; // @[Mux.scala 31:69:@50126.4]
  assign _T_6825 = _T_6779 ? _T_6801 : _T_6824; // @[Mux.scala 31:69:@50127.4]
  assign _T_6826 = _T_6778 ? _T_6799 : _T_6825; // @[Mux.scala 31:69:@50128.4]
  assign _T_6827 = _T_6777 ? _T_6797 : _T_6826; // @[Mux.scala 31:69:@50129.4]
  assign _T_6828 = _T_6776 ? _T_6795 : _T_6827; // @[Mux.scala 31:69:@50130.4]
  assign _T_6829 = _T_6775 ? _T_6793 : _T_6828; // @[Mux.scala 31:69:@50131.4]
  assign _T_6830 = _T_6774 ? _T_6791 : _T_6829; // @[Mux.scala 31:69:@50132.4]
  assign _T_6831 = _T_6773 ? _T_6789 : _T_6830; // @[Mux.scala 31:69:@50133.4]
  assign _T_6839 = _T_5924 & _T_3798; // @[MemPrimitives.scala 110:228:@50142.4]
  assign _T_6845 = _T_5930 & _T_3804; // @[MemPrimitives.scala 110:228:@50146.4]
  assign _T_6851 = _T_5936 & _T_3810; // @[MemPrimitives.scala 110:228:@50150.4]
  assign _T_6857 = _T_5942 & _T_3816; // @[MemPrimitives.scala 110:228:@50154.4]
  assign _T_6863 = _T_5948 & _T_3822; // @[MemPrimitives.scala 110:228:@50158.4]
  assign _T_6869 = _T_5954 & _T_3828; // @[MemPrimitives.scala 110:228:@50162.4]
  assign _T_6875 = _T_5960 & _T_3834; // @[MemPrimitives.scala 110:228:@50166.4]
  assign _T_6881 = _T_5966 & _T_3840; // @[MemPrimitives.scala 110:228:@50170.4]
  assign _T_6887 = _T_5972 & _T_3846; // @[MemPrimitives.scala 110:228:@50174.4]
  assign _T_6893 = _T_5978 & _T_3852; // @[MemPrimitives.scala 110:228:@50178.4]
  assign _T_6899 = _T_5984 & _T_3858; // @[MemPrimitives.scala 110:228:@50182.4]
  assign _T_6905 = _T_5990 & _T_3864; // @[MemPrimitives.scala 110:228:@50186.4]
  assign _T_6911 = _T_5996 & _T_3870; // @[MemPrimitives.scala 110:228:@50190.4]
  assign _T_6917 = _T_6002 & _T_3876; // @[MemPrimitives.scala 110:228:@50194.4]
  assign _T_6923 = _T_6008 & _T_3882; // @[MemPrimitives.scala 110:228:@50198.4]
  assign _T_6925 = StickySelects_27_io_outs_0; // @[MemPrimitives.scala 123:41:@50218.4]
  assign _T_6926 = StickySelects_27_io_outs_1; // @[MemPrimitives.scala 123:41:@50219.4]
  assign _T_6927 = StickySelects_27_io_outs_2; // @[MemPrimitives.scala 123:41:@50220.4]
  assign _T_6928 = StickySelects_27_io_outs_3; // @[MemPrimitives.scala 123:41:@50221.4]
  assign _T_6929 = StickySelects_27_io_outs_4; // @[MemPrimitives.scala 123:41:@50222.4]
  assign _T_6930 = StickySelects_27_io_outs_5; // @[MemPrimitives.scala 123:41:@50223.4]
  assign _T_6931 = StickySelects_27_io_outs_6; // @[MemPrimitives.scala 123:41:@50224.4]
  assign _T_6932 = StickySelects_27_io_outs_7; // @[MemPrimitives.scala 123:41:@50225.4]
  assign _T_6933 = StickySelects_27_io_outs_8; // @[MemPrimitives.scala 123:41:@50226.4]
  assign _T_6934 = StickySelects_27_io_outs_9; // @[MemPrimitives.scala 123:41:@50227.4]
  assign _T_6935 = StickySelects_27_io_outs_10; // @[MemPrimitives.scala 123:41:@50228.4]
  assign _T_6936 = StickySelects_27_io_outs_11; // @[MemPrimitives.scala 123:41:@50229.4]
  assign _T_6937 = StickySelects_27_io_outs_12; // @[MemPrimitives.scala 123:41:@50230.4]
  assign _T_6938 = StickySelects_27_io_outs_13; // @[MemPrimitives.scala 123:41:@50231.4]
  assign _T_6939 = StickySelects_27_io_outs_14; // @[MemPrimitives.scala 123:41:@50232.4]
  assign _T_6941 = {_T_6925,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@50234.4]
  assign _T_6943 = {_T_6926,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@50236.4]
  assign _T_6945 = {_T_6927,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@50238.4]
  assign _T_6947 = {_T_6928,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@50240.4]
  assign _T_6949 = {_T_6929,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@50242.4]
  assign _T_6951 = {_T_6930,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@50244.4]
  assign _T_6953 = {_T_6931,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@50246.4]
  assign _T_6955 = {_T_6932,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@50248.4]
  assign _T_6957 = {_T_6933,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@50250.4]
  assign _T_6959 = {_T_6934,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@50252.4]
  assign _T_6961 = {_T_6935,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@50254.4]
  assign _T_6963 = {_T_6936,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@50256.4]
  assign _T_6965 = {_T_6937,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@50258.4]
  assign _T_6967 = {_T_6938,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@50260.4]
  assign _T_6969 = {_T_6939,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@50262.4]
  assign _T_6970 = _T_6938 ? _T_6967 : _T_6969; // @[Mux.scala 31:69:@50263.4]
  assign _T_6971 = _T_6937 ? _T_6965 : _T_6970; // @[Mux.scala 31:69:@50264.4]
  assign _T_6972 = _T_6936 ? _T_6963 : _T_6971; // @[Mux.scala 31:69:@50265.4]
  assign _T_6973 = _T_6935 ? _T_6961 : _T_6972; // @[Mux.scala 31:69:@50266.4]
  assign _T_6974 = _T_6934 ? _T_6959 : _T_6973; // @[Mux.scala 31:69:@50267.4]
  assign _T_6975 = _T_6933 ? _T_6957 : _T_6974; // @[Mux.scala 31:69:@50268.4]
  assign _T_6976 = _T_6932 ? _T_6955 : _T_6975; // @[Mux.scala 31:69:@50269.4]
  assign _T_6977 = _T_6931 ? _T_6953 : _T_6976; // @[Mux.scala 31:69:@50270.4]
  assign _T_6978 = _T_6930 ? _T_6951 : _T_6977; // @[Mux.scala 31:69:@50271.4]
  assign _T_6979 = _T_6929 ? _T_6949 : _T_6978; // @[Mux.scala 31:69:@50272.4]
  assign _T_6980 = _T_6928 ? _T_6947 : _T_6979; // @[Mux.scala 31:69:@50273.4]
  assign _T_6981 = _T_6927 ? _T_6945 : _T_6980; // @[Mux.scala 31:69:@50274.4]
  assign _T_6982 = _T_6926 ? _T_6943 : _T_6981; // @[Mux.scala 31:69:@50275.4]
  assign _T_6983 = _T_6925 ? _T_6941 : _T_6982; // @[Mux.scala 31:69:@50276.4]
  assign _T_6991 = _T_5772 & _T_3950; // @[MemPrimitives.scala 110:228:@50285.4]
  assign _T_6997 = _T_5778 & _T_3956; // @[MemPrimitives.scala 110:228:@50289.4]
  assign _T_7003 = _T_5784 & _T_3962; // @[MemPrimitives.scala 110:228:@50293.4]
  assign _T_7009 = _T_5790 & _T_3968; // @[MemPrimitives.scala 110:228:@50297.4]
  assign _T_7015 = _T_5796 & _T_3974; // @[MemPrimitives.scala 110:228:@50301.4]
  assign _T_7021 = _T_5802 & _T_3980; // @[MemPrimitives.scala 110:228:@50305.4]
  assign _T_7027 = _T_5808 & _T_3986; // @[MemPrimitives.scala 110:228:@50309.4]
  assign _T_7033 = _T_5814 & _T_3992; // @[MemPrimitives.scala 110:228:@50313.4]
  assign _T_7039 = _T_5820 & _T_3998; // @[MemPrimitives.scala 110:228:@50317.4]
  assign _T_7045 = _T_5826 & _T_4004; // @[MemPrimitives.scala 110:228:@50321.4]
  assign _T_7051 = _T_5832 & _T_4010; // @[MemPrimitives.scala 110:228:@50325.4]
  assign _T_7057 = _T_5838 & _T_4016; // @[MemPrimitives.scala 110:228:@50329.4]
  assign _T_7063 = _T_5844 & _T_4022; // @[MemPrimitives.scala 110:228:@50333.4]
  assign _T_7069 = _T_5850 & _T_4028; // @[MemPrimitives.scala 110:228:@50337.4]
  assign _T_7075 = _T_5856 & _T_4034; // @[MemPrimitives.scala 110:228:@50341.4]
  assign _T_7077 = StickySelects_28_io_outs_0; // @[MemPrimitives.scala 123:41:@50361.4]
  assign _T_7078 = StickySelects_28_io_outs_1; // @[MemPrimitives.scala 123:41:@50362.4]
  assign _T_7079 = StickySelects_28_io_outs_2; // @[MemPrimitives.scala 123:41:@50363.4]
  assign _T_7080 = StickySelects_28_io_outs_3; // @[MemPrimitives.scala 123:41:@50364.4]
  assign _T_7081 = StickySelects_28_io_outs_4; // @[MemPrimitives.scala 123:41:@50365.4]
  assign _T_7082 = StickySelects_28_io_outs_5; // @[MemPrimitives.scala 123:41:@50366.4]
  assign _T_7083 = StickySelects_28_io_outs_6; // @[MemPrimitives.scala 123:41:@50367.4]
  assign _T_7084 = StickySelects_28_io_outs_7; // @[MemPrimitives.scala 123:41:@50368.4]
  assign _T_7085 = StickySelects_28_io_outs_8; // @[MemPrimitives.scala 123:41:@50369.4]
  assign _T_7086 = StickySelects_28_io_outs_9; // @[MemPrimitives.scala 123:41:@50370.4]
  assign _T_7087 = StickySelects_28_io_outs_10; // @[MemPrimitives.scala 123:41:@50371.4]
  assign _T_7088 = StickySelects_28_io_outs_11; // @[MemPrimitives.scala 123:41:@50372.4]
  assign _T_7089 = StickySelects_28_io_outs_12; // @[MemPrimitives.scala 123:41:@50373.4]
  assign _T_7090 = StickySelects_28_io_outs_13; // @[MemPrimitives.scala 123:41:@50374.4]
  assign _T_7091 = StickySelects_28_io_outs_14; // @[MemPrimitives.scala 123:41:@50375.4]
  assign _T_7093 = {_T_7077,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@50377.4]
  assign _T_7095 = {_T_7078,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@50379.4]
  assign _T_7097 = {_T_7079,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@50381.4]
  assign _T_7099 = {_T_7080,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@50383.4]
  assign _T_7101 = {_T_7081,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@50385.4]
  assign _T_7103 = {_T_7082,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@50387.4]
  assign _T_7105 = {_T_7083,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@50389.4]
  assign _T_7107 = {_T_7084,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@50391.4]
  assign _T_7109 = {_T_7085,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@50393.4]
  assign _T_7111 = {_T_7086,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@50395.4]
  assign _T_7113 = {_T_7087,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@50397.4]
  assign _T_7115 = {_T_7088,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@50399.4]
  assign _T_7117 = {_T_7089,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@50401.4]
  assign _T_7119 = {_T_7090,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@50403.4]
  assign _T_7121 = {_T_7091,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@50405.4]
  assign _T_7122 = _T_7090 ? _T_7119 : _T_7121; // @[Mux.scala 31:69:@50406.4]
  assign _T_7123 = _T_7089 ? _T_7117 : _T_7122; // @[Mux.scala 31:69:@50407.4]
  assign _T_7124 = _T_7088 ? _T_7115 : _T_7123; // @[Mux.scala 31:69:@50408.4]
  assign _T_7125 = _T_7087 ? _T_7113 : _T_7124; // @[Mux.scala 31:69:@50409.4]
  assign _T_7126 = _T_7086 ? _T_7111 : _T_7125; // @[Mux.scala 31:69:@50410.4]
  assign _T_7127 = _T_7085 ? _T_7109 : _T_7126; // @[Mux.scala 31:69:@50411.4]
  assign _T_7128 = _T_7084 ? _T_7107 : _T_7127; // @[Mux.scala 31:69:@50412.4]
  assign _T_7129 = _T_7083 ? _T_7105 : _T_7128; // @[Mux.scala 31:69:@50413.4]
  assign _T_7130 = _T_7082 ? _T_7103 : _T_7129; // @[Mux.scala 31:69:@50414.4]
  assign _T_7131 = _T_7081 ? _T_7101 : _T_7130; // @[Mux.scala 31:69:@50415.4]
  assign _T_7132 = _T_7080 ? _T_7099 : _T_7131; // @[Mux.scala 31:69:@50416.4]
  assign _T_7133 = _T_7079 ? _T_7097 : _T_7132; // @[Mux.scala 31:69:@50417.4]
  assign _T_7134 = _T_7078 ? _T_7095 : _T_7133; // @[Mux.scala 31:69:@50418.4]
  assign _T_7135 = _T_7077 ? _T_7093 : _T_7134; // @[Mux.scala 31:69:@50419.4]
  assign _T_7143 = _T_5924 & _T_4102; // @[MemPrimitives.scala 110:228:@50428.4]
  assign _T_7149 = _T_5930 & _T_4108; // @[MemPrimitives.scala 110:228:@50432.4]
  assign _T_7155 = _T_5936 & _T_4114; // @[MemPrimitives.scala 110:228:@50436.4]
  assign _T_7161 = _T_5942 & _T_4120; // @[MemPrimitives.scala 110:228:@50440.4]
  assign _T_7167 = _T_5948 & _T_4126; // @[MemPrimitives.scala 110:228:@50444.4]
  assign _T_7173 = _T_5954 & _T_4132; // @[MemPrimitives.scala 110:228:@50448.4]
  assign _T_7179 = _T_5960 & _T_4138; // @[MemPrimitives.scala 110:228:@50452.4]
  assign _T_7185 = _T_5966 & _T_4144; // @[MemPrimitives.scala 110:228:@50456.4]
  assign _T_7191 = _T_5972 & _T_4150; // @[MemPrimitives.scala 110:228:@50460.4]
  assign _T_7197 = _T_5978 & _T_4156; // @[MemPrimitives.scala 110:228:@50464.4]
  assign _T_7203 = _T_5984 & _T_4162; // @[MemPrimitives.scala 110:228:@50468.4]
  assign _T_7209 = _T_5990 & _T_4168; // @[MemPrimitives.scala 110:228:@50472.4]
  assign _T_7215 = _T_5996 & _T_4174; // @[MemPrimitives.scala 110:228:@50476.4]
  assign _T_7221 = _T_6002 & _T_4180; // @[MemPrimitives.scala 110:228:@50480.4]
  assign _T_7227 = _T_6008 & _T_4186; // @[MemPrimitives.scala 110:228:@50484.4]
  assign _T_7229 = StickySelects_29_io_outs_0; // @[MemPrimitives.scala 123:41:@50504.4]
  assign _T_7230 = StickySelects_29_io_outs_1; // @[MemPrimitives.scala 123:41:@50505.4]
  assign _T_7231 = StickySelects_29_io_outs_2; // @[MemPrimitives.scala 123:41:@50506.4]
  assign _T_7232 = StickySelects_29_io_outs_3; // @[MemPrimitives.scala 123:41:@50507.4]
  assign _T_7233 = StickySelects_29_io_outs_4; // @[MemPrimitives.scala 123:41:@50508.4]
  assign _T_7234 = StickySelects_29_io_outs_5; // @[MemPrimitives.scala 123:41:@50509.4]
  assign _T_7235 = StickySelects_29_io_outs_6; // @[MemPrimitives.scala 123:41:@50510.4]
  assign _T_7236 = StickySelects_29_io_outs_7; // @[MemPrimitives.scala 123:41:@50511.4]
  assign _T_7237 = StickySelects_29_io_outs_8; // @[MemPrimitives.scala 123:41:@50512.4]
  assign _T_7238 = StickySelects_29_io_outs_9; // @[MemPrimitives.scala 123:41:@50513.4]
  assign _T_7239 = StickySelects_29_io_outs_10; // @[MemPrimitives.scala 123:41:@50514.4]
  assign _T_7240 = StickySelects_29_io_outs_11; // @[MemPrimitives.scala 123:41:@50515.4]
  assign _T_7241 = StickySelects_29_io_outs_12; // @[MemPrimitives.scala 123:41:@50516.4]
  assign _T_7242 = StickySelects_29_io_outs_13; // @[MemPrimitives.scala 123:41:@50517.4]
  assign _T_7243 = StickySelects_29_io_outs_14; // @[MemPrimitives.scala 123:41:@50518.4]
  assign _T_7245 = {_T_7229,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@50520.4]
  assign _T_7247 = {_T_7230,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@50522.4]
  assign _T_7249 = {_T_7231,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@50524.4]
  assign _T_7251 = {_T_7232,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@50526.4]
  assign _T_7253 = {_T_7233,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@50528.4]
  assign _T_7255 = {_T_7234,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@50530.4]
  assign _T_7257 = {_T_7235,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@50532.4]
  assign _T_7259 = {_T_7236,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@50534.4]
  assign _T_7261 = {_T_7237,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@50536.4]
  assign _T_7263 = {_T_7238,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@50538.4]
  assign _T_7265 = {_T_7239,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@50540.4]
  assign _T_7267 = {_T_7240,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@50542.4]
  assign _T_7269 = {_T_7241,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@50544.4]
  assign _T_7271 = {_T_7242,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@50546.4]
  assign _T_7273 = {_T_7243,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@50548.4]
  assign _T_7274 = _T_7242 ? _T_7271 : _T_7273; // @[Mux.scala 31:69:@50549.4]
  assign _T_7275 = _T_7241 ? _T_7269 : _T_7274; // @[Mux.scala 31:69:@50550.4]
  assign _T_7276 = _T_7240 ? _T_7267 : _T_7275; // @[Mux.scala 31:69:@50551.4]
  assign _T_7277 = _T_7239 ? _T_7265 : _T_7276; // @[Mux.scala 31:69:@50552.4]
  assign _T_7278 = _T_7238 ? _T_7263 : _T_7277; // @[Mux.scala 31:69:@50553.4]
  assign _T_7279 = _T_7237 ? _T_7261 : _T_7278; // @[Mux.scala 31:69:@50554.4]
  assign _T_7280 = _T_7236 ? _T_7259 : _T_7279; // @[Mux.scala 31:69:@50555.4]
  assign _T_7281 = _T_7235 ? _T_7257 : _T_7280; // @[Mux.scala 31:69:@50556.4]
  assign _T_7282 = _T_7234 ? _T_7255 : _T_7281; // @[Mux.scala 31:69:@50557.4]
  assign _T_7283 = _T_7233 ? _T_7253 : _T_7282; // @[Mux.scala 31:69:@50558.4]
  assign _T_7284 = _T_7232 ? _T_7251 : _T_7283; // @[Mux.scala 31:69:@50559.4]
  assign _T_7285 = _T_7231 ? _T_7249 : _T_7284; // @[Mux.scala 31:69:@50560.4]
  assign _T_7286 = _T_7230 ? _T_7247 : _T_7285; // @[Mux.scala 31:69:@50561.4]
  assign _T_7287 = _T_7229 ? _T_7245 : _T_7286; // @[Mux.scala 31:69:@50562.4]
  assign _T_7292 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50569.4]
  assign _T_7295 = _T_7292 & _T_2734; // @[MemPrimitives.scala 110:228:@50571.4]
  assign _T_7298 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50573.4]
  assign _T_7301 = _T_7298 & _T_2740; // @[MemPrimitives.scala 110:228:@50575.4]
  assign _T_7304 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50577.4]
  assign _T_7307 = _T_7304 & _T_2746; // @[MemPrimitives.scala 110:228:@50579.4]
  assign _T_7310 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50581.4]
  assign _T_7313 = _T_7310 & _T_2752; // @[MemPrimitives.scala 110:228:@50583.4]
  assign _T_7316 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50585.4]
  assign _T_7319 = _T_7316 & _T_2758; // @[MemPrimitives.scala 110:228:@50587.4]
  assign _T_7322 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50589.4]
  assign _T_7325 = _T_7322 & _T_2764; // @[MemPrimitives.scala 110:228:@50591.4]
  assign _T_7328 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50593.4]
  assign _T_7331 = _T_7328 & _T_2770; // @[MemPrimitives.scala 110:228:@50595.4]
  assign _T_7334 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50597.4]
  assign _T_7337 = _T_7334 & _T_2776; // @[MemPrimitives.scala 110:228:@50599.4]
  assign _T_7340 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50601.4]
  assign _T_7343 = _T_7340 & _T_2782; // @[MemPrimitives.scala 110:228:@50603.4]
  assign _T_7346 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50605.4]
  assign _T_7349 = _T_7346 & _T_2788; // @[MemPrimitives.scala 110:228:@50607.4]
  assign _T_7352 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50609.4]
  assign _T_7355 = _T_7352 & _T_2794; // @[MemPrimitives.scala 110:228:@50611.4]
  assign _T_7358 = io_rPort_19_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50613.4]
  assign _T_7361 = _T_7358 & _T_2800; // @[MemPrimitives.scala 110:228:@50615.4]
  assign _T_7364 = io_rPort_22_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50617.4]
  assign _T_7367 = _T_7364 & _T_2806; // @[MemPrimitives.scala 110:228:@50619.4]
  assign _T_7370 = io_rPort_26_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50621.4]
  assign _T_7373 = _T_7370 & _T_2812; // @[MemPrimitives.scala 110:228:@50623.4]
  assign _T_7376 = io_rPort_29_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50625.4]
  assign _T_7379 = _T_7376 & _T_2818; // @[MemPrimitives.scala 110:228:@50627.4]
  assign _T_7381 = StickySelects_30_io_outs_0; // @[MemPrimitives.scala 123:41:@50647.4]
  assign _T_7382 = StickySelects_30_io_outs_1; // @[MemPrimitives.scala 123:41:@50648.4]
  assign _T_7383 = StickySelects_30_io_outs_2; // @[MemPrimitives.scala 123:41:@50649.4]
  assign _T_7384 = StickySelects_30_io_outs_3; // @[MemPrimitives.scala 123:41:@50650.4]
  assign _T_7385 = StickySelects_30_io_outs_4; // @[MemPrimitives.scala 123:41:@50651.4]
  assign _T_7386 = StickySelects_30_io_outs_5; // @[MemPrimitives.scala 123:41:@50652.4]
  assign _T_7387 = StickySelects_30_io_outs_6; // @[MemPrimitives.scala 123:41:@50653.4]
  assign _T_7388 = StickySelects_30_io_outs_7; // @[MemPrimitives.scala 123:41:@50654.4]
  assign _T_7389 = StickySelects_30_io_outs_8; // @[MemPrimitives.scala 123:41:@50655.4]
  assign _T_7390 = StickySelects_30_io_outs_9; // @[MemPrimitives.scala 123:41:@50656.4]
  assign _T_7391 = StickySelects_30_io_outs_10; // @[MemPrimitives.scala 123:41:@50657.4]
  assign _T_7392 = StickySelects_30_io_outs_11; // @[MemPrimitives.scala 123:41:@50658.4]
  assign _T_7393 = StickySelects_30_io_outs_12; // @[MemPrimitives.scala 123:41:@50659.4]
  assign _T_7394 = StickySelects_30_io_outs_13; // @[MemPrimitives.scala 123:41:@50660.4]
  assign _T_7395 = StickySelects_30_io_outs_14; // @[MemPrimitives.scala 123:41:@50661.4]
  assign _T_7397 = {_T_7381,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@50663.4]
  assign _T_7399 = {_T_7382,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@50665.4]
  assign _T_7401 = {_T_7383,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@50667.4]
  assign _T_7403 = {_T_7384,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@50669.4]
  assign _T_7405 = {_T_7385,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@50671.4]
  assign _T_7407 = {_T_7386,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@50673.4]
  assign _T_7409 = {_T_7387,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@50675.4]
  assign _T_7411 = {_T_7388,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@50677.4]
  assign _T_7413 = {_T_7389,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@50679.4]
  assign _T_7415 = {_T_7390,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@50681.4]
  assign _T_7417 = {_T_7391,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@50683.4]
  assign _T_7419 = {_T_7392,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@50685.4]
  assign _T_7421 = {_T_7393,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@50687.4]
  assign _T_7423 = {_T_7394,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@50689.4]
  assign _T_7425 = {_T_7395,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@50691.4]
  assign _T_7426 = _T_7394 ? _T_7423 : _T_7425; // @[Mux.scala 31:69:@50692.4]
  assign _T_7427 = _T_7393 ? _T_7421 : _T_7426; // @[Mux.scala 31:69:@50693.4]
  assign _T_7428 = _T_7392 ? _T_7419 : _T_7427; // @[Mux.scala 31:69:@50694.4]
  assign _T_7429 = _T_7391 ? _T_7417 : _T_7428; // @[Mux.scala 31:69:@50695.4]
  assign _T_7430 = _T_7390 ? _T_7415 : _T_7429; // @[Mux.scala 31:69:@50696.4]
  assign _T_7431 = _T_7389 ? _T_7413 : _T_7430; // @[Mux.scala 31:69:@50697.4]
  assign _T_7432 = _T_7388 ? _T_7411 : _T_7431; // @[Mux.scala 31:69:@50698.4]
  assign _T_7433 = _T_7387 ? _T_7409 : _T_7432; // @[Mux.scala 31:69:@50699.4]
  assign _T_7434 = _T_7386 ? _T_7407 : _T_7433; // @[Mux.scala 31:69:@50700.4]
  assign _T_7435 = _T_7385 ? _T_7405 : _T_7434; // @[Mux.scala 31:69:@50701.4]
  assign _T_7436 = _T_7384 ? _T_7403 : _T_7435; // @[Mux.scala 31:69:@50702.4]
  assign _T_7437 = _T_7383 ? _T_7401 : _T_7436; // @[Mux.scala 31:69:@50703.4]
  assign _T_7438 = _T_7382 ? _T_7399 : _T_7437; // @[Mux.scala 31:69:@50704.4]
  assign _T_7439 = _T_7381 ? _T_7397 : _T_7438; // @[Mux.scala 31:69:@50705.4]
  assign _T_7444 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50712.4]
  assign _T_7447 = _T_7444 & _T_2886; // @[MemPrimitives.scala 110:228:@50714.4]
  assign _T_7450 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50716.4]
  assign _T_7453 = _T_7450 & _T_2892; // @[MemPrimitives.scala 110:228:@50718.4]
  assign _T_7456 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50720.4]
  assign _T_7459 = _T_7456 & _T_2898; // @[MemPrimitives.scala 110:228:@50722.4]
  assign _T_7462 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50724.4]
  assign _T_7465 = _T_7462 & _T_2904; // @[MemPrimitives.scala 110:228:@50726.4]
  assign _T_7468 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50728.4]
  assign _T_7471 = _T_7468 & _T_2910; // @[MemPrimitives.scala 110:228:@50730.4]
  assign _T_7474 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50732.4]
  assign _T_7477 = _T_7474 & _T_2916; // @[MemPrimitives.scala 110:228:@50734.4]
  assign _T_7480 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50736.4]
  assign _T_7483 = _T_7480 & _T_2922; // @[MemPrimitives.scala 110:228:@50738.4]
  assign _T_7486 = io_rPort_18_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50740.4]
  assign _T_7489 = _T_7486 & _T_2928; // @[MemPrimitives.scala 110:228:@50742.4]
  assign _T_7492 = io_rPort_20_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50744.4]
  assign _T_7495 = _T_7492 & _T_2934; // @[MemPrimitives.scala 110:228:@50746.4]
  assign _T_7498 = io_rPort_21_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50748.4]
  assign _T_7501 = _T_7498 & _T_2940; // @[MemPrimitives.scala 110:228:@50750.4]
  assign _T_7504 = io_rPort_23_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50752.4]
  assign _T_7507 = _T_7504 & _T_2946; // @[MemPrimitives.scala 110:228:@50754.4]
  assign _T_7510 = io_rPort_24_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50756.4]
  assign _T_7513 = _T_7510 & _T_2952; // @[MemPrimitives.scala 110:228:@50758.4]
  assign _T_7516 = io_rPort_25_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50760.4]
  assign _T_7519 = _T_7516 & _T_2958; // @[MemPrimitives.scala 110:228:@50762.4]
  assign _T_7522 = io_rPort_27_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50764.4]
  assign _T_7525 = _T_7522 & _T_2964; // @[MemPrimitives.scala 110:228:@50766.4]
  assign _T_7528 = io_rPort_28_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@50768.4]
  assign _T_7531 = _T_7528 & _T_2970; // @[MemPrimitives.scala 110:228:@50770.4]
  assign _T_7533 = StickySelects_31_io_outs_0; // @[MemPrimitives.scala 123:41:@50790.4]
  assign _T_7534 = StickySelects_31_io_outs_1; // @[MemPrimitives.scala 123:41:@50791.4]
  assign _T_7535 = StickySelects_31_io_outs_2; // @[MemPrimitives.scala 123:41:@50792.4]
  assign _T_7536 = StickySelects_31_io_outs_3; // @[MemPrimitives.scala 123:41:@50793.4]
  assign _T_7537 = StickySelects_31_io_outs_4; // @[MemPrimitives.scala 123:41:@50794.4]
  assign _T_7538 = StickySelects_31_io_outs_5; // @[MemPrimitives.scala 123:41:@50795.4]
  assign _T_7539 = StickySelects_31_io_outs_6; // @[MemPrimitives.scala 123:41:@50796.4]
  assign _T_7540 = StickySelects_31_io_outs_7; // @[MemPrimitives.scala 123:41:@50797.4]
  assign _T_7541 = StickySelects_31_io_outs_8; // @[MemPrimitives.scala 123:41:@50798.4]
  assign _T_7542 = StickySelects_31_io_outs_9; // @[MemPrimitives.scala 123:41:@50799.4]
  assign _T_7543 = StickySelects_31_io_outs_10; // @[MemPrimitives.scala 123:41:@50800.4]
  assign _T_7544 = StickySelects_31_io_outs_11; // @[MemPrimitives.scala 123:41:@50801.4]
  assign _T_7545 = StickySelects_31_io_outs_12; // @[MemPrimitives.scala 123:41:@50802.4]
  assign _T_7546 = StickySelects_31_io_outs_13; // @[MemPrimitives.scala 123:41:@50803.4]
  assign _T_7547 = StickySelects_31_io_outs_14; // @[MemPrimitives.scala 123:41:@50804.4]
  assign _T_7549 = {_T_7533,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@50806.4]
  assign _T_7551 = {_T_7534,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@50808.4]
  assign _T_7553 = {_T_7535,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@50810.4]
  assign _T_7555 = {_T_7536,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@50812.4]
  assign _T_7557 = {_T_7537,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@50814.4]
  assign _T_7559 = {_T_7538,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@50816.4]
  assign _T_7561 = {_T_7539,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@50818.4]
  assign _T_7563 = {_T_7540,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@50820.4]
  assign _T_7565 = {_T_7541,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@50822.4]
  assign _T_7567 = {_T_7542,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@50824.4]
  assign _T_7569 = {_T_7543,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@50826.4]
  assign _T_7571 = {_T_7544,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@50828.4]
  assign _T_7573 = {_T_7545,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@50830.4]
  assign _T_7575 = {_T_7546,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@50832.4]
  assign _T_7577 = {_T_7547,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@50834.4]
  assign _T_7578 = _T_7546 ? _T_7575 : _T_7577; // @[Mux.scala 31:69:@50835.4]
  assign _T_7579 = _T_7545 ? _T_7573 : _T_7578; // @[Mux.scala 31:69:@50836.4]
  assign _T_7580 = _T_7544 ? _T_7571 : _T_7579; // @[Mux.scala 31:69:@50837.4]
  assign _T_7581 = _T_7543 ? _T_7569 : _T_7580; // @[Mux.scala 31:69:@50838.4]
  assign _T_7582 = _T_7542 ? _T_7567 : _T_7581; // @[Mux.scala 31:69:@50839.4]
  assign _T_7583 = _T_7541 ? _T_7565 : _T_7582; // @[Mux.scala 31:69:@50840.4]
  assign _T_7584 = _T_7540 ? _T_7563 : _T_7583; // @[Mux.scala 31:69:@50841.4]
  assign _T_7585 = _T_7539 ? _T_7561 : _T_7584; // @[Mux.scala 31:69:@50842.4]
  assign _T_7586 = _T_7538 ? _T_7559 : _T_7585; // @[Mux.scala 31:69:@50843.4]
  assign _T_7587 = _T_7537 ? _T_7557 : _T_7586; // @[Mux.scala 31:69:@50844.4]
  assign _T_7588 = _T_7536 ? _T_7555 : _T_7587; // @[Mux.scala 31:69:@50845.4]
  assign _T_7589 = _T_7535 ? _T_7553 : _T_7588; // @[Mux.scala 31:69:@50846.4]
  assign _T_7590 = _T_7534 ? _T_7551 : _T_7589; // @[Mux.scala 31:69:@50847.4]
  assign _T_7591 = _T_7533 ? _T_7549 : _T_7590; // @[Mux.scala 31:69:@50848.4]
  assign _T_7599 = _T_7292 & _T_3038; // @[MemPrimitives.scala 110:228:@50857.4]
  assign _T_7605 = _T_7298 & _T_3044; // @[MemPrimitives.scala 110:228:@50861.4]
  assign _T_7611 = _T_7304 & _T_3050; // @[MemPrimitives.scala 110:228:@50865.4]
  assign _T_7617 = _T_7310 & _T_3056; // @[MemPrimitives.scala 110:228:@50869.4]
  assign _T_7623 = _T_7316 & _T_3062; // @[MemPrimitives.scala 110:228:@50873.4]
  assign _T_7629 = _T_7322 & _T_3068; // @[MemPrimitives.scala 110:228:@50877.4]
  assign _T_7635 = _T_7328 & _T_3074; // @[MemPrimitives.scala 110:228:@50881.4]
  assign _T_7641 = _T_7334 & _T_3080; // @[MemPrimitives.scala 110:228:@50885.4]
  assign _T_7647 = _T_7340 & _T_3086; // @[MemPrimitives.scala 110:228:@50889.4]
  assign _T_7653 = _T_7346 & _T_3092; // @[MemPrimitives.scala 110:228:@50893.4]
  assign _T_7659 = _T_7352 & _T_3098; // @[MemPrimitives.scala 110:228:@50897.4]
  assign _T_7665 = _T_7358 & _T_3104; // @[MemPrimitives.scala 110:228:@50901.4]
  assign _T_7671 = _T_7364 & _T_3110; // @[MemPrimitives.scala 110:228:@50905.4]
  assign _T_7677 = _T_7370 & _T_3116; // @[MemPrimitives.scala 110:228:@50909.4]
  assign _T_7683 = _T_7376 & _T_3122; // @[MemPrimitives.scala 110:228:@50913.4]
  assign _T_7685 = StickySelects_32_io_outs_0; // @[MemPrimitives.scala 123:41:@50933.4]
  assign _T_7686 = StickySelects_32_io_outs_1; // @[MemPrimitives.scala 123:41:@50934.4]
  assign _T_7687 = StickySelects_32_io_outs_2; // @[MemPrimitives.scala 123:41:@50935.4]
  assign _T_7688 = StickySelects_32_io_outs_3; // @[MemPrimitives.scala 123:41:@50936.4]
  assign _T_7689 = StickySelects_32_io_outs_4; // @[MemPrimitives.scala 123:41:@50937.4]
  assign _T_7690 = StickySelects_32_io_outs_5; // @[MemPrimitives.scala 123:41:@50938.4]
  assign _T_7691 = StickySelects_32_io_outs_6; // @[MemPrimitives.scala 123:41:@50939.4]
  assign _T_7692 = StickySelects_32_io_outs_7; // @[MemPrimitives.scala 123:41:@50940.4]
  assign _T_7693 = StickySelects_32_io_outs_8; // @[MemPrimitives.scala 123:41:@50941.4]
  assign _T_7694 = StickySelects_32_io_outs_9; // @[MemPrimitives.scala 123:41:@50942.4]
  assign _T_7695 = StickySelects_32_io_outs_10; // @[MemPrimitives.scala 123:41:@50943.4]
  assign _T_7696 = StickySelects_32_io_outs_11; // @[MemPrimitives.scala 123:41:@50944.4]
  assign _T_7697 = StickySelects_32_io_outs_12; // @[MemPrimitives.scala 123:41:@50945.4]
  assign _T_7698 = StickySelects_32_io_outs_13; // @[MemPrimitives.scala 123:41:@50946.4]
  assign _T_7699 = StickySelects_32_io_outs_14; // @[MemPrimitives.scala 123:41:@50947.4]
  assign _T_7701 = {_T_7685,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@50949.4]
  assign _T_7703 = {_T_7686,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@50951.4]
  assign _T_7705 = {_T_7687,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@50953.4]
  assign _T_7707 = {_T_7688,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@50955.4]
  assign _T_7709 = {_T_7689,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@50957.4]
  assign _T_7711 = {_T_7690,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@50959.4]
  assign _T_7713 = {_T_7691,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@50961.4]
  assign _T_7715 = {_T_7692,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@50963.4]
  assign _T_7717 = {_T_7693,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@50965.4]
  assign _T_7719 = {_T_7694,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@50967.4]
  assign _T_7721 = {_T_7695,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@50969.4]
  assign _T_7723 = {_T_7696,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@50971.4]
  assign _T_7725 = {_T_7697,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@50973.4]
  assign _T_7727 = {_T_7698,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@50975.4]
  assign _T_7729 = {_T_7699,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@50977.4]
  assign _T_7730 = _T_7698 ? _T_7727 : _T_7729; // @[Mux.scala 31:69:@50978.4]
  assign _T_7731 = _T_7697 ? _T_7725 : _T_7730; // @[Mux.scala 31:69:@50979.4]
  assign _T_7732 = _T_7696 ? _T_7723 : _T_7731; // @[Mux.scala 31:69:@50980.4]
  assign _T_7733 = _T_7695 ? _T_7721 : _T_7732; // @[Mux.scala 31:69:@50981.4]
  assign _T_7734 = _T_7694 ? _T_7719 : _T_7733; // @[Mux.scala 31:69:@50982.4]
  assign _T_7735 = _T_7693 ? _T_7717 : _T_7734; // @[Mux.scala 31:69:@50983.4]
  assign _T_7736 = _T_7692 ? _T_7715 : _T_7735; // @[Mux.scala 31:69:@50984.4]
  assign _T_7737 = _T_7691 ? _T_7713 : _T_7736; // @[Mux.scala 31:69:@50985.4]
  assign _T_7738 = _T_7690 ? _T_7711 : _T_7737; // @[Mux.scala 31:69:@50986.4]
  assign _T_7739 = _T_7689 ? _T_7709 : _T_7738; // @[Mux.scala 31:69:@50987.4]
  assign _T_7740 = _T_7688 ? _T_7707 : _T_7739; // @[Mux.scala 31:69:@50988.4]
  assign _T_7741 = _T_7687 ? _T_7705 : _T_7740; // @[Mux.scala 31:69:@50989.4]
  assign _T_7742 = _T_7686 ? _T_7703 : _T_7741; // @[Mux.scala 31:69:@50990.4]
  assign _T_7743 = _T_7685 ? _T_7701 : _T_7742; // @[Mux.scala 31:69:@50991.4]
  assign _T_7751 = _T_7444 & _T_3190; // @[MemPrimitives.scala 110:228:@51000.4]
  assign _T_7757 = _T_7450 & _T_3196; // @[MemPrimitives.scala 110:228:@51004.4]
  assign _T_7763 = _T_7456 & _T_3202; // @[MemPrimitives.scala 110:228:@51008.4]
  assign _T_7769 = _T_7462 & _T_3208; // @[MemPrimitives.scala 110:228:@51012.4]
  assign _T_7775 = _T_7468 & _T_3214; // @[MemPrimitives.scala 110:228:@51016.4]
  assign _T_7781 = _T_7474 & _T_3220; // @[MemPrimitives.scala 110:228:@51020.4]
  assign _T_7787 = _T_7480 & _T_3226; // @[MemPrimitives.scala 110:228:@51024.4]
  assign _T_7793 = _T_7486 & _T_3232; // @[MemPrimitives.scala 110:228:@51028.4]
  assign _T_7799 = _T_7492 & _T_3238; // @[MemPrimitives.scala 110:228:@51032.4]
  assign _T_7805 = _T_7498 & _T_3244; // @[MemPrimitives.scala 110:228:@51036.4]
  assign _T_7811 = _T_7504 & _T_3250; // @[MemPrimitives.scala 110:228:@51040.4]
  assign _T_7817 = _T_7510 & _T_3256; // @[MemPrimitives.scala 110:228:@51044.4]
  assign _T_7823 = _T_7516 & _T_3262; // @[MemPrimitives.scala 110:228:@51048.4]
  assign _T_7829 = _T_7522 & _T_3268; // @[MemPrimitives.scala 110:228:@51052.4]
  assign _T_7835 = _T_7528 & _T_3274; // @[MemPrimitives.scala 110:228:@51056.4]
  assign _T_7837 = StickySelects_33_io_outs_0; // @[MemPrimitives.scala 123:41:@51076.4]
  assign _T_7838 = StickySelects_33_io_outs_1; // @[MemPrimitives.scala 123:41:@51077.4]
  assign _T_7839 = StickySelects_33_io_outs_2; // @[MemPrimitives.scala 123:41:@51078.4]
  assign _T_7840 = StickySelects_33_io_outs_3; // @[MemPrimitives.scala 123:41:@51079.4]
  assign _T_7841 = StickySelects_33_io_outs_4; // @[MemPrimitives.scala 123:41:@51080.4]
  assign _T_7842 = StickySelects_33_io_outs_5; // @[MemPrimitives.scala 123:41:@51081.4]
  assign _T_7843 = StickySelects_33_io_outs_6; // @[MemPrimitives.scala 123:41:@51082.4]
  assign _T_7844 = StickySelects_33_io_outs_7; // @[MemPrimitives.scala 123:41:@51083.4]
  assign _T_7845 = StickySelects_33_io_outs_8; // @[MemPrimitives.scala 123:41:@51084.4]
  assign _T_7846 = StickySelects_33_io_outs_9; // @[MemPrimitives.scala 123:41:@51085.4]
  assign _T_7847 = StickySelects_33_io_outs_10; // @[MemPrimitives.scala 123:41:@51086.4]
  assign _T_7848 = StickySelects_33_io_outs_11; // @[MemPrimitives.scala 123:41:@51087.4]
  assign _T_7849 = StickySelects_33_io_outs_12; // @[MemPrimitives.scala 123:41:@51088.4]
  assign _T_7850 = StickySelects_33_io_outs_13; // @[MemPrimitives.scala 123:41:@51089.4]
  assign _T_7851 = StickySelects_33_io_outs_14; // @[MemPrimitives.scala 123:41:@51090.4]
  assign _T_7853 = {_T_7837,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@51092.4]
  assign _T_7855 = {_T_7838,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@51094.4]
  assign _T_7857 = {_T_7839,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@51096.4]
  assign _T_7859 = {_T_7840,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@51098.4]
  assign _T_7861 = {_T_7841,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@51100.4]
  assign _T_7863 = {_T_7842,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@51102.4]
  assign _T_7865 = {_T_7843,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@51104.4]
  assign _T_7867 = {_T_7844,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@51106.4]
  assign _T_7869 = {_T_7845,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@51108.4]
  assign _T_7871 = {_T_7846,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@51110.4]
  assign _T_7873 = {_T_7847,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@51112.4]
  assign _T_7875 = {_T_7848,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@51114.4]
  assign _T_7877 = {_T_7849,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@51116.4]
  assign _T_7879 = {_T_7850,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@51118.4]
  assign _T_7881 = {_T_7851,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@51120.4]
  assign _T_7882 = _T_7850 ? _T_7879 : _T_7881; // @[Mux.scala 31:69:@51121.4]
  assign _T_7883 = _T_7849 ? _T_7877 : _T_7882; // @[Mux.scala 31:69:@51122.4]
  assign _T_7884 = _T_7848 ? _T_7875 : _T_7883; // @[Mux.scala 31:69:@51123.4]
  assign _T_7885 = _T_7847 ? _T_7873 : _T_7884; // @[Mux.scala 31:69:@51124.4]
  assign _T_7886 = _T_7846 ? _T_7871 : _T_7885; // @[Mux.scala 31:69:@51125.4]
  assign _T_7887 = _T_7845 ? _T_7869 : _T_7886; // @[Mux.scala 31:69:@51126.4]
  assign _T_7888 = _T_7844 ? _T_7867 : _T_7887; // @[Mux.scala 31:69:@51127.4]
  assign _T_7889 = _T_7843 ? _T_7865 : _T_7888; // @[Mux.scala 31:69:@51128.4]
  assign _T_7890 = _T_7842 ? _T_7863 : _T_7889; // @[Mux.scala 31:69:@51129.4]
  assign _T_7891 = _T_7841 ? _T_7861 : _T_7890; // @[Mux.scala 31:69:@51130.4]
  assign _T_7892 = _T_7840 ? _T_7859 : _T_7891; // @[Mux.scala 31:69:@51131.4]
  assign _T_7893 = _T_7839 ? _T_7857 : _T_7892; // @[Mux.scala 31:69:@51132.4]
  assign _T_7894 = _T_7838 ? _T_7855 : _T_7893; // @[Mux.scala 31:69:@51133.4]
  assign _T_7895 = _T_7837 ? _T_7853 : _T_7894; // @[Mux.scala 31:69:@51134.4]
  assign _T_7903 = _T_7292 & _T_3342; // @[MemPrimitives.scala 110:228:@51143.4]
  assign _T_7909 = _T_7298 & _T_3348; // @[MemPrimitives.scala 110:228:@51147.4]
  assign _T_7915 = _T_7304 & _T_3354; // @[MemPrimitives.scala 110:228:@51151.4]
  assign _T_7921 = _T_7310 & _T_3360; // @[MemPrimitives.scala 110:228:@51155.4]
  assign _T_7927 = _T_7316 & _T_3366; // @[MemPrimitives.scala 110:228:@51159.4]
  assign _T_7933 = _T_7322 & _T_3372; // @[MemPrimitives.scala 110:228:@51163.4]
  assign _T_7939 = _T_7328 & _T_3378; // @[MemPrimitives.scala 110:228:@51167.4]
  assign _T_7945 = _T_7334 & _T_3384; // @[MemPrimitives.scala 110:228:@51171.4]
  assign _T_7951 = _T_7340 & _T_3390; // @[MemPrimitives.scala 110:228:@51175.4]
  assign _T_7957 = _T_7346 & _T_3396; // @[MemPrimitives.scala 110:228:@51179.4]
  assign _T_7963 = _T_7352 & _T_3402; // @[MemPrimitives.scala 110:228:@51183.4]
  assign _T_7969 = _T_7358 & _T_3408; // @[MemPrimitives.scala 110:228:@51187.4]
  assign _T_7975 = _T_7364 & _T_3414; // @[MemPrimitives.scala 110:228:@51191.4]
  assign _T_7981 = _T_7370 & _T_3420; // @[MemPrimitives.scala 110:228:@51195.4]
  assign _T_7987 = _T_7376 & _T_3426; // @[MemPrimitives.scala 110:228:@51199.4]
  assign _T_7989 = StickySelects_34_io_outs_0; // @[MemPrimitives.scala 123:41:@51219.4]
  assign _T_7990 = StickySelects_34_io_outs_1; // @[MemPrimitives.scala 123:41:@51220.4]
  assign _T_7991 = StickySelects_34_io_outs_2; // @[MemPrimitives.scala 123:41:@51221.4]
  assign _T_7992 = StickySelects_34_io_outs_3; // @[MemPrimitives.scala 123:41:@51222.4]
  assign _T_7993 = StickySelects_34_io_outs_4; // @[MemPrimitives.scala 123:41:@51223.4]
  assign _T_7994 = StickySelects_34_io_outs_5; // @[MemPrimitives.scala 123:41:@51224.4]
  assign _T_7995 = StickySelects_34_io_outs_6; // @[MemPrimitives.scala 123:41:@51225.4]
  assign _T_7996 = StickySelects_34_io_outs_7; // @[MemPrimitives.scala 123:41:@51226.4]
  assign _T_7997 = StickySelects_34_io_outs_8; // @[MemPrimitives.scala 123:41:@51227.4]
  assign _T_7998 = StickySelects_34_io_outs_9; // @[MemPrimitives.scala 123:41:@51228.4]
  assign _T_7999 = StickySelects_34_io_outs_10; // @[MemPrimitives.scala 123:41:@51229.4]
  assign _T_8000 = StickySelects_34_io_outs_11; // @[MemPrimitives.scala 123:41:@51230.4]
  assign _T_8001 = StickySelects_34_io_outs_12; // @[MemPrimitives.scala 123:41:@51231.4]
  assign _T_8002 = StickySelects_34_io_outs_13; // @[MemPrimitives.scala 123:41:@51232.4]
  assign _T_8003 = StickySelects_34_io_outs_14; // @[MemPrimitives.scala 123:41:@51233.4]
  assign _T_8005 = {_T_7989,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@51235.4]
  assign _T_8007 = {_T_7990,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@51237.4]
  assign _T_8009 = {_T_7991,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@51239.4]
  assign _T_8011 = {_T_7992,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@51241.4]
  assign _T_8013 = {_T_7993,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@51243.4]
  assign _T_8015 = {_T_7994,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@51245.4]
  assign _T_8017 = {_T_7995,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@51247.4]
  assign _T_8019 = {_T_7996,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@51249.4]
  assign _T_8021 = {_T_7997,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@51251.4]
  assign _T_8023 = {_T_7998,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@51253.4]
  assign _T_8025 = {_T_7999,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@51255.4]
  assign _T_8027 = {_T_8000,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@51257.4]
  assign _T_8029 = {_T_8001,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@51259.4]
  assign _T_8031 = {_T_8002,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@51261.4]
  assign _T_8033 = {_T_8003,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@51263.4]
  assign _T_8034 = _T_8002 ? _T_8031 : _T_8033; // @[Mux.scala 31:69:@51264.4]
  assign _T_8035 = _T_8001 ? _T_8029 : _T_8034; // @[Mux.scala 31:69:@51265.4]
  assign _T_8036 = _T_8000 ? _T_8027 : _T_8035; // @[Mux.scala 31:69:@51266.4]
  assign _T_8037 = _T_7999 ? _T_8025 : _T_8036; // @[Mux.scala 31:69:@51267.4]
  assign _T_8038 = _T_7998 ? _T_8023 : _T_8037; // @[Mux.scala 31:69:@51268.4]
  assign _T_8039 = _T_7997 ? _T_8021 : _T_8038; // @[Mux.scala 31:69:@51269.4]
  assign _T_8040 = _T_7996 ? _T_8019 : _T_8039; // @[Mux.scala 31:69:@51270.4]
  assign _T_8041 = _T_7995 ? _T_8017 : _T_8040; // @[Mux.scala 31:69:@51271.4]
  assign _T_8042 = _T_7994 ? _T_8015 : _T_8041; // @[Mux.scala 31:69:@51272.4]
  assign _T_8043 = _T_7993 ? _T_8013 : _T_8042; // @[Mux.scala 31:69:@51273.4]
  assign _T_8044 = _T_7992 ? _T_8011 : _T_8043; // @[Mux.scala 31:69:@51274.4]
  assign _T_8045 = _T_7991 ? _T_8009 : _T_8044; // @[Mux.scala 31:69:@51275.4]
  assign _T_8046 = _T_7990 ? _T_8007 : _T_8045; // @[Mux.scala 31:69:@51276.4]
  assign _T_8047 = _T_7989 ? _T_8005 : _T_8046; // @[Mux.scala 31:69:@51277.4]
  assign _T_8055 = _T_7444 & _T_3494; // @[MemPrimitives.scala 110:228:@51286.4]
  assign _T_8061 = _T_7450 & _T_3500; // @[MemPrimitives.scala 110:228:@51290.4]
  assign _T_8067 = _T_7456 & _T_3506; // @[MemPrimitives.scala 110:228:@51294.4]
  assign _T_8073 = _T_7462 & _T_3512; // @[MemPrimitives.scala 110:228:@51298.4]
  assign _T_8079 = _T_7468 & _T_3518; // @[MemPrimitives.scala 110:228:@51302.4]
  assign _T_8085 = _T_7474 & _T_3524; // @[MemPrimitives.scala 110:228:@51306.4]
  assign _T_8091 = _T_7480 & _T_3530; // @[MemPrimitives.scala 110:228:@51310.4]
  assign _T_8097 = _T_7486 & _T_3536; // @[MemPrimitives.scala 110:228:@51314.4]
  assign _T_8103 = _T_7492 & _T_3542; // @[MemPrimitives.scala 110:228:@51318.4]
  assign _T_8109 = _T_7498 & _T_3548; // @[MemPrimitives.scala 110:228:@51322.4]
  assign _T_8115 = _T_7504 & _T_3554; // @[MemPrimitives.scala 110:228:@51326.4]
  assign _T_8121 = _T_7510 & _T_3560; // @[MemPrimitives.scala 110:228:@51330.4]
  assign _T_8127 = _T_7516 & _T_3566; // @[MemPrimitives.scala 110:228:@51334.4]
  assign _T_8133 = _T_7522 & _T_3572; // @[MemPrimitives.scala 110:228:@51338.4]
  assign _T_8139 = _T_7528 & _T_3578; // @[MemPrimitives.scala 110:228:@51342.4]
  assign _T_8141 = StickySelects_35_io_outs_0; // @[MemPrimitives.scala 123:41:@51362.4]
  assign _T_8142 = StickySelects_35_io_outs_1; // @[MemPrimitives.scala 123:41:@51363.4]
  assign _T_8143 = StickySelects_35_io_outs_2; // @[MemPrimitives.scala 123:41:@51364.4]
  assign _T_8144 = StickySelects_35_io_outs_3; // @[MemPrimitives.scala 123:41:@51365.4]
  assign _T_8145 = StickySelects_35_io_outs_4; // @[MemPrimitives.scala 123:41:@51366.4]
  assign _T_8146 = StickySelects_35_io_outs_5; // @[MemPrimitives.scala 123:41:@51367.4]
  assign _T_8147 = StickySelects_35_io_outs_6; // @[MemPrimitives.scala 123:41:@51368.4]
  assign _T_8148 = StickySelects_35_io_outs_7; // @[MemPrimitives.scala 123:41:@51369.4]
  assign _T_8149 = StickySelects_35_io_outs_8; // @[MemPrimitives.scala 123:41:@51370.4]
  assign _T_8150 = StickySelects_35_io_outs_9; // @[MemPrimitives.scala 123:41:@51371.4]
  assign _T_8151 = StickySelects_35_io_outs_10; // @[MemPrimitives.scala 123:41:@51372.4]
  assign _T_8152 = StickySelects_35_io_outs_11; // @[MemPrimitives.scala 123:41:@51373.4]
  assign _T_8153 = StickySelects_35_io_outs_12; // @[MemPrimitives.scala 123:41:@51374.4]
  assign _T_8154 = StickySelects_35_io_outs_13; // @[MemPrimitives.scala 123:41:@51375.4]
  assign _T_8155 = StickySelects_35_io_outs_14; // @[MemPrimitives.scala 123:41:@51376.4]
  assign _T_8157 = {_T_8141,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@51378.4]
  assign _T_8159 = {_T_8142,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@51380.4]
  assign _T_8161 = {_T_8143,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@51382.4]
  assign _T_8163 = {_T_8144,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@51384.4]
  assign _T_8165 = {_T_8145,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@51386.4]
  assign _T_8167 = {_T_8146,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@51388.4]
  assign _T_8169 = {_T_8147,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@51390.4]
  assign _T_8171 = {_T_8148,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@51392.4]
  assign _T_8173 = {_T_8149,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@51394.4]
  assign _T_8175 = {_T_8150,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@51396.4]
  assign _T_8177 = {_T_8151,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@51398.4]
  assign _T_8179 = {_T_8152,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@51400.4]
  assign _T_8181 = {_T_8153,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@51402.4]
  assign _T_8183 = {_T_8154,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@51404.4]
  assign _T_8185 = {_T_8155,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@51406.4]
  assign _T_8186 = _T_8154 ? _T_8183 : _T_8185; // @[Mux.scala 31:69:@51407.4]
  assign _T_8187 = _T_8153 ? _T_8181 : _T_8186; // @[Mux.scala 31:69:@51408.4]
  assign _T_8188 = _T_8152 ? _T_8179 : _T_8187; // @[Mux.scala 31:69:@51409.4]
  assign _T_8189 = _T_8151 ? _T_8177 : _T_8188; // @[Mux.scala 31:69:@51410.4]
  assign _T_8190 = _T_8150 ? _T_8175 : _T_8189; // @[Mux.scala 31:69:@51411.4]
  assign _T_8191 = _T_8149 ? _T_8173 : _T_8190; // @[Mux.scala 31:69:@51412.4]
  assign _T_8192 = _T_8148 ? _T_8171 : _T_8191; // @[Mux.scala 31:69:@51413.4]
  assign _T_8193 = _T_8147 ? _T_8169 : _T_8192; // @[Mux.scala 31:69:@51414.4]
  assign _T_8194 = _T_8146 ? _T_8167 : _T_8193; // @[Mux.scala 31:69:@51415.4]
  assign _T_8195 = _T_8145 ? _T_8165 : _T_8194; // @[Mux.scala 31:69:@51416.4]
  assign _T_8196 = _T_8144 ? _T_8163 : _T_8195; // @[Mux.scala 31:69:@51417.4]
  assign _T_8197 = _T_8143 ? _T_8161 : _T_8196; // @[Mux.scala 31:69:@51418.4]
  assign _T_8198 = _T_8142 ? _T_8159 : _T_8197; // @[Mux.scala 31:69:@51419.4]
  assign _T_8199 = _T_8141 ? _T_8157 : _T_8198; // @[Mux.scala 31:69:@51420.4]
  assign _T_8207 = _T_7292 & _T_3646; // @[MemPrimitives.scala 110:228:@51429.4]
  assign _T_8213 = _T_7298 & _T_3652; // @[MemPrimitives.scala 110:228:@51433.4]
  assign _T_8219 = _T_7304 & _T_3658; // @[MemPrimitives.scala 110:228:@51437.4]
  assign _T_8225 = _T_7310 & _T_3664; // @[MemPrimitives.scala 110:228:@51441.4]
  assign _T_8231 = _T_7316 & _T_3670; // @[MemPrimitives.scala 110:228:@51445.4]
  assign _T_8237 = _T_7322 & _T_3676; // @[MemPrimitives.scala 110:228:@51449.4]
  assign _T_8243 = _T_7328 & _T_3682; // @[MemPrimitives.scala 110:228:@51453.4]
  assign _T_8249 = _T_7334 & _T_3688; // @[MemPrimitives.scala 110:228:@51457.4]
  assign _T_8255 = _T_7340 & _T_3694; // @[MemPrimitives.scala 110:228:@51461.4]
  assign _T_8261 = _T_7346 & _T_3700; // @[MemPrimitives.scala 110:228:@51465.4]
  assign _T_8267 = _T_7352 & _T_3706; // @[MemPrimitives.scala 110:228:@51469.4]
  assign _T_8273 = _T_7358 & _T_3712; // @[MemPrimitives.scala 110:228:@51473.4]
  assign _T_8279 = _T_7364 & _T_3718; // @[MemPrimitives.scala 110:228:@51477.4]
  assign _T_8285 = _T_7370 & _T_3724; // @[MemPrimitives.scala 110:228:@51481.4]
  assign _T_8291 = _T_7376 & _T_3730; // @[MemPrimitives.scala 110:228:@51485.4]
  assign _T_8293 = StickySelects_36_io_outs_0; // @[MemPrimitives.scala 123:41:@51505.4]
  assign _T_8294 = StickySelects_36_io_outs_1; // @[MemPrimitives.scala 123:41:@51506.4]
  assign _T_8295 = StickySelects_36_io_outs_2; // @[MemPrimitives.scala 123:41:@51507.4]
  assign _T_8296 = StickySelects_36_io_outs_3; // @[MemPrimitives.scala 123:41:@51508.4]
  assign _T_8297 = StickySelects_36_io_outs_4; // @[MemPrimitives.scala 123:41:@51509.4]
  assign _T_8298 = StickySelects_36_io_outs_5; // @[MemPrimitives.scala 123:41:@51510.4]
  assign _T_8299 = StickySelects_36_io_outs_6; // @[MemPrimitives.scala 123:41:@51511.4]
  assign _T_8300 = StickySelects_36_io_outs_7; // @[MemPrimitives.scala 123:41:@51512.4]
  assign _T_8301 = StickySelects_36_io_outs_8; // @[MemPrimitives.scala 123:41:@51513.4]
  assign _T_8302 = StickySelects_36_io_outs_9; // @[MemPrimitives.scala 123:41:@51514.4]
  assign _T_8303 = StickySelects_36_io_outs_10; // @[MemPrimitives.scala 123:41:@51515.4]
  assign _T_8304 = StickySelects_36_io_outs_11; // @[MemPrimitives.scala 123:41:@51516.4]
  assign _T_8305 = StickySelects_36_io_outs_12; // @[MemPrimitives.scala 123:41:@51517.4]
  assign _T_8306 = StickySelects_36_io_outs_13; // @[MemPrimitives.scala 123:41:@51518.4]
  assign _T_8307 = StickySelects_36_io_outs_14; // @[MemPrimitives.scala 123:41:@51519.4]
  assign _T_8309 = {_T_8293,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@51521.4]
  assign _T_8311 = {_T_8294,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@51523.4]
  assign _T_8313 = {_T_8295,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@51525.4]
  assign _T_8315 = {_T_8296,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@51527.4]
  assign _T_8317 = {_T_8297,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@51529.4]
  assign _T_8319 = {_T_8298,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@51531.4]
  assign _T_8321 = {_T_8299,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@51533.4]
  assign _T_8323 = {_T_8300,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@51535.4]
  assign _T_8325 = {_T_8301,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@51537.4]
  assign _T_8327 = {_T_8302,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@51539.4]
  assign _T_8329 = {_T_8303,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@51541.4]
  assign _T_8331 = {_T_8304,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@51543.4]
  assign _T_8333 = {_T_8305,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@51545.4]
  assign _T_8335 = {_T_8306,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@51547.4]
  assign _T_8337 = {_T_8307,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@51549.4]
  assign _T_8338 = _T_8306 ? _T_8335 : _T_8337; // @[Mux.scala 31:69:@51550.4]
  assign _T_8339 = _T_8305 ? _T_8333 : _T_8338; // @[Mux.scala 31:69:@51551.4]
  assign _T_8340 = _T_8304 ? _T_8331 : _T_8339; // @[Mux.scala 31:69:@51552.4]
  assign _T_8341 = _T_8303 ? _T_8329 : _T_8340; // @[Mux.scala 31:69:@51553.4]
  assign _T_8342 = _T_8302 ? _T_8327 : _T_8341; // @[Mux.scala 31:69:@51554.4]
  assign _T_8343 = _T_8301 ? _T_8325 : _T_8342; // @[Mux.scala 31:69:@51555.4]
  assign _T_8344 = _T_8300 ? _T_8323 : _T_8343; // @[Mux.scala 31:69:@51556.4]
  assign _T_8345 = _T_8299 ? _T_8321 : _T_8344; // @[Mux.scala 31:69:@51557.4]
  assign _T_8346 = _T_8298 ? _T_8319 : _T_8345; // @[Mux.scala 31:69:@51558.4]
  assign _T_8347 = _T_8297 ? _T_8317 : _T_8346; // @[Mux.scala 31:69:@51559.4]
  assign _T_8348 = _T_8296 ? _T_8315 : _T_8347; // @[Mux.scala 31:69:@51560.4]
  assign _T_8349 = _T_8295 ? _T_8313 : _T_8348; // @[Mux.scala 31:69:@51561.4]
  assign _T_8350 = _T_8294 ? _T_8311 : _T_8349; // @[Mux.scala 31:69:@51562.4]
  assign _T_8351 = _T_8293 ? _T_8309 : _T_8350; // @[Mux.scala 31:69:@51563.4]
  assign _T_8359 = _T_7444 & _T_3798; // @[MemPrimitives.scala 110:228:@51572.4]
  assign _T_8365 = _T_7450 & _T_3804; // @[MemPrimitives.scala 110:228:@51576.4]
  assign _T_8371 = _T_7456 & _T_3810; // @[MemPrimitives.scala 110:228:@51580.4]
  assign _T_8377 = _T_7462 & _T_3816; // @[MemPrimitives.scala 110:228:@51584.4]
  assign _T_8383 = _T_7468 & _T_3822; // @[MemPrimitives.scala 110:228:@51588.4]
  assign _T_8389 = _T_7474 & _T_3828; // @[MemPrimitives.scala 110:228:@51592.4]
  assign _T_8395 = _T_7480 & _T_3834; // @[MemPrimitives.scala 110:228:@51596.4]
  assign _T_8401 = _T_7486 & _T_3840; // @[MemPrimitives.scala 110:228:@51600.4]
  assign _T_8407 = _T_7492 & _T_3846; // @[MemPrimitives.scala 110:228:@51604.4]
  assign _T_8413 = _T_7498 & _T_3852; // @[MemPrimitives.scala 110:228:@51608.4]
  assign _T_8419 = _T_7504 & _T_3858; // @[MemPrimitives.scala 110:228:@51612.4]
  assign _T_8425 = _T_7510 & _T_3864; // @[MemPrimitives.scala 110:228:@51616.4]
  assign _T_8431 = _T_7516 & _T_3870; // @[MemPrimitives.scala 110:228:@51620.4]
  assign _T_8437 = _T_7522 & _T_3876; // @[MemPrimitives.scala 110:228:@51624.4]
  assign _T_8443 = _T_7528 & _T_3882; // @[MemPrimitives.scala 110:228:@51628.4]
  assign _T_8445 = StickySelects_37_io_outs_0; // @[MemPrimitives.scala 123:41:@51648.4]
  assign _T_8446 = StickySelects_37_io_outs_1; // @[MemPrimitives.scala 123:41:@51649.4]
  assign _T_8447 = StickySelects_37_io_outs_2; // @[MemPrimitives.scala 123:41:@51650.4]
  assign _T_8448 = StickySelects_37_io_outs_3; // @[MemPrimitives.scala 123:41:@51651.4]
  assign _T_8449 = StickySelects_37_io_outs_4; // @[MemPrimitives.scala 123:41:@51652.4]
  assign _T_8450 = StickySelects_37_io_outs_5; // @[MemPrimitives.scala 123:41:@51653.4]
  assign _T_8451 = StickySelects_37_io_outs_6; // @[MemPrimitives.scala 123:41:@51654.4]
  assign _T_8452 = StickySelects_37_io_outs_7; // @[MemPrimitives.scala 123:41:@51655.4]
  assign _T_8453 = StickySelects_37_io_outs_8; // @[MemPrimitives.scala 123:41:@51656.4]
  assign _T_8454 = StickySelects_37_io_outs_9; // @[MemPrimitives.scala 123:41:@51657.4]
  assign _T_8455 = StickySelects_37_io_outs_10; // @[MemPrimitives.scala 123:41:@51658.4]
  assign _T_8456 = StickySelects_37_io_outs_11; // @[MemPrimitives.scala 123:41:@51659.4]
  assign _T_8457 = StickySelects_37_io_outs_12; // @[MemPrimitives.scala 123:41:@51660.4]
  assign _T_8458 = StickySelects_37_io_outs_13; // @[MemPrimitives.scala 123:41:@51661.4]
  assign _T_8459 = StickySelects_37_io_outs_14; // @[MemPrimitives.scala 123:41:@51662.4]
  assign _T_8461 = {_T_8445,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@51664.4]
  assign _T_8463 = {_T_8446,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@51666.4]
  assign _T_8465 = {_T_8447,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@51668.4]
  assign _T_8467 = {_T_8448,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@51670.4]
  assign _T_8469 = {_T_8449,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@51672.4]
  assign _T_8471 = {_T_8450,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@51674.4]
  assign _T_8473 = {_T_8451,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@51676.4]
  assign _T_8475 = {_T_8452,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@51678.4]
  assign _T_8477 = {_T_8453,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@51680.4]
  assign _T_8479 = {_T_8454,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@51682.4]
  assign _T_8481 = {_T_8455,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@51684.4]
  assign _T_8483 = {_T_8456,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@51686.4]
  assign _T_8485 = {_T_8457,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@51688.4]
  assign _T_8487 = {_T_8458,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@51690.4]
  assign _T_8489 = {_T_8459,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@51692.4]
  assign _T_8490 = _T_8458 ? _T_8487 : _T_8489; // @[Mux.scala 31:69:@51693.4]
  assign _T_8491 = _T_8457 ? _T_8485 : _T_8490; // @[Mux.scala 31:69:@51694.4]
  assign _T_8492 = _T_8456 ? _T_8483 : _T_8491; // @[Mux.scala 31:69:@51695.4]
  assign _T_8493 = _T_8455 ? _T_8481 : _T_8492; // @[Mux.scala 31:69:@51696.4]
  assign _T_8494 = _T_8454 ? _T_8479 : _T_8493; // @[Mux.scala 31:69:@51697.4]
  assign _T_8495 = _T_8453 ? _T_8477 : _T_8494; // @[Mux.scala 31:69:@51698.4]
  assign _T_8496 = _T_8452 ? _T_8475 : _T_8495; // @[Mux.scala 31:69:@51699.4]
  assign _T_8497 = _T_8451 ? _T_8473 : _T_8496; // @[Mux.scala 31:69:@51700.4]
  assign _T_8498 = _T_8450 ? _T_8471 : _T_8497; // @[Mux.scala 31:69:@51701.4]
  assign _T_8499 = _T_8449 ? _T_8469 : _T_8498; // @[Mux.scala 31:69:@51702.4]
  assign _T_8500 = _T_8448 ? _T_8467 : _T_8499; // @[Mux.scala 31:69:@51703.4]
  assign _T_8501 = _T_8447 ? _T_8465 : _T_8500; // @[Mux.scala 31:69:@51704.4]
  assign _T_8502 = _T_8446 ? _T_8463 : _T_8501; // @[Mux.scala 31:69:@51705.4]
  assign _T_8503 = _T_8445 ? _T_8461 : _T_8502; // @[Mux.scala 31:69:@51706.4]
  assign _T_8511 = _T_7292 & _T_3950; // @[MemPrimitives.scala 110:228:@51715.4]
  assign _T_8517 = _T_7298 & _T_3956; // @[MemPrimitives.scala 110:228:@51719.4]
  assign _T_8523 = _T_7304 & _T_3962; // @[MemPrimitives.scala 110:228:@51723.4]
  assign _T_8529 = _T_7310 & _T_3968; // @[MemPrimitives.scala 110:228:@51727.4]
  assign _T_8535 = _T_7316 & _T_3974; // @[MemPrimitives.scala 110:228:@51731.4]
  assign _T_8541 = _T_7322 & _T_3980; // @[MemPrimitives.scala 110:228:@51735.4]
  assign _T_8547 = _T_7328 & _T_3986; // @[MemPrimitives.scala 110:228:@51739.4]
  assign _T_8553 = _T_7334 & _T_3992; // @[MemPrimitives.scala 110:228:@51743.4]
  assign _T_8559 = _T_7340 & _T_3998; // @[MemPrimitives.scala 110:228:@51747.4]
  assign _T_8565 = _T_7346 & _T_4004; // @[MemPrimitives.scala 110:228:@51751.4]
  assign _T_8571 = _T_7352 & _T_4010; // @[MemPrimitives.scala 110:228:@51755.4]
  assign _T_8577 = _T_7358 & _T_4016; // @[MemPrimitives.scala 110:228:@51759.4]
  assign _T_8583 = _T_7364 & _T_4022; // @[MemPrimitives.scala 110:228:@51763.4]
  assign _T_8589 = _T_7370 & _T_4028; // @[MemPrimitives.scala 110:228:@51767.4]
  assign _T_8595 = _T_7376 & _T_4034; // @[MemPrimitives.scala 110:228:@51771.4]
  assign _T_8597 = StickySelects_38_io_outs_0; // @[MemPrimitives.scala 123:41:@51791.4]
  assign _T_8598 = StickySelects_38_io_outs_1; // @[MemPrimitives.scala 123:41:@51792.4]
  assign _T_8599 = StickySelects_38_io_outs_2; // @[MemPrimitives.scala 123:41:@51793.4]
  assign _T_8600 = StickySelects_38_io_outs_3; // @[MemPrimitives.scala 123:41:@51794.4]
  assign _T_8601 = StickySelects_38_io_outs_4; // @[MemPrimitives.scala 123:41:@51795.4]
  assign _T_8602 = StickySelects_38_io_outs_5; // @[MemPrimitives.scala 123:41:@51796.4]
  assign _T_8603 = StickySelects_38_io_outs_6; // @[MemPrimitives.scala 123:41:@51797.4]
  assign _T_8604 = StickySelects_38_io_outs_7; // @[MemPrimitives.scala 123:41:@51798.4]
  assign _T_8605 = StickySelects_38_io_outs_8; // @[MemPrimitives.scala 123:41:@51799.4]
  assign _T_8606 = StickySelects_38_io_outs_9; // @[MemPrimitives.scala 123:41:@51800.4]
  assign _T_8607 = StickySelects_38_io_outs_10; // @[MemPrimitives.scala 123:41:@51801.4]
  assign _T_8608 = StickySelects_38_io_outs_11; // @[MemPrimitives.scala 123:41:@51802.4]
  assign _T_8609 = StickySelects_38_io_outs_12; // @[MemPrimitives.scala 123:41:@51803.4]
  assign _T_8610 = StickySelects_38_io_outs_13; // @[MemPrimitives.scala 123:41:@51804.4]
  assign _T_8611 = StickySelects_38_io_outs_14; // @[MemPrimitives.scala 123:41:@51805.4]
  assign _T_8613 = {_T_8597,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@51807.4]
  assign _T_8615 = {_T_8598,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@51809.4]
  assign _T_8617 = {_T_8599,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@51811.4]
  assign _T_8619 = {_T_8600,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@51813.4]
  assign _T_8621 = {_T_8601,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@51815.4]
  assign _T_8623 = {_T_8602,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@51817.4]
  assign _T_8625 = {_T_8603,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@51819.4]
  assign _T_8627 = {_T_8604,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@51821.4]
  assign _T_8629 = {_T_8605,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@51823.4]
  assign _T_8631 = {_T_8606,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@51825.4]
  assign _T_8633 = {_T_8607,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@51827.4]
  assign _T_8635 = {_T_8608,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@51829.4]
  assign _T_8637 = {_T_8609,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@51831.4]
  assign _T_8639 = {_T_8610,io_rPort_26_backpressure,io_rPort_26_ofs_0}; // @[Cat.scala 30:58:@51833.4]
  assign _T_8641 = {_T_8611,io_rPort_29_backpressure,io_rPort_29_ofs_0}; // @[Cat.scala 30:58:@51835.4]
  assign _T_8642 = _T_8610 ? _T_8639 : _T_8641; // @[Mux.scala 31:69:@51836.4]
  assign _T_8643 = _T_8609 ? _T_8637 : _T_8642; // @[Mux.scala 31:69:@51837.4]
  assign _T_8644 = _T_8608 ? _T_8635 : _T_8643; // @[Mux.scala 31:69:@51838.4]
  assign _T_8645 = _T_8607 ? _T_8633 : _T_8644; // @[Mux.scala 31:69:@51839.4]
  assign _T_8646 = _T_8606 ? _T_8631 : _T_8645; // @[Mux.scala 31:69:@51840.4]
  assign _T_8647 = _T_8605 ? _T_8629 : _T_8646; // @[Mux.scala 31:69:@51841.4]
  assign _T_8648 = _T_8604 ? _T_8627 : _T_8647; // @[Mux.scala 31:69:@51842.4]
  assign _T_8649 = _T_8603 ? _T_8625 : _T_8648; // @[Mux.scala 31:69:@51843.4]
  assign _T_8650 = _T_8602 ? _T_8623 : _T_8649; // @[Mux.scala 31:69:@51844.4]
  assign _T_8651 = _T_8601 ? _T_8621 : _T_8650; // @[Mux.scala 31:69:@51845.4]
  assign _T_8652 = _T_8600 ? _T_8619 : _T_8651; // @[Mux.scala 31:69:@51846.4]
  assign _T_8653 = _T_8599 ? _T_8617 : _T_8652; // @[Mux.scala 31:69:@51847.4]
  assign _T_8654 = _T_8598 ? _T_8615 : _T_8653; // @[Mux.scala 31:69:@51848.4]
  assign _T_8655 = _T_8597 ? _T_8613 : _T_8654; // @[Mux.scala 31:69:@51849.4]
  assign _T_8663 = _T_7444 & _T_4102; // @[MemPrimitives.scala 110:228:@51858.4]
  assign _T_8669 = _T_7450 & _T_4108; // @[MemPrimitives.scala 110:228:@51862.4]
  assign _T_8675 = _T_7456 & _T_4114; // @[MemPrimitives.scala 110:228:@51866.4]
  assign _T_8681 = _T_7462 & _T_4120; // @[MemPrimitives.scala 110:228:@51870.4]
  assign _T_8687 = _T_7468 & _T_4126; // @[MemPrimitives.scala 110:228:@51874.4]
  assign _T_8693 = _T_7474 & _T_4132; // @[MemPrimitives.scala 110:228:@51878.4]
  assign _T_8699 = _T_7480 & _T_4138; // @[MemPrimitives.scala 110:228:@51882.4]
  assign _T_8705 = _T_7486 & _T_4144; // @[MemPrimitives.scala 110:228:@51886.4]
  assign _T_8711 = _T_7492 & _T_4150; // @[MemPrimitives.scala 110:228:@51890.4]
  assign _T_8717 = _T_7498 & _T_4156; // @[MemPrimitives.scala 110:228:@51894.4]
  assign _T_8723 = _T_7504 & _T_4162; // @[MemPrimitives.scala 110:228:@51898.4]
  assign _T_8729 = _T_7510 & _T_4168; // @[MemPrimitives.scala 110:228:@51902.4]
  assign _T_8735 = _T_7516 & _T_4174; // @[MemPrimitives.scala 110:228:@51906.4]
  assign _T_8741 = _T_7522 & _T_4180; // @[MemPrimitives.scala 110:228:@51910.4]
  assign _T_8747 = _T_7528 & _T_4186; // @[MemPrimitives.scala 110:228:@51914.4]
  assign _T_8749 = StickySelects_39_io_outs_0; // @[MemPrimitives.scala 123:41:@51934.4]
  assign _T_8750 = StickySelects_39_io_outs_1; // @[MemPrimitives.scala 123:41:@51935.4]
  assign _T_8751 = StickySelects_39_io_outs_2; // @[MemPrimitives.scala 123:41:@51936.4]
  assign _T_8752 = StickySelects_39_io_outs_3; // @[MemPrimitives.scala 123:41:@51937.4]
  assign _T_8753 = StickySelects_39_io_outs_4; // @[MemPrimitives.scala 123:41:@51938.4]
  assign _T_8754 = StickySelects_39_io_outs_5; // @[MemPrimitives.scala 123:41:@51939.4]
  assign _T_8755 = StickySelects_39_io_outs_6; // @[MemPrimitives.scala 123:41:@51940.4]
  assign _T_8756 = StickySelects_39_io_outs_7; // @[MemPrimitives.scala 123:41:@51941.4]
  assign _T_8757 = StickySelects_39_io_outs_8; // @[MemPrimitives.scala 123:41:@51942.4]
  assign _T_8758 = StickySelects_39_io_outs_9; // @[MemPrimitives.scala 123:41:@51943.4]
  assign _T_8759 = StickySelects_39_io_outs_10; // @[MemPrimitives.scala 123:41:@51944.4]
  assign _T_8760 = StickySelects_39_io_outs_11; // @[MemPrimitives.scala 123:41:@51945.4]
  assign _T_8761 = StickySelects_39_io_outs_12; // @[MemPrimitives.scala 123:41:@51946.4]
  assign _T_8762 = StickySelects_39_io_outs_13; // @[MemPrimitives.scala 123:41:@51947.4]
  assign _T_8763 = StickySelects_39_io_outs_14; // @[MemPrimitives.scala 123:41:@51948.4]
  assign _T_8765 = {_T_8749,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@51950.4]
  assign _T_8767 = {_T_8750,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@51952.4]
  assign _T_8769 = {_T_8751,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@51954.4]
  assign _T_8771 = {_T_8752,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@51956.4]
  assign _T_8773 = {_T_8753,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@51958.4]
  assign _T_8775 = {_T_8754,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@51960.4]
  assign _T_8777 = {_T_8755,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@51962.4]
  assign _T_8779 = {_T_8756,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@51964.4]
  assign _T_8781 = {_T_8757,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@51966.4]
  assign _T_8783 = {_T_8758,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@51968.4]
  assign _T_8785 = {_T_8759,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@51970.4]
  assign _T_8787 = {_T_8760,io_rPort_24_backpressure,io_rPort_24_ofs_0}; // @[Cat.scala 30:58:@51972.4]
  assign _T_8789 = {_T_8761,io_rPort_25_backpressure,io_rPort_25_ofs_0}; // @[Cat.scala 30:58:@51974.4]
  assign _T_8791 = {_T_8762,io_rPort_27_backpressure,io_rPort_27_ofs_0}; // @[Cat.scala 30:58:@51976.4]
  assign _T_8793 = {_T_8763,io_rPort_28_backpressure,io_rPort_28_ofs_0}; // @[Cat.scala 30:58:@51978.4]
  assign _T_8794 = _T_8762 ? _T_8791 : _T_8793; // @[Mux.scala 31:69:@51979.4]
  assign _T_8795 = _T_8761 ? _T_8789 : _T_8794; // @[Mux.scala 31:69:@51980.4]
  assign _T_8796 = _T_8760 ? _T_8787 : _T_8795; // @[Mux.scala 31:69:@51981.4]
  assign _T_8797 = _T_8759 ? _T_8785 : _T_8796; // @[Mux.scala 31:69:@51982.4]
  assign _T_8798 = _T_8758 ? _T_8783 : _T_8797; // @[Mux.scala 31:69:@51983.4]
  assign _T_8799 = _T_8757 ? _T_8781 : _T_8798; // @[Mux.scala 31:69:@51984.4]
  assign _T_8800 = _T_8756 ? _T_8779 : _T_8799; // @[Mux.scala 31:69:@51985.4]
  assign _T_8801 = _T_8755 ? _T_8777 : _T_8800; // @[Mux.scala 31:69:@51986.4]
  assign _T_8802 = _T_8754 ? _T_8775 : _T_8801; // @[Mux.scala 31:69:@51987.4]
  assign _T_8803 = _T_8753 ? _T_8773 : _T_8802; // @[Mux.scala 31:69:@51988.4]
  assign _T_8804 = _T_8752 ? _T_8771 : _T_8803; // @[Mux.scala 31:69:@51989.4]
  assign _T_8805 = _T_8751 ? _T_8769 : _T_8804; // @[Mux.scala 31:69:@51990.4]
  assign _T_8806 = _T_8750 ? _T_8767 : _T_8805; // @[Mux.scala 31:69:@51991.4]
  assign _T_8807 = _T_8749 ? _T_8765 : _T_8806; // @[Mux.scala 31:69:@51992.4]
  assign _T_8967 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@52209.4 package.scala 96:25:@52210.4]
  assign _T_8971 = _T_8967 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@52219.4]
  assign _T_8964 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@52201.4 package.scala 96:25:@52202.4]
  assign _T_8972 = _T_8964 ? Mem1D_34_io_output : _T_8971; // @[Mux.scala 31:69:@52220.4]
  assign _T_8961 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@52193.4 package.scala 96:25:@52194.4]
  assign _T_8973 = _T_8961 ? Mem1D_32_io_output : _T_8972; // @[Mux.scala 31:69:@52221.4]
  assign _T_8958 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@52185.4 package.scala 96:25:@52186.4]
  assign _T_8974 = _T_8958 ? Mem1D_30_io_output : _T_8973; // @[Mux.scala 31:69:@52222.4]
  assign _T_8955 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@52177.4 package.scala 96:25:@52178.4]
  assign _T_8975 = _T_8955 ? Mem1D_28_io_output : _T_8974; // @[Mux.scala 31:69:@52223.4]
  assign _T_8952 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@52169.4 package.scala 96:25:@52170.4]
  assign _T_8976 = _T_8952 ? Mem1D_26_io_output : _T_8975; // @[Mux.scala 31:69:@52224.4]
  assign _T_8949 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@52161.4 package.scala 96:25:@52162.4]
  assign _T_8977 = _T_8949 ? Mem1D_24_io_output : _T_8976; // @[Mux.scala 31:69:@52225.4]
  assign _T_8946 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@52153.4 package.scala 96:25:@52154.4]
  assign _T_8978 = _T_8946 ? Mem1D_22_io_output : _T_8977; // @[Mux.scala 31:69:@52226.4]
  assign _T_8943 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@52145.4 package.scala 96:25:@52146.4]
  assign _T_8979 = _T_8943 ? Mem1D_20_io_output : _T_8978; // @[Mux.scala 31:69:@52227.4]
  assign _T_8940 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@52137.4 package.scala 96:25:@52138.4]
  assign _T_8980 = _T_8940 ? Mem1D_18_io_output : _T_8979; // @[Mux.scala 31:69:@52228.4]
  assign _T_8937 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@52129.4 package.scala 96:25:@52130.4]
  assign _T_8981 = _T_8937 ? Mem1D_16_io_output : _T_8980; // @[Mux.scala 31:69:@52229.4]
  assign _T_8934 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@52121.4 package.scala 96:25:@52122.4]
  assign _T_8982 = _T_8934 ? Mem1D_14_io_output : _T_8981; // @[Mux.scala 31:69:@52230.4]
  assign _T_8931 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@52113.4 package.scala 96:25:@52114.4]
  assign _T_8983 = _T_8931 ? Mem1D_12_io_output : _T_8982; // @[Mux.scala 31:69:@52231.4]
  assign _T_8928 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@52105.4 package.scala 96:25:@52106.4]
  assign _T_8984 = _T_8928 ? Mem1D_10_io_output : _T_8983; // @[Mux.scala 31:69:@52232.4]
  assign _T_8925 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@52097.4 package.scala 96:25:@52098.4]
  assign _T_8985 = _T_8925 ? Mem1D_8_io_output : _T_8984; // @[Mux.scala 31:69:@52233.4]
  assign _T_8922 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@52089.4 package.scala 96:25:@52090.4]
  assign _T_8986 = _T_8922 ? Mem1D_6_io_output : _T_8985; // @[Mux.scala 31:69:@52234.4]
  assign _T_8919 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@52081.4 package.scala 96:25:@52082.4]
  assign _T_8987 = _T_8919 ? Mem1D_4_io_output : _T_8986; // @[Mux.scala 31:69:@52235.4]
  assign _T_8916 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@52073.4 package.scala 96:25:@52074.4]
  assign _T_8988 = _T_8916 ? Mem1D_2_io_output : _T_8987; // @[Mux.scala 31:69:@52236.4]
  assign _T_8913 = RetimeWrapper_io_out; // @[package.scala 96:25:@52065.4 package.scala 96:25:@52066.4]
  assign _T_9146 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@52449.4 package.scala 96:25:@52450.4]
  assign _T_9150 = _T_9146 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@52459.4]
  assign _T_9143 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@52441.4 package.scala 96:25:@52442.4]
  assign _T_9151 = _T_9143 ? Mem1D_34_io_output : _T_9150; // @[Mux.scala 31:69:@52460.4]
  assign _T_9140 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@52433.4 package.scala 96:25:@52434.4]
  assign _T_9152 = _T_9140 ? Mem1D_32_io_output : _T_9151; // @[Mux.scala 31:69:@52461.4]
  assign _T_9137 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@52425.4 package.scala 96:25:@52426.4]
  assign _T_9153 = _T_9137 ? Mem1D_30_io_output : _T_9152; // @[Mux.scala 31:69:@52462.4]
  assign _T_9134 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@52417.4 package.scala 96:25:@52418.4]
  assign _T_9154 = _T_9134 ? Mem1D_28_io_output : _T_9153; // @[Mux.scala 31:69:@52463.4]
  assign _T_9131 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@52409.4 package.scala 96:25:@52410.4]
  assign _T_9155 = _T_9131 ? Mem1D_26_io_output : _T_9154; // @[Mux.scala 31:69:@52464.4]
  assign _T_9128 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@52401.4 package.scala 96:25:@52402.4]
  assign _T_9156 = _T_9128 ? Mem1D_24_io_output : _T_9155; // @[Mux.scala 31:69:@52465.4]
  assign _T_9125 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@52393.4 package.scala 96:25:@52394.4]
  assign _T_9157 = _T_9125 ? Mem1D_22_io_output : _T_9156; // @[Mux.scala 31:69:@52466.4]
  assign _T_9122 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@52385.4 package.scala 96:25:@52386.4]
  assign _T_9158 = _T_9122 ? Mem1D_20_io_output : _T_9157; // @[Mux.scala 31:69:@52467.4]
  assign _T_9119 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@52377.4 package.scala 96:25:@52378.4]
  assign _T_9159 = _T_9119 ? Mem1D_18_io_output : _T_9158; // @[Mux.scala 31:69:@52468.4]
  assign _T_9116 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@52369.4 package.scala 96:25:@52370.4]
  assign _T_9160 = _T_9116 ? Mem1D_16_io_output : _T_9159; // @[Mux.scala 31:69:@52469.4]
  assign _T_9113 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@52361.4 package.scala 96:25:@52362.4]
  assign _T_9161 = _T_9113 ? Mem1D_14_io_output : _T_9160; // @[Mux.scala 31:69:@52470.4]
  assign _T_9110 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@52353.4 package.scala 96:25:@52354.4]
  assign _T_9162 = _T_9110 ? Mem1D_12_io_output : _T_9161; // @[Mux.scala 31:69:@52471.4]
  assign _T_9107 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@52345.4 package.scala 96:25:@52346.4]
  assign _T_9163 = _T_9107 ? Mem1D_10_io_output : _T_9162; // @[Mux.scala 31:69:@52472.4]
  assign _T_9104 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@52337.4 package.scala 96:25:@52338.4]
  assign _T_9164 = _T_9104 ? Mem1D_8_io_output : _T_9163; // @[Mux.scala 31:69:@52473.4]
  assign _T_9101 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@52329.4 package.scala 96:25:@52330.4]
  assign _T_9165 = _T_9101 ? Mem1D_6_io_output : _T_9164; // @[Mux.scala 31:69:@52474.4]
  assign _T_9098 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@52321.4 package.scala 96:25:@52322.4]
  assign _T_9166 = _T_9098 ? Mem1D_4_io_output : _T_9165; // @[Mux.scala 31:69:@52475.4]
  assign _T_9095 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@52313.4 package.scala 96:25:@52314.4]
  assign _T_9167 = _T_9095 ? Mem1D_2_io_output : _T_9166; // @[Mux.scala 31:69:@52476.4]
  assign _T_9092 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@52305.4 package.scala 96:25:@52306.4]
  assign _T_9325 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@52689.4 package.scala 96:25:@52690.4]
  assign _T_9329 = _T_9325 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@52699.4]
  assign _T_9322 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@52681.4 package.scala 96:25:@52682.4]
  assign _T_9330 = _T_9322 ? Mem1D_35_io_output : _T_9329; // @[Mux.scala 31:69:@52700.4]
  assign _T_9319 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@52673.4 package.scala 96:25:@52674.4]
  assign _T_9331 = _T_9319 ? Mem1D_33_io_output : _T_9330; // @[Mux.scala 31:69:@52701.4]
  assign _T_9316 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@52665.4 package.scala 96:25:@52666.4]
  assign _T_9332 = _T_9316 ? Mem1D_31_io_output : _T_9331; // @[Mux.scala 31:69:@52702.4]
  assign _T_9313 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@52657.4 package.scala 96:25:@52658.4]
  assign _T_9333 = _T_9313 ? Mem1D_29_io_output : _T_9332; // @[Mux.scala 31:69:@52703.4]
  assign _T_9310 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@52649.4 package.scala 96:25:@52650.4]
  assign _T_9334 = _T_9310 ? Mem1D_27_io_output : _T_9333; // @[Mux.scala 31:69:@52704.4]
  assign _T_9307 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@52641.4 package.scala 96:25:@52642.4]
  assign _T_9335 = _T_9307 ? Mem1D_25_io_output : _T_9334; // @[Mux.scala 31:69:@52705.4]
  assign _T_9304 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@52633.4 package.scala 96:25:@52634.4]
  assign _T_9336 = _T_9304 ? Mem1D_23_io_output : _T_9335; // @[Mux.scala 31:69:@52706.4]
  assign _T_9301 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@52625.4 package.scala 96:25:@52626.4]
  assign _T_9337 = _T_9301 ? Mem1D_21_io_output : _T_9336; // @[Mux.scala 31:69:@52707.4]
  assign _T_9298 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@52617.4 package.scala 96:25:@52618.4]
  assign _T_9338 = _T_9298 ? Mem1D_19_io_output : _T_9337; // @[Mux.scala 31:69:@52708.4]
  assign _T_9295 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@52609.4 package.scala 96:25:@52610.4]
  assign _T_9339 = _T_9295 ? Mem1D_17_io_output : _T_9338; // @[Mux.scala 31:69:@52709.4]
  assign _T_9292 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@52601.4 package.scala 96:25:@52602.4]
  assign _T_9340 = _T_9292 ? Mem1D_15_io_output : _T_9339; // @[Mux.scala 31:69:@52710.4]
  assign _T_9289 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@52593.4 package.scala 96:25:@52594.4]
  assign _T_9341 = _T_9289 ? Mem1D_13_io_output : _T_9340; // @[Mux.scala 31:69:@52711.4]
  assign _T_9286 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@52585.4 package.scala 96:25:@52586.4]
  assign _T_9342 = _T_9286 ? Mem1D_11_io_output : _T_9341; // @[Mux.scala 31:69:@52712.4]
  assign _T_9283 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@52577.4 package.scala 96:25:@52578.4]
  assign _T_9343 = _T_9283 ? Mem1D_9_io_output : _T_9342; // @[Mux.scala 31:69:@52713.4]
  assign _T_9280 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@52569.4 package.scala 96:25:@52570.4]
  assign _T_9344 = _T_9280 ? Mem1D_7_io_output : _T_9343; // @[Mux.scala 31:69:@52714.4]
  assign _T_9277 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@52561.4 package.scala 96:25:@52562.4]
  assign _T_9345 = _T_9277 ? Mem1D_5_io_output : _T_9344; // @[Mux.scala 31:69:@52715.4]
  assign _T_9274 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@52553.4 package.scala 96:25:@52554.4]
  assign _T_9346 = _T_9274 ? Mem1D_3_io_output : _T_9345; // @[Mux.scala 31:69:@52716.4]
  assign _T_9271 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@52545.4 package.scala 96:25:@52546.4]
  assign _T_9504 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@52929.4 package.scala 96:25:@52930.4]
  assign _T_9508 = _T_9504 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@52939.4]
  assign _T_9501 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@52921.4 package.scala 96:25:@52922.4]
  assign _T_9509 = _T_9501 ? Mem1D_34_io_output : _T_9508; // @[Mux.scala 31:69:@52940.4]
  assign _T_9498 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@52913.4 package.scala 96:25:@52914.4]
  assign _T_9510 = _T_9498 ? Mem1D_32_io_output : _T_9509; // @[Mux.scala 31:69:@52941.4]
  assign _T_9495 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@52905.4 package.scala 96:25:@52906.4]
  assign _T_9511 = _T_9495 ? Mem1D_30_io_output : _T_9510; // @[Mux.scala 31:69:@52942.4]
  assign _T_9492 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@52897.4 package.scala 96:25:@52898.4]
  assign _T_9512 = _T_9492 ? Mem1D_28_io_output : _T_9511; // @[Mux.scala 31:69:@52943.4]
  assign _T_9489 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@52889.4 package.scala 96:25:@52890.4]
  assign _T_9513 = _T_9489 ? Mem1D_26_io_output : _T_9512; // @[Mux.scala 31:69:@52944.4]
  assign _T_9486 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@52881.4 package.scala 96:25:@52882.4]
  assign _T_9514 = _T_9486 ? Mem1D_24_io_output : _T_9513; // @[Mux.scala 31:69:@52945.4]
  assign _T_9483 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@52873.4 package.scala 96:25:@52874.4]
  assign _T_9515 = _T_9483 ? Mem1D_22_io_output : _T_9514; // @[Mux.scala 31:69:@52946.4]
  assign _T_9480 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@52865.4 package.scala 96:25:@52866.4]
  assign _T_9516 = _T_9480 ? Mem1D_20_io_output : _T_9515; // @[Mux.scala 31:69:@52947.4]
  assign _T_9477 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@52857.4 package.scala 96:25:@52858.4]
  assign _T_9517 = _T_9477 ? Mem1D_18_io_output : _T_9516; // @[Mux.scala 31:69:@52948.4]
  assign _T_9474 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@52849.4 package.scala 96:25:@52850.4]
  assign _T_9518 = _T_9474 ? Mem1D_16_io_output : _T_9517; // @[Mux.scala 31:69:@52949.4]
  assign _T_9471 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@52841.4 package.scala 96:25:@52842.4]
  assign _T_9519 = _T_9471 ? Mem1D_14_io_output : _T_9518; // @[Mux.scala 31:69:@52950.4]
  assign _T_9468 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@52833.4 package.scala 96:25:@52834.4]
  assign _T_9520 = _T_9468 ? Mem1D_12_io_output : _T_9519; // @[Mux.scala 31:69:@52951.4]
  assign _T_9465 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@52825.4 package.scala 96:25:@52826.4]
  assign _T_9521 = _T_9465 ? Mem1D_10_io_output : _T_9520; // @[Mux.scala 31:69:@52952.4]
  assign _T_9462 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@52817.4 package.scala 96:25:@52818.4]
  assign _T_9522 = _T_9462 ? Mem1D_8_io_output : _T_9521; // @[Mux.scala 31:69:@52953.4]
  assign _T_9459 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@52809.4 package.scala 96:25:@52810.4]
  assign _T_9523 = _T_9459 ? Mem1D_6_io_output : _T_9522; // @[Mux.scala 31:69:@52954.4]
  assign _T_9456 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@52801.4 package.scala 96:25:@52802.4]
  assign _T_9524 = _T_9456 ? Mem1D_4_io_output : _T_9523; // @[Mux.scala 31:69:@52955.4]
  assign _T_9453 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@52793.4 package.scala 96:25:@52794.4]
  assign _T_9525 = _T_9453 ? Mem1D_2_io_output : _T_9524; // @[Mux.scala 31:69:@52956.4]
  assign _T_9450 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@52785.4 package.scala 96:25:@52786.4]
  assign _T_9683 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@53169.4 package.scala 96:25:@53170.4]
  assign _T_9687 = _T_9683 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@53179.4]
  assign _T_9680 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@53161.4 package.scala 96:25:@53162.4]
  assign _T_9688 = _T_9680 ? Mem1D_34_io_output : _T_9687; // @[Mux.scala 31:69:@53180.4]
  assign _T_9677 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@53153.4 package.scala 96:25:@53154.4]
  assign _T_9689 = _T_9677 ? Mem1D_32_io_output : _T_9688; // @[Mux.scala 31:69:@53181.4]
  assign _T_9674 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@53145.4 package.scala 96:25:@53146.4]
  assign _T_9690 = _T_9674 ? Mem1D_30_io_output : _T_9689; // @[Mux.scala 31:69:@53182.4]
  assign _T_9671 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@53137.4 package.scala 96:25:@53138.4]
  assign _T_9691 = _T_9671 ? Mem1D_28_io_output : _T_9690; // @[Mux.scala 31:69:@53183.4]
  assign _T_9668 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@53129.4 package.scala 96:25:@53130.4]
  assign _T_9692 = _T_9668 ? Mem1D_26_io_output : _T_9691; // @[Mux.scala 31:69:@53184.4]
  assign _T_9665 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@53121.4 package.scala 96:25:@53122.4]
  assign _T_9693 = _T_9665 ? Mem1D_24_io_output : _T_9692; // @[Mux.scala 31:69:@53185.4]
  assign _T_9662 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@53113.4 package.scala 96:25:@53114.4]
  assign _T_9694 = _T_9662 ? Mem1D_22_io_output : _T_9693; // @[Mux.scala 31:69:@53186.4]
  assign _T_9659 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@53105.4 package.scala 96:25:@53106.4]
  assign _T_9695 = _T_9659 ? Mem1D_20_io_output : _T_9694; // @[Mux.scala 31:69:@53187.4]
  assign _T_9656 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@53097.4 package.scala 96:25:@53098.4]
  assign _T_9696 = _T_9656 ? Mem1D_18_io_output : _T_9695; // @[Mux.scala 31:69:@53188.4]
  assign _T_9653 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@53089.4 package.scala 96:25:@53090.4]
  assign _T_9697 = _T_9653 ? Mem1D_16_io_output : _T_9696; // @[Mux.scala 31:69:@53189.4]
  assign _T_9650 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@53081.4 package.scala 96:25:@53082.4]
  assign _T_9698 = _T_9650 ? Mem1D_14_io_output : _T_9697; // @[Mux.scala 31:69:@53190.4]
  assign _T_9647 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@53073.4 package.scala 96:25:@53074.4]
  assign _T_9699 = _T_9647 ? Mem1D_12_io_output : _T_9698; // @[Mux.scala 31:69:@53191.4]
  assign _T_9644 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@53065.4 package.scala 96:25:@53066.4]
  assign _T_9700 = _T_9644 ? Mem1D_10_io_output : _T_9699; // @[Mux.scala 31:69:@53192.4]
  assign _T_9641 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@53057.4 package.scala 96:25:@53058.4]
  assign _T_9701 = _T_9641 ? Mem1D_8_io_output : _T_9700; // @[Mux.scala 31:69:@53193.4]
  assign _T_9638 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@53049.4 package.scala 96:25:@53050.4]
  assign _T_9702 = _T_9638 ? Mem1D_6_io_output : _T_9701; // @[Mux.scala 31:69:@53194.4]
  assign _T_9635 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@53041.4 package.scala 96:25:@53042.4]
  assign _T_9703 = _T_9635 ? Mem1D_4_io_output : _T_9702; // @[Mux.scala 31:69:@53195.4]
  assign _T_9632 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@53033.4 package.scala 96:25:@53034.4]
  assign _T_9704 = _T_9632 ? Mem1D_2_io_output : _T_9703; // @[Mux.scala 31:69:@53196.4]
  assign _T_9629 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@53025.4 package.scala 96:25:@53026.4]
  assign _T_9862 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@53409.4 package.scala 96:25:@53410.4]
  assign _T_9866 = _T_9862 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@53419.4]
  assign _T_9859 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@53401.4 package.scala 96:25:@53402.4]
  assign _T_9867 = _T_9859 ? Mem1D_34_io_output : _T_9866; // @[Mux.scala 31:69:@53420.4]
  assign _T_9856 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@53393.4 package.scala 96:25:@53394.4]
  assign _T_9868 = _T_9856 ? Mem1D_32_io_output : _T_9867; // @[Mux.scala 31:69:@53421.4]
  assign _T_9853 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@53385.4 package.scala 96:25:@53386.4]
  assign _T_9869 = _T_9853 ? Mem1D_30_io_output : _T_9868; // @[Mux.scala 31:69:@53422.4]
  assign _T_9850 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@53377.4 package.scala 96:25:@53378.4]
  assign _T_9870 = _T_9850 ? Mem1D_28_io_output : _T_9869; // @[Mux.scala 31:69:@53423.4]
  assign _T_9847 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@53369.4 package.scala 96:25:@53370.4]
  assign _T_9871 = _T_9847 ? Mem1D_26_io_output : _T_9870; // @[Mux.scala 31:69:@53424.4]
  assign _T_9844 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@53361.4 package.scala 96:25:@53362.4]
  assign _T_9872 = _T_9844 ? Mem1D_24_io_output : _T_9871; // @[Mux.scala 31:69:@53425.4]
  assign _T_9841 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@53353.4 package.scala 96:25:@53354.4]
  assign _T_9873 = _T_9841 ? Mem1D_22_io_output : _T_9872; // @[Mux.scala 31:69:@53426.4]
  assign _T_9838 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@53345.4 package.scala 96:25:@53346.4]
  assign _T_9874 = _T_9838 ? Mem1D_20_io_output : _T_9873; // @[Mux.scala 31:69:@53427.4]
  assign _T_9835 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@53337.4 package.scala 96:25:@53338.4]
  assign _T_9875 = _T_9835 ? Mem1D_18_io_output : _T_9874; // @[Mux.scala 31:69:@53428.4]
  assign _T_9832 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@53329.4 package.scala 96:25:@53330.4]
  assign _T_9876 = _T_9832 ? Mem1D_16_io_output : _T_9875; // @[Mux.scala 31:69:@53429.4]
  assign _T_9829 = RetimeWrapper_107_io_out; // @[package.scala 96:25:@53321.4 package.scala 96:25:@53322.4]
  assign _T_9877 = _T_9829 ? Mem1D_14_io_output : _T_9876; // @[Mux.scala 31:69:@53430.4]
  assign _T_9826 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@53313.4 package.scala 96:25:@53314.4]
  assign _T_9878 = _T_9826 ? Mem1D_12_io_output : _T_9877; // @[Mux.scala 31:69:@53431.4]
  assign _T_9823 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@53305.4 package.scala 96:25:@53306.4]
  assign _T_9879 = _T_9823 ? Mem1D_10_io_output : _T_9878; // @[Mux.scala 31:69:@53432.4]
  assign _T_9820 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@53297.4 package.scala 96:25:@53298.4]
  assign _T_9880 = _T_9820 ? Mem1D_8_io_output : _T_9879; // @[Mux.scala 31:69:@53433.4]
  assign _T_9817 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@53289.4 package.scala 96:25:@53290.4]
  assign _T_9881 = _T_9817 ? Mem1D_6_io_output : _T_9880; // @[Mux.scala 31:69:@53434.4]
  assign _T_9814 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@53281.4 package.scala 96:25:@53282.4]
  assign _T_9882 = _T_9814 ? Mem1D_4_io_output : _T_9881; // @[Mux.scala 31:69:@53435.4]
  assign _T_9811 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@53273.4 package.scala 96:25:@53274.4]
  assign _T_9883 = _T_9811 ? Mem1D_2_io_output : _T_9882; // @[Mux.scala 31:69:@53436.4]
  assign _T_9808 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@53265.4 package.scala 96:25:@53266.4]
  assign _T_10041 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@53649.4 package.scala 96:25:@53650.4]
  assign _T_10045 = _T_10041 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@53659.4]
  assign _T_10038 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@53641.4 package.scala 96:25:@53642.4]
  assign _T_10046 = _T_10038 ? Mem1D_35_io_output : _T_10045; // @[Mux.scala 31:69:@53660.4]
  assign _T_10035 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@53633.4 package.scala 96:25:@53634.4]
  assign _T_10047 = _T_10035 ? Mem1D_33_io_output : _T_10046; // @[Mux.scala 31:69:@53661.4]
  assign _T_10032 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@53625.4 package.scala 96:25:@53626.4]
  assign _T_10048 = _T_10032 ? Mem1D_31_io_output : _T_10047; // @[Mux.scala 31:69:@53662.4]
  assign _T_10029 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@53617.4 package.scala 96:25:@53618.4]
  assign _T_10049 = _T_10029 ? Mem1D_29_io_output : _T_10048; // @[Mux.scala 31:69:@53663.4]
  assign _T_10026 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@53609.4 package.scala 96:25:@53610.4]
  assign _T_10050 = _T_10026 ? Mem1D_27_io_output : _T_10049; // @[Mux.scala 31:69:@53664.4]
  assign _T_10023 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@53601.4 package.scala 96:25:@53602.4]
  assign _T_10051 = _T_10023 ? Mem1D_25_io_output : _T_10050; // @[Mux.scala 31:69:@53665.4]
  assign _T_10020 = RetimeWrapper_131_io_out; // @[package.scala 96:25:@53593.4 package.scala 96:25:@53594.4]
  assign _T_10052 = _T_10020 ? Mem1D_23_io_output : _T_10051; // @[Mux.scala 31:69:@53666.4]
  assign _T_10017 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@53585.4 package.scala 96:25:@53586.4]
  assign _T_10053 = _T_10017 ? Mem1D_21_io_output : _T_10052; // @[Mux.scala 31:69:@53667.4]
  assign _T_10014 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@53577.4 package.scala 96:25:@53578.4]
  assign _T_10054 = _T_10014 ? Mem1D_19_io_output : _T_10053; // @[Mux.scala 31:69:@53668.4]
  assign _T_10011 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@53569.4 package.scala 96:25:@53570.4]
  assign _T_10055 = _T_10011 ? Mem1D_17_io_output : _T_10054; // @[Mux.scala 31:69:@53669.4]
  assign _T_10008 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@53561.4 package.scala 96:25:@53562.4]
  assign _T_10056 = _T_10008 ? Mem1D_15_io_output : _T_10055; // @[Mux.scala 31:69:@53670.4]
  assign _T_10005 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@53553.4 package.scala 96:25:@53554.4]
  assign _T_10057 = _T_10005 ? Mem1D_13_io_output : _T_10056; // @[Mux.scala 31:69:@53671.4]
  assign _T_10002 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@53545.4 package.scala 96:25:@53546.4]
  assign _T_10058 = _T_10002 ? Mem1D_11_io_output : _T_10057; // @[Mux.scala 31:69:@53672.4]
  assign _T_9999 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@53537.4 package.scala 96:25:@53538.4]
  assign _T_10059 = _T_9999 ? Mem1D_9_io_output : _T_10058; // @[Mux.scala 31:69:@53673.4]
  assign _T_9996 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@53529.4 package.scala 96:25:@53530.4]
  assign _T_10060 = _T_9996 ? Mem1D_7_io_output : _T_10059; // @[Mux.scala 31:69:@53674.4]
  assign _T_9993 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@53521.4 package.scala 96:25:@53522.4]
  assign _T_10061 = _T_9993 ? Mem1D_5_io_output : _T_10060; // @[Mux.scala 31:69:@53675.4]
  assign _T_9990 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@53513.4 package.scala 96:25:@53514.4]
  assign _T_10062 = _T_9990 ? Mem1D_3_io_output : _T_10061; // @[Mux.scala 31:69:@53676.4]
  assign _T_9987 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@53505.4 package.scala 96:25:@53506.4]
  assign _T_10220 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@53889.4 package.scala 96:25:@53890.4]
  assign _T_10224 = _T_10220 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@53899.4]
  assign _T_10217 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@53881.4 package.scala 96:25:@53882.4]
  assign _T_10225 = _T_10217 ? Mem1D_35_io_output : _T_10224; // @[Mux.scala 31:69:@53900.4]
  assign _T_10214 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@53873.4 package.scala 96:25:@53874.4]
  assign _T_10226 = _T_10214 ? Mem1D_33_io_output : _T_10225; // @[Mux.scala 31:69:@53901.4]
  assign _T_10211 = RetimeWrapper_155_io_out; // @[package.scala 96:25:@53865.4 package.scala 96:25:@53866.4]
  assign _T_10227 = _T_10211 ? Mem1D_31_io_output : _T_10226; // @[Mux.scala 31:69:@53902.4]
  assign _T_10208 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@53857.4 package.scala 96:25:@53858.4]
  assign _T_10228 = _T_10208 ? Mem1D_29_io_output : _T_10227; // @[Mux.scala 31:69:@53903.4]
  assign _T_10205 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@53849.4 package.scala 96:25:@53850.4]
  assign _T_10229 = _T_10205 ? Mem1D_27_io_output : _T_10228; // @[Mux.scala 31:69:@53904.4]
  assign _T_10202 = RetimeWrapper_152_io_out; // @[package.scala 96:25:@53841.4 package.scala 96:25:@53842.4]
  assign _T_10230 = _T_10202 ? Mem1D_25_io_output : _T_10229; // @[Mux.scala 31:69:@53905.4]
  assign _T_10199 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@53833.4 package.scala 96:25:@53834.4]
  assign _T_10231 = _T_10199 ? Mem1D_23_io_output : _T_10230; // @[Mux.scala 31:69:@53906.4]
  assign _T_10196 = RetimeWrapper_150_io_out; // @[package.scala 96:25:@53825.4 package.scala 96:25:@53826.4]
  assign _T_10232 = _T_10196 ? Mem1D_21_io_output : _T_10231; // @[Mux.scala 31:69:@53907.4]
  assign _T_10193 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@53817.4 package.scala 96:25:@53818.4]
  assign _T_10233 = _T_10193 ? Mem1D_19_io_output : _T_10232; // @[Mux.scala 31:69:@53908.4]
  assign _T_10190 = RetimeWrapper_148_io_out; // @[package.scala 96:25:@53809.4 package.scala 96:25:@53810.4]
  assign _T_10234 = _T_10190 ? Mem1D_17_io_output : _T_10233; // @[Mux.scala 31:69:@53909.4]
  assign _T_10187 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@53801.4 package.scala 96:25:@53802.4]
  assign _T_10235 = _T_10187 ? Mem1D_15_io_output : _T_10234; // @[Mux.scala 31:69:@53910.4]
  assign _T_10184 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@53793.4 package.scala 96:25:@53794.4]
  assign _T_10236 = _T_10184 ? Mem1D_13_io_output : _T_10235; // @[Mux.scala 31:69:@53911.4]
  assign _T_10181 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@53785.4 package.scala 96:25:@53786.4]
  assign _T_10237 = _T_10181 ? Mem1D_11_io_output : _T_10236; // @[Mux.scala 31:69:@53912.4]
  assign _T_10178 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@53777.4 package.scala 96:25:@53778.4]
  assign _T_10238 = _T_10178 ? Mem1D_9_io_output : _T_10237; // @[Mux.scala 31:69:@53913.4]
  assign _T_10175 = RetimeWrapper_143_io_out; // @[package.scala 96:25:@53769.4 package.scala 96:25:@53770.4]
  assign _T_10239 = _T_10175 ? Mem1D_7_io_output : _T_10238; // @[Mux.scala 31:69:@53914.4]
  assign _T_10172 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@53761.4 package.scala 96:25:@53762.4]
  assign _T_10240 = _T_10172 ? Mem1D_5_io_output : _T_10239; // @[Mux.scala 31:69:@53915.4]
  assign _T_10169 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@53753.4 package.scala 96:25:@53754.4]
  assign _T_10241 = _T_10169 ? Mem1D_3_io_output : _T_10240; // @[Mux.scala 31:69:@53916.4]
  assign _T_10166 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@53745.4 package.scala 96:25:@53746.4]
  assign _T_10399 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@54129.4 package.scala 96:25:@54130.4]
  assign _T_10403 = _T_10399 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@54139.4]
  assign _T_10396 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@54121.4 package.scala 96:25:@54122.4]
  assign _T_10404 = _T_10396 ? Mem1D_35_io_output : _T_10403; // @[Mux.scala 31:69:@54140.4]
  assign _T_10393 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@54113.4 package.scala 96:25:@54114.4]
  assign _T_10405 = _T_10393 ? Mem1D_33_io_output : _T_10404; // @[Mux.scala 31:69:@54141.4]
  assign _T_10390 = RetimeWrapper_175_io_out; // @[package.scala 96:25:@54105.4 package.scala 96:25:@54106.4]
  assign _T_10406 = _T_10390 ? Mem1D_31_io_output : _T_10405; // @[Mux.scala 31:69:@54142.4]
  assign _T_10387 = RetimeWrapper_174_io_out; // @[package.scala 96:25:@54097.4 package.scala 96:25:@54098.4]
  assign _T_10407 = _T_10387 ? Mem1D_29_io_output : _T_10406; // @[Mux.scala 31:69:@54143.4]
  assign _T_10384 = RetimeWrapper_173_io_out; // @[package.scala 96:25:@54089.4 package.scala 96:25:@54090.4]
  assign _T_10408 = _T_10384 ? Mem1D_27_io_output : _T_10407; // @[Mux.scala 31:69:@54144.4]
  assign _T_10381 = RetimeWrapper_172_io_out; // @[package.scala 96:25:@54081.4 package.scala 96:25:@54082.4]
  assign _T_10409 = _T_10381 ? Mem1D_25_io_output : _T_10408; // @[Mux.scala 31:69:@54145.4]
  assign _T_10378 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@54073.4 package.scala 96:25:@54074.4]
  assign _T_10410 = _T_10378 ? Mem1D_23_io_output : _T_10409; // @[Mux.scala 31:69:@54146.4]
  assign _T_10375 = RetimeWrapper_170_io_out; // @[package.scala 96:25:@54065.4 package.scala 96:25:@54066.4]
  assign _T_10411 = _T_10375 ? Mem1D_21_io_output : _T_10410; // @[Mux.scala 31:69:@54147.4]
  assign _T_10372 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@54057.4 package.scala 96:25:@54058.4]
  assign _T_10412 = _T_10372 ? Mem1D_19_io_output : _T_10411; // @[Mux.scala 31:69:@54148.4]
  assign _T_10369 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@54049.4 package.scala 96:25:@54050.4]
  assign _T_10413 = _T_10369 ? Mem1D_17_io_output : _T_10412; // @[Mux.scala 31:69:@54149.4]
  assign _T_10366 = RetimeWrapper_167_io_out; // @[package.scala 96:25:@54041.4 package.scala 96:25:@54042.4]
  assign _T_10414 = _T_10366 ? Mem1D_15_io_output : _T_10413; // @[Mux.scala 31:69:@54150.4]
  assign _T_10363 = RetimeWrapper_166_io_out; // @[package.scala 96:25:@54033.4 package.scala 96:25:@54034.4]
  assign _T_10415 = _T_10363 ? Mem1D_13_io_output : _T_10414; // @[Mux.scala 31:69:@54151.4]
  assign _T_10360 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@54025.4 package.scala 96:25:@54026.4]
  assign _T_10416 = _T_10360 ? Mem1D_11_io_output : _T_10415; // @[Mux.scala 31:69:@54152.4]
  assign _T_10357 = RetimeWrapper_164_io_out; // @[package.scala 96:25:@54017.4 package.scala 96:25:@54018.4]
  assign _T_10417 = _T_10357 ? Mem1D_9_io_output : _T_10416; // @[Mux.scala 31:69:@54153.4]
  assign _T_10354 = RetimeWrapper_163_io_out; // @[package.scala 96:25:@54009.4 package.scala 96:25:@54010.4]
  assign _T_10418 = _T_10354 ? Mem1D_7_io_output : _T_10417; // @[Mux.scala 31:69:@54154.4]
  assign _T_10351 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@54001.4 package.scala 96:25:@54002.4]
  assign _T_10419 = _T_10351 ? Mem1D_5_io_output : _T_10418; // @[Mux.scala 31:69:@54155.4]
  assign _T_10348 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@53993.4 package.scala 96:25:@53994.4]
  assign _T_10420 = _T_10348 ? Mem1D_3_io_output : _T_10419; // @[Mux.scala 31:69:@54156.4]
  assign _T_10345 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@53985.4 package.scala 96:25:@53986.4]
  assign _T_10578 = RetimeWrapper_198_io_out; // @[package.scala 96:25:@54369.4 package.scala 96:25:@54370.4]
  assign _T_10582 = _T_10578 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@54379.4]
  assign _T_10575 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@54361.4 package.scala 96:25:@54362.4]
  assign _T_10583 = _T_10575 ? Mem1D_34_io_output : _T_10582; // @[Mux.scala 31:69:@54380.4]
  assign _T_10572 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@54353.4 package.scala 96:25:@54354.4]
  assign _T_10584 = _T_10572 ? Mem1D_32_io_output : _T_10583; // @[Mux.scala 31:69:@54381.4]
  assign _T_10569 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@54345.4 package.scala 96:25:@54346.4]
  assign _T_10585 = _T_10569 ? Mem1D_30_io_output : _T_10584; // @[Mux.scala 31:69:@54382.4]
  assign _T_10566 = RetimeWrapper_194_io_out; // @[package.scala 96:25:@54337.4 package.scala 96:25:@54338.4]
  assign _T_10586 = _T_10566 ? Mem1D_28_io_output : _T_10585; // @[Mux.scala 31:69:@54383.4]
  assign _T_10563 = RetimeWrapper_193_io_out; // @[package.scala 96:25:@54329.4 package.scala 96:25:@54330.4]
  assign _T_10587 = _T_10563 ? Mem1D_26_io_output : _T_10586; // @[Mux.scala 31:69:@54384.4]
  assign _T_10560 = RetimeWrapper_192_io_out; // @[package.scala 96:25:@54321.4 package.scala 96:25:@54322.4]
  assign _T_10588 = _T_10560 ? Mem1D_24_io_output : _T_10587; // @[Mux.scala 31:69:@54385.4]
  assign _T_10557 = RetimeWrapper_191_io_out; // @[package.scala 96:25:@54313.4 package.scala 96:25:@54314.4]
  assign _T_10589 = _T_10557 ? Mem1D_22_io_output : _T_10588; // @[Mux.scala 31:69:@54386.4]
  assign _T_10554 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@54305.4 package.scala 96:25:@54306.4]
  assign _T_10590 = _T_10554 ? Mem1D_20_io_output : _T_10589; // @[Mux.scala 31:69:@54387.4]
  assign _T_10551 = RetimeWrapper_189_io_out; // @[package.scala 96:25:@54297.4 package.scala 96:25:@54298.4]
  assign _T_10591 = _T_10551 ? Mem1D_18_io_output : _T_10590; // @[Mux.scala 31:69:@54388.4]
  assign _T_10548 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@54289.4 package.scala 96:25:@54290.4]
  assign _T_10592 = _T_10548 ? Mem1D_16_io_output : _T_10591; // @[Mux.scala 31:69:@54389.4]
  assign _T_10545 = RetimeWrapper_187_io_out; // @[package.scala 96:25:@54281.4 package.scala 96:25:@54282.4]
  assign _T_10593 = _T_10545 ? Mem1D_14_io_output : _T_10592; // @[Mux.scala 31:69:@54390.4]
  assign _T_10542 = RetimeWrapper_186_io_out; // @[package.scala 96:25:@54273.4 package.scala 96:25:@54274.4]
  assign _T_10594 = _T_10542 ? Mem1D_12_io_output : _T_10593; // @[Mux.scala 31:69:@54391.4]
  assign _T_10539 = RetimeWrapper_185_io_out; // @[package.scala 96:25:@54265.4 package.scala 96:25:@54266.4]
  assign _T_10595 = _T_10539 ? Mem1D_10_io_output : _T_10594; // @[Mux.scala 31:69:@54392.4]
  assign _T_10536 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@54257.4 package.scala 96:25:@54258.4]
  assign _T_10596 = _T_10536 ? Mem1D_8_io_output : _T_10595; // @[Mux.scala 31:69:@54393.4]
  assign _T_10533 = RetimeWrapper_183_io_out; // @[package.scala 96:25:@54249.4 package.scala 96:25:@54250.4]
  assign _T_10597 = _T_10533 ? Mem1D_6_io_output : _T_10596; // @[Mux.scala 31:69:@54394.4]
  assign _T_10530 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@54241.4 package.scala 96:25:@54242.4]
  assign _T_10598 = _T_10530 ? Mem1D_4_io_output : _T_10597; // @[Mux.scala 31:69:@54395.4]
  assign _T_10527 = RetimeWrapper_181_io_out; // @[package.scala 96:25:@54233.4 package.scala 96:25:@54234.4]
  assign _T_10599 = _T_10527 ? Mem1D_2_io_output : _T_10598; // @[Mux.scala 31:69:@54396.4]
  assign _T_10524 = RetimeWrapper_180_io_out; // @[package.scala 96:25:@54225.4 package.scala 96:25:@54226.4]
  assign _T_10757 = RetimeWrapper_218_io_out; // @[package.scala 96:25:@54609.4 package.scala 96:25:@54610.4]
  assign _T_10761 = _T_10757 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@54619.4]
  assign _T_10754 = RetimeWrapper_217_io_out; // @[package.scala 96:25:@54601.4 package.scala 96:25:@54602.4]
  assign _T_10762 = _T_10754 ? Mem1D_34_io_output : _T_10761; // @[Mux.scala 31:69:@54620.4]
  assign _T_10751 = RetimeWrapper_216_io_out; // @[package.scala 96:25:@54593.4 package.scala 96:25:@54594.4]
  assign _T_10763 = _T_10751 ? Mem1D_32_io_output : _T_10762; // @[Mux.scala 31:69:@54621.4]
  assign _T_10748 = RetimeWrapper_215_io_out; // @[package.scala 96:25:@54585.4 package.scala 96:25:@54586.4]
  assign _T_10764 = _T_10748 ? Mem1D_30_io_output : _T_10763; // @[Mux.scala 31:69:@54622.4]
  assign _T_10745 = RetimeWrapper_214_io_out; // @[package.scala 96:25:@54577.4 package.scala 96:25:@54578.4]
  assign _T_10765 = _T_10745 ? Mem1D_28_io_output : _T_10764; // @[Mux.scala 31:69:@54623.4]
  assign _T_10742 = RetimeWrapper_213_io_out; // @[package.scala 96:25:@54569.4 package.scala 96:25:@54570.4]
  assign _T_10766 = _T_10742 ? Mem1D_26_io_output : _T_10765; // @[Mux.scala 31:69:@54624.4]
  assign _T_10739 = RetimeWrapper_212_io_out; // @[package.scala 96:25:@54561.4 package.scala 96:25:@54562.4]
  assign _T_10767 = _T_10739 ? Mem1D_24_io_output : _T_10766; // @[Mux.scala 31:69:@54625.4]
  assign _T_10736 = RetimeWrapper_211_io_out; // @[package.scala 96:25:@54553.4 package.scala 96:25:@54554.4]
  assign _T_10768 = _T_10736 ? Mem1D_22_io_output : _T_10767; // @[Mux.scala 31:69:@54626.4]
  assign _T_10733 = RetimeWrapper_210_io_out; // @[package.scala 96:25:@54545.4 package.scala 96:25:@54546.4]
  assign _T_10769 = _T_10733 ? Mem1D_20_io_output : _T_10768; // @[Mux.scala 31:69:@54627.4]
  assign _T_10730 = RetimeWrapper_209_io_out; // @[package.scala 96:25:@54537.4 package.scala 96:25:@54538.4]
  assign _T_10770 = _T_10730 ? Mem1D_18_io_output : _T_10769; // @[Mux.scala 31:69:@54628.4]
  assign _T_10727 = RetimeWrapper_208_io_out; // @[package.scala 96:25:@54529.4 package.scala 96:25:@54530.4]
  assign _T_10771 = _T_10727 ? Mem1D_16_io_output : _T_10770; // @[Mux.scala 31:69:@54629.4]
  assign _T_10724 = RetimeWrapper_207_io_out; // @[package.scala 96:25:@54521.4 package.scala 96:25:@54522.4]
  assign _T_10772 = _T_10724 ? Mem1D_14_io_output : _T_10771; // @[Mux.scala 31:69:@54630.4]
  assign _T_10721 = RetimeWrapper_206_io_out; // @[package.scala 96:25:@54513.4 package.scala 96:25:@54514.4]
  assign _T_10773 = _T_10721 ? Mem1D_12_io_output : _T_10772; // @[Mux.scala 31:69:@54631.4]
  assign _T_10718 = RetimeWrapper_205_io_out; // @[package.scala 96:25:@54505.4 package.scala 96:25:@54506.4]
  assign _T_10774 = _T_10718 ? Mem1D_10_io_output : _T_10773; // @[Mux.scala 31:69:@54632.4]
  assign _T_10715 = RetimeWrapper_204_io_out; // @[package.scala 96:25:@54497.4 package.scala 96:25:@54498.4]
  assign _T_10775 = _T_10715 ? Mem1D_8_io_output : _T_10774; // @[Mux.scala 31:69:@54633.4]
  assign _T_10712 = RetimeWrapper_203_io_out; // @[package.scala 96:25:@54489.4 package.scala 96:25:@54490.4]
  assign _T_10776 = _T_10712 ? Mem1D_6_io_output : _T_10775; // @[Mux.scala 31:69:@54634.4]
  assign _T_10709 = RetimeWrapper_202_io_out; // @[package.scala 96:25:@54481.4 package.scala 96:25:@54482.4]
  assign _T_10777 = _T_10709 ? Mem1D_4_io_output : _T_10776; // @[Mux.scala 31:69:@54635.4]
  assign _T_10706 = RetimeWrapper_201_io_out; // @[package.scala 96:25:@54473.4 package.scala 96:25:@54474.4]
  assign _T_10778 = _T_10706 ? Mem1D_2_io_output : _T_10777; // @[Mux.scala 31:69:@54636.4]
  assign _T_10703 = RetimeWrapper_200_io_out; // @[package.scala 96:25:@54465.4 package.scala 96:25:@54466.4]
  assign _T_10936 = RetimeWrapper_238_io_out; // @[package.scala 96:25:@54849.4 package.scala 96:25:@54850.4]
  assign _T_10940 = _T_10936 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@54859.4]
  assign _T_10933 = RetimeWrapper_237_io_out; // @[package.scala 96:25:@54841.4 package.scala 96:25:@54842.4]
  assign _T_10941 = _T_10933 ? Mem1D_35_io_output : _T_10940; // @[Mux.scala 31:69:@54860.4]
  assign _T_10930 = RetimeWrapper_236_io_out; // @[package.scala 96:25:@54833.4 package.scala 96:25:@54834.4]
  assign _T_10942 = _T_10930 ? Mem1D_33_io_output : _T_10941; // @[Mux.scala 31:69:@54861.4]
  assign _T_10927 = RetimeWrapper_235_io_out; // @[package.scala 96:25:@54825.4 package.scala 96:25:@54826.4]
  assign _T_10943 = _T_10927 ? Mem1D_31_io_output : _T_10942; // @[Mux.scala 31:69:@54862.4]
  assign _T_10924 = RetimeWrapper_234_io_out; // @[package.scala 96:25:@54817.4 package.scala 96:25:@54818.4]
  assign _T_10944 = _T_10924 ? Mem1D_29_io_output : _T_10943; // @[Mux.scala 31:69:@54863.4]
  assign _T_10921 = RetimeWrapper_233_io_out; // @[package.scala 96:25:@54809.4 package.scala 96:25:@54810.4]
  assign _T_10945 = _T_10921 ? Mem1D_27_io_output : _T_10944; // @[Mux.scala 31:69:@54864.4]
  assign _T_10918 = RetimeWrapper_232_io_out; // @[package.scala 96:25:@54801.4 package.scala 96:25:@54802.4]
  assign _T_10946 = _T_10918 ? Mem1D_25_io_output : _T_10945; // @[Mux.scala 31:69:@54865.4]
  assign _T_10915 = RetimeWrapper_231_io_out; // @[package.scala 96:25:@54793.4 package.scala 96:25:@54794.4]
  assign _T_10947 = _T_10915 ? Mem1D_23_io_output : _T_10946; // @[Mux.scala 31:69:@54866.4]
  assign _T_10912 = RetimeWrapper_230_io_out; // @[package.scala 96:25:@54785.4 package.scala 96:25:@54786.4]
  assign _T_10948 = _T_10912 ? Mem1D_21_io_output : _T_10947; // @[Mux.scala 31:69:@54867.4]
  assign _T_10909 = RetimeWrapper_229_io_out; // @[package.scala 96:25:@54777.4 package.scala 96:25:@54778.4]
  assign _T_10949 = _T_10909 ? Mem1D_19_io_output : _T_10948; // @[Mux.scala 31:69:@54868.4]
  assign _T_10906 = RetimeWrapper_228_io_out; // @[package.scala 96:25:@54769.4 package.scala 96:25:@54770.4]
  assign _T_10950 = _T_10906 ? Mem1D_17_io_output : _T_10949; // @[Mux.scala 31:69:@54869.4]
  assign _T_10903 = RetimeWrapper_227_io_out; // @[package.scala 96:25:@54761.4 package.scala 96:25:@54762.4]
  assign _T_10951 = _T_10903 ? Mem1D_15_io_output : _T_10950; // @[Mux.scala 31:69:@54870.4]
  assign _T_10900 = RetimeWrapper_226_io_out; // @[package.scala 96:25:@54753.4 package.scala 96:25:@54754.4]
  assign _T_10952 = _T_10900 ? Mem1D_13_io_output : _T_10951; // @[Mux.scala 31:69:@54871.4]
  assign _T_10897 = RetimeWrapper_225_io_out; // @[package.scala 96:25:@54745.4 package.scala 96:25:@54746.4]
  assign _T_10953 = _T_10897 ? Mem1D_11_io_output : _T_10952; // @[Mux.scala 31:69:@54872.4]
  assign _T_10894 = RetimeWrapper_224_io_out; // @[package.scala 96:25:@54737.4 package.scala 96:25:@54738.4]
  assign _T_10954 = _T_10894 ? Mem1D_9_io_output : _T_10953; // @[Mux.scala 31:69:@54873.4]
  assign _T_10891 = RetimeWrapper_223_io_out; // @[package.scala 96:25:@54729.4 package.scala 96:25:@54730.4]
  assign _T_10955 = _T_10891 ? Mem1D_7_io_output : _T_10954; // @[Mux.scala 31:69:@54874.4]
  assign _T_10888 = RetimeWrapper_222_io_out; // @[package.scala 96:25:@54721.4 package.scala 96:25:@54722.4]
  assign _T_10956 = _T_10888 ? Mem1D_5_io_output : _T_10955; // @[Mux.scala 31:69:@54875.4]
  assign _T_10885 = RetimeWrapper_221_io_out; // @[package.scala 96:25:@54713.4 package.scala 96:25:@54714.4]
  assign _T_10957 = _T_10885 ? Mem1D_3_io_output : _T_10956; // @[Mux.scala 31:69:@54876.4]
  assign _T_10882 = RetimeWrapper_220_io_out; // @[package.scala 96:25:@54705.4 package.scala 96:25:@54706.4]
  assign _T_11115 = RetimeWrapper_258_io_out; // @[package.scala 96:25:@55089.4 package.scala 96:25:@55090.4]
  assign _T_11119 = _T_11115 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@55099.4]
  assign _T_11112 = RetimeWrapper_257_io_out; // @[package.scala 96:25:@55081.4 package.scala 96:25:@55082.4]
  assign _T_11120 = _T_11112 ? Mem1D_35_io_output : _T_11119; // @[Mux.scala 31:69:@55100.4]
  assign _T_11109 = RetimeWrapper_256_io_out; // @[package.scala 96:25:@55073.4 package.scala 96:25:@55074.4]
  assign _T_11121 = _T_11109 ? Mem1D_33_io_output : _T_11120; // @[Mux.scala 31:69:@55101.4]
  assign _T_11106 = RetimeWrapper_255_io_out; // @[package.scala 96:25:@55065.4 package.scala 96:25:@55066.4]
  assign _T_11122 = _T_11106 ? Mem1D_31_io_output : _T_11121; // @[Mux.scala 31:69:@55102.4]
  assign _T_11103 = RetimeWrapper_254_io_out; // @[package.scala 96:25:@55057.4 package.scala 96:25:@55058.4]
  assign _T_11123 = _T_11103 ? Mem1D_29_io_output : _T_11122; // @[Mux.scala 31:69:@55103.4]
  assign _T_11100 = RetimeWrapper_253_io_out; // @[package.scala 96:25:@55049.4 package.scala 96:25:@55050.4]
  assign _T_11124 = _T_11100 ? Mem1D_27_io_output : _T_11123; // @[Mux.scala 31:69:@55104.4]
  assign _T_11097 = RetimeWrapper_252_io_out; // @[package.scala 96:25:@55041.4 package.scala 96:25:@55042.4]
  assign _T_11125 = _T_11097 ? Mem1D_25_io_output : _T_11124; // @[Mux.scala 31:69:@55105.4]
  assign _T_11094 = RetimeWrapper_251_io_out; // @[package.scala 96:25:@55033.4 package.scala 96:25:@55034.4]
  assign _T_11126 = _T_11094 ? Mem1D_23_io_output : _T_11125; // @[Mux.scala 31:69:@55106.4]
  assign _T_11091 = RetimeWrapper_250_io_out; // @[package.scala 96:25:@55025.4 package.scala 96:25:@55026.4]
  assign _T_11127 = _T_11091 ? Mem1D_21_io_output : _T_11126; // @[Mux.scala 31:69:@55107.4]
  assign _T_11088 = RetimeWrapper_249_io_out; // @[package.scala 96:25:@55017.4 package.scala 96:25:@55018.4]
  assign _T_11128 = _T_11088 ? Mem1D_19_io_output : _T_11127; // @[Mux.scala 31:69:@55108.4]
  assign _T_11085 = RetimeWrapper_248_io_out; // @[package.scala 96:25:@55009.4 package.scala 96:25:@55010.4]
  assign _T_11129 = _T_11085 ? Mem1D_17_io_output : _T_11128; // @[Mux.scala 31:69:@55109.4]
  assign _T_11082 = RetimeWrapper_247_io_out; // @[package.scala 96:25:@55001.4 package.scala 96:25:@55002.4]
  assign _T_11130 = _T_11082 ? Mem1D_15_io_output : _T_11129; // @[Mux.scala 31:69:@55110.4]
  assign _T_11079 = RetimeWrapper_246_io_out; // @[package.scala 96:25:@54993.4 package.scala 96:25:@54994.4]
  assign _T_11131 = _T_11079 ? Mem1D_13_io_output : _T_11130; // @[Mux.scala 31:69:@55111.4]
  assign _T_11076 = RetimeWrapper_245_io_out; // @[package.scala 96:25:@54985.4 package.scala 96:25:@54986.4]
  assign _T_11132 = _T_11076 ? Mem1D_11_io_output : _T_11131; // @[Mux.scala 31:69:@55112.4]
  assign _T_11073 = RetimeWrapper_244_io_out; // @[package.scala 96:25:@54977.4 package.scala 96:25:@54978.4]
  assign _T_11133 = _T_11073 ? Mem1D_9_io_output : _T_11132; // @[Mux.scala 31:69:@55113.4]
  assign _T_11070 = RetimeWrapper_243_io_out; // @[package.scala 96:25:@54969.4 package.scala 96:25:@54970.4]
  assign _T_11134 = _T_11070 ? Mem1D_7_io_output : _T_11133; // @[Mux.scala 31:69:@55114.4]
  assign _T_11067 = RetimeWrapper_242_io_out; // @[package.scala 96:25:@54961.4 package.scala 96:25:@54962.4]
  assign _T_11135 = _T_11067 ? Mem1D_5_io_output : _T_11134; // @[Mux.scala 31:69:@55115.4]
  assign _T_11064 = RetimeWrapper_241_io_out; // @[package.scala 96:25:@54953.4 package.scala 96:25:@54954.4]
  assign _T_11136 = _T_11064 ? Mem1D_3_io_output : _T_11135; // @[Mux.scala 31:69:@55116.4]
  assign _T_11061 = RetimeWrapper_240_io_out; // @[package.scala 96:25:@54945.4 package.scala 96:25:@54946.4]
  assign _T_11294 = RetimeWrapper_278_io_out; // @[package.scala 96:25:@55329.4 package.scala 96:25:@55330.4]
  assign _T_11298 = _T_11294 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@55339.4]
  assign _T_11291 = RetimeWrapper_277_io_out; // @[package.scala 96:25:@55321.4 package.scala 96:25:@55322.4]
  assign _T_11299 = _T_11291 ? Mem1D_34_io_output : _T_11298; // @[Mux.scala 31:69:@55340.4]
  assign _T_11288 = RetimeWrapper_276_io_out; // @[package.scala 96:25:@55313.4 package.scala 96:25:@55314.4]
  assign _T_11300 = _T_11288 ? Mem1D_32_io_output : _T_11299; // @[Mux.scala 31:69:@55341.4]
  assign _T_11285 = RetimeWrapper_275_io_out; // @[package.scala 96:25:@55305.4 package.scala 96:25:@55306.4]
  assign _T_11301 = _T_11285 ? Mem1D_30_io_output : _T_11300; // @[Mux.scala 31:69:@55342.4]
  assign _T_11282 = RetimeWrapper_274_io_out; // @[package.scala 96:25:@55297.4 package.scala 96:25:@55298.4]
  assign _T_11302 = _T_11282 ? Mem1D_28_io_output : _T_11301; // @[Mux.scala 31:69:@55343.4]
  assign _T_11279 = RetimeWrapper_273_io_out; // @[package.scala 96:25:@55289.4 package.scala 96:25:@55290.4]
  assign _T_11303 = _T_11279 ? Mem1D_26_io_output : _T_11302; // @[Mux.scala 31:69:@55344.4]
  assign _T_11276 = RetimeWrapper_272_io_out; // @[package.scala 96:25:@55281.4 package.scala 96:25:@55282.4]
  assign _T_11304 = _T_11276 ? Mem1D_24_io_output : _T_11303; // @[Mux.scala 31:69:@55345.4]
  assign _T_11273 = RetimeWrapper_271_io_out; // @[package.scala 96:25:@55273.4 package.scala 96:25:@55274.4]
  assign _T_11305 = _T_11273 ? Mem1D_22_io_output : _T_11304; // @[Mux.scala 31:69:@55346.4]
  assign _T_11270 = RetimeWrapper_270_io_out; // @[package.scala 96:25:@55265.4 package.scala 96:25:@55266.4]
  assign _T_11306 = _T_11270 ? Mem1D_20_io_output : _T_11305; // @[Mux.scala 31:69:@55347.4]
  assign _T_11267 = RetimeWrapper_269_io_out; // @[package.scala 96:25:@55257.4 package.scala 96:25:@55258.4]
  assign _T_11307 = _T_11267 ? Mem1D_18_io_output : _T_11306; // @[Mux.scala 31:69:@55348.4]
  assign _T_11264 = RetimeWrapper_268_io_out; // @[package.scala 96:25:@55249.4 package.scala 96:25:@55250.4]
  assign _T_11308 = _T_11264 ? Mem1D_16_io_output : _T_11307; // @[Mux.scala 31:69:@55349.4]
  assign _T_11261 = RetimeWrapper_267_io_out; // @[package.scala 96:25:@55241.4 package.scala 96:25:@55242.4]
  assign _T_11309 = _T_11261 ? Mem1D_14_io_output : _T_11308; // @[Mux.scala 31:69:@55350.4]
  assign _T_11258 = RetimeWrapper_266_io_out; // @[package.scala 96:25:@55233.4 package.scala 96:25:@55234.4]
  assign _T_11310 = _T_11258 ? Mem1D_12_io_output : _T_11309; // @[Mux.scala 31:69:@55351.4]
  assign _T_11255 = RetimeWrapper_265_io_out; // @[package.scala 96:25:@55225.4 package.scala 96:25:@55226.4]
  assign _T_11311 = _T_11255 ? Mem1D_10_io_output : _T_11310; // @[Mux.scala 31:69:@55352.4]
  assign _T_11252 = RetimeWrapper_264_io_out; // @[package.scala 96:25:@55217.4 package.scala 96:25:@55218.4]
  assign _T_11312 = _T_11252 ? Mem1D_8_io_output : _T_11311; // @[Mux.scala 31:69:@55353.4]
  assign _T_11249 = RetimeWrapper_263_io_out; // @[package.scala 96:25:@55209.4 package.scala 96:25:@55210.4]
  assign _T_11313 = _T_11249 ? Mem1D_6_io_output : _T_11312; // @[Mux.scala 31:69:@55354.4]
  assign _T_11246 = RetimeWrapper_262_io_out; // @[package.scala 96:25:@55201.4 package.scala 96:25:@55202.4]
  assign _T_11314 = _T_11246 ? Mem1D_4_io_output : _T_11313; // @[Mux.scala 31:69:@55355.4]
  assign _T_11243 = RetimeWrapper_261_io_out; // @[package.scala 96:25:@55193.4 package.scala 96:25:@55194.4]
  assign _T_11315 = _T_11243 ? Mem1D_2_io_output : _T_11314; // @[Mux.scala 31:69:@55356.4]
  assign _T_11240 = RetimeWrapper_260_io_out; // @[package.scala 96:25:@55185.4 package.scala 96:25:@55186.4]
  assign _T_11473 = RetimeWrapper_298_io_out; // @[package.scala 96:25:@55569.4 package.scala 96:25:@55570.4]
  assign _T_11477 = _T_11473 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@55579.4]
  assign _T_11470 = RetimeWrapper_297_io_out; // @[package.scala 96:25:@55561.4 package.scala 96:25:@55562.4]
  assign _T_11478 = _T_11470 ? Mem1D_35_io_output : _T_11477; // @[Mux.scala 31:69:@55580.4]
  assign _T_11467 = RetimeWrapper_296_io_out; // @[package.scala 96:25:@55553.4 package.scala 96:25:@55554.4]
  assign _T_11479 = _T_11467 ? Mem1D_33_io_output : _T_11478; // @[Mux.scala 31:69:@55581.4]
  assign _T_11464 = RetimeWrapper_295_io_out; // @[package.scala 96:25:@55545.4 package.scala 96:25:@55546.4]
  assign _T_11480 = _T_11464 ? Mem1D_31_io_output : _T_11479; // @[Mux.scala 31:69:@55582.4]
  assign _T_11461 = RetimeWrapper_294_io_out; // @[package.scala 96:25:@55537.4 package.scala 96:25:@55538.4]
  assign _T_11481 = _T_11461 ? Mem1D_29_io_output : _T_11480; // @[Mux.scala 31:69:@55583.4]
  assign _T_11458 = RetimeWrapper_293_io_out; // @[package.scala 96:25:@55529.4 package.scala 96:25:@55530.4]
  assign _T_11482 = _T_11458 ? Mem1D_27_io_output : _T_11481; // @[Mux.scala 31:69:@55584.4]
  assign _T_11455 = RetimeWrapper_292_io_out; // @[package.scala 96:25:@55521.4 package.scala 96:25:@55522.4]
  assign _T_11483 = _T_11455 ? Mem1D_25_io_output : _T_11482; // @[Mux.scala 31:69:@55585.4]
  assign _T_11452 = RetimeWrapper_291_io_out; // @[package.scala 96:25:@55513.4 package.scala 96:25:@55514.4]
  assign _T_11484 = _T_11452 ? Mem1D_23_io_output : _T_11483; // @[Mux.scala 31:69:@55586.4]
  assign _T_11449 = RetimeWrapper_290_io_out; // @[package.scala 96:25:@55505.4 package.scala 96:25:@55506.4]
  assign _T_11485 = _T_11449 ? Mem1D_21_io_output : _T_11484; // @[Mux.scala 31:69:@55587.4]
  assign _T_11446 = RetimeWrapper_289_io_out; // @[package.scala 96:25:@55497.4 package.scala 96:25:@55498.4]
  assign _T_11486 = _T_11446 ? Mem1D_19_io_output : _T_11485; // @[Mux.scala 31:69:@55588.4]
  assign _T_11443 = RetimeWrapper_288_io_out; // @[package.scala 96:25:@55489.4 package.scala 96:25:@55490.4]
  assign _T_11487 = _T_11443 ? Mem1D_17_io_output : _T_11486; // @[Mux.scala 31:69:@55589.4]
  assign _T_11440 = RetimeWrapper_287_io_out; // @[package.scala 96:25:@55481.4 package.scala 96:25:@55482.4]
  assign _T_11488 = _T_11440 ? Mem1D_15_io_output : _T_11487; // @[Mux.scala 31:69:@55590.4]
  assign _T_11437 = RetimeWrapper_286_io_out; // @[package.scala 96:25:@55473.4 package.scala 96:25:@55474.4]
  assign _T_11489 = _T_11437 ? Mem1D_13_io_output : _T_11488; // @[Mux.scala 31:69:@55591.4]
  assign _T_11434 = RetimeWrapper_285_io_out; // @[package.scala 96:25:@55465.4 package.scala 96:25:@55466.4]
  assign _T_11490 = _T_11434 ? Mem1D_11_io_output : _T_11489; // @[Mux.scala 31:69:@55592.4]
  assign _T_11431 = RetimeWrapper_284_io_out; // @[package.scala 96:25:@55457.4 package.scala 96:25:@55458.4]
  assign _T_11491 = _T_11431 ? Mem1D_9_io_output : _T_11490; // @[Mux.scala 31:69:@55593.4]
  assign _T_11428 = RetimeWrapper_283_io_out; // @[package.scala 96:25:@55449.4 package.scala 96:25:@55450.4]
  assign _T_11492 = _T_11428 ? Mem1D_7_io_output : _T_11491; // @[Mux.scala 31:69:@55594.4]
  assign _T_11425 = RetimeWrapper_282_io_out; // @[package.scala 96:25:@55441.4 package.scala 96:25:@55442.4]
  assign _T_11493 = _T_11425 ? Mem1D_5_io_output : _T_11492; // @[Mux.scala 31:69:@55595.4]
  assign _T_11422 = RetimeWrapper_281_io_out; // @[package.scala 96:25:@55433.4 package.scala 96:25:@55434.4]
  assign _T_11494 = _T_11422 ? Mem1D_3_io_output : _T_11493; // @[Mux.scala 31:69:@55596.4]
  assign _T_11419 = RetimeWrapper_280_io_out; // @[package.scala 96:25:@55425.4 package.scala 96:25:@55426.4]
  assign _T_11652 = RetimeWrapper_318_io_out; // @[package.scala 96:25:@55809.4 package.scala 96:25:@55810.4]
  assign _T_11656 = _T_11652 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@55819.4]
  assign _T_11649 = RetimeWrapper_317_io_out; // @[package.scala 96:25:@55801.4 package.scala 96:25:@55802.4]
  assign _T_11657 = _T_11649 ? Mem1D_34_io_output : _T_11656; // @[Mux.scala 31:69:@55820.4]
  assign _T_11646 = RetimeWrapper_316_io_out; // @[package.scala 96:25:@55793.4 package.scala 96:25:@55794.4]
  assign _T_11658 = _T_11646 ? Mem1D_32_io_output : _T_11657; // @[Mux.scala 31:69:@55821.4]
  assign _T_11643 = RetimeWrapper_315_io_out; // @[package.scala 96:25:@55785.4 package.scala 96:25:@55786.4]
  assign _T_11659 = _T_11643 ? Mem1D_30_io_output : _T_11658; // @[Mux.scala 31:69:@55822.4]
  assign _T_11640 = RetimeWrapper_314_io_out; // @[package.scala 96:25:@55777.4 package.scala 96:25:@55778.4]
  assign _T_11660 = _T_11640 ? Mem1D_28_io_output : _T_11659; // @[Mux.scala 31:69:@55823.4]
  assign _T_11637 = RetimeWrapper_313_io_out; // @[package.scala 96:25:@55769.4 package.scala 96:25:@55770.4]
  assign _T_11661 = _T_11637 ? Mem1D_26_io_output : _T_11660; // @[Mux.scala 31:69:@55824.4]
  assign _T_11634 = RetimeWrapper_312_io_out; // @[package.scala 96:25:@55761.4 package.scala 96:25:@55762.4]
  assign _T_11662 = _T_11634 ? Mem1D_24_io_output : _T_11661; // @[Mux.scala 31:69:@55825.4]
  assign _T_11631 = RetimeWrapper_311_io_out; // @[package.scala 96:25:@55753.4 package.scala 96:25:@55754.4]
  assign _T_11663 = _T_11631 ? Mem1D_22_io_output : _T_11662; // @[Mux.scala 31:69:@55826.4]
  assign _T_11628 = RetimeWrapper_310_io_out; // @[package.scala 96:25:@55745.4 package.scala 96:25:@55746.4]
  assign _T_11664 = _T_11628 ? Mem1D_20_io_output : _T_11663; // @[Mux.scala 31:69:@55827.4]
  assign _T_11625 = RetimeWrapper_309_io_out; // @[package.scala 96:25:@55737.4 package.scala 96:25:@55738.4]
  assign _T_11665 = _T_11625 ? Mem1D_18_io_output : _T_11664; // @[Mux.scala 31:69:@55828.4]
  assign _T_11622 = RetimeWrapper_308_io_out; // @[package.scala 96:25:@55729.4 package.scala 96:25:@55730.4]
  assign _T_11666 = _T_11622 ? Mem1D_16_io_output : _T_11665; // @[Mux.scala 31:69:@55829.4]
  assign _T_11619 = RetimeWrapper_307_io_out; // @[package.scala 96:25:@55721.4 package.scala 96:25:@55722.4]
  assign _T_11667 = _T_11619 ? Mem1D_14_io_output : _T_11666; // @[Mux.scala 31:69:@55830.4]
  assign _T_11616 = RetimeWrapper_306_io_out; // @[package.scala 96:25:@55713.4 package.scala 96:25:@55714.4]
  assign _T_11668 = _T_11616 ? Mem1D_12_io_output : _T_11667; // @[Mux.scala 31:69:@55831.4]
  assign _T_11613 = RetimeWrapper_305_io_out; // @[package.scala 96:25:@55705.4 package.scala 96:25:@55706.4]
  assign _T_11669 = _T_11613 ? Mem1D_10_io_output : _T_11668; // @[Mux.scala 31:69:@55832.4]
  assign _T_11610 = RetimeWrapper_304_io_out; // @[package.scala 96:25:@55697.4 package.scala 96:25:@55698.4]
  assign _T_11670 = _T_11610 ? Mem1D_8_io_output : _T_11669; // @[Mux.scala 31:69:@55833.4]
  assign _T_11607 = RetimeWrapper_303_io_out; // @[package.scala 96:25:@55689.4 package.scala 96:25:@55690.4]
  assign _T_11671 = _T_11607 ? Mem1D_6_io_output : _T_11670; // @[Mux.scala 31:69:@55834.4]
  assign _T_11604 = RetimeWrapper_302_io_out; // @[package.scala 96:25:@55681.4 package.scala 96:25:@55682.4]
  assign _T_11672 = _T_11604 ? Mem1D_4_io_output : _T_11671; // @[Mux.scala 31:69:@55835.4]
  assign _T_11601 = RetimeWrapper_301_io_out; // @[package.scala 96:25:@55673.4 package.scala 96:25:@55674.4]
  assign _T_11673 = _T_11601 ? Mem1D_2_io_output : _T_11672; // @[Mux.scala 31:69:@55836.4]
  assign _T_11598 = RetimeWrapper_300_io_out; // @[package.scala 96:25:@55665.4 package.scala 96:25:@55666.4]
  assign _T_11831 = RetimeWrapper_338_io_out; // @[package.scala 96:25:@56049.4 package.scala 96:25:@56050.4]
  assign _T_11835 = _T_11831 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@56059.4]
  assign _T_11828 = RetimeWrapper_337_io_out; // @[package.scala 96:25:@56041.4 package.scala 96:25:@56042.4]
  assign _T_11836 = _T_11828 ? Mem1D_34_io_output : _T_11835; // @[Mux.scala 31:69:@56060.4]
  assign _T_11825 = RetimeWrapper_336_io_out; // @[package.scala 96:25:@56033.4 package.scala 96:25:@56034.4]
  assign _T_11837 = _T_11825 ? Mem1D_32_io_output : _T_11836; // @[Mux.scala 31:69:@56061.4]
  assign _T_11822 = RetimeWrapper_335_io_out; // @[package.scala 96:25:@56025.4 package.scala 96:25:@56026.4]
  assign _T_11838 = _T_11822 ? Mem1D_30_io_output : _T_11837; // @[Mux.scala 31:69:@56062.4]
  assign _T_11819 = RetimeWrapper_334_io_out; // @[package.scala 96:25:@56017.4 package.scala 96:25:@56018.4]
  assign _T_11839 = _T_11819 ? Mem1D_28_io_output : _T_11838; // @[Mux.scala 31:69:@56063.4]
  assign _T_11816 = RetimeWrapper_333_io_out; // @[package.scala 96:25:@56009.4 package.scala 96:25:@56010.4]
  assign _T_11840 = _T_11816 ? Mem1D_26_io_output : _T_11839; // @[Mux.scala 31:69:@56064.4]
  assign _T_11813 = RetimeWrapper_332_io_out; // @[package.scala 96:25:@56001.4 package.scala 96:25:@56002.4]
  assign _T_11841 = _T_11813 ? Mem1D_24_io_output : _T_11840; // @[Mux.scala 31:69:@56065.4]
  assign _T_11810 = RetimeWrapper_331_io_out; // @[package.scala 96:25:@55993.4 package.scala 96:25:@55994.4]
  assign _T_11842 = _T_11810 ? Mem1D_22_io_output : _T_11841; // @[Mux.scala 31:69:@56066.4]
  assign _T_11807 = RetimeWrapper_330_io_out; // @[package.scala 96:25:@55985.4 package.scala 96:25:@55986.4]
  assign _T_11843 = _T_11807 ? Mem1D_20_io_output : _T_11842; // @[Mux.scala 31:69:@56067.4]
  assign _T_11804 = RetimeWrapper_329_io_out; // @[package.scala 96:25:@55977.4 package.scala 96:25:@55978.4]
  assign _T_11844 = _T_11804 ? Mem1D_18_io_output : _T_11843; // @[Mux.scala 31:69:@56068.4]
  assign _T_11801 = RetimeWrapper_328_io_out; // @[package.scala 96:25:@55969.4 package.scala 96:25:@55970.4]
  assign _T_11845 = _T_11801 ? Mem1D_16_io_output : _T_11844; // @[Mux.scala 31:69:@56069.4]
  assign _T_11798 = RetimeWrapper_327_io_out; // @[package.scala 96:25:@55961.4 package.scala 96:25:@55962.4]
  assign _T_11846 = _T_11798 ? Mem1D_14_io_output : _T_11845; // @[Mux.scala 31:69:@56070.4]
  assign _T_11795 = RetimeWrapper_326_io_out; // @[package.scala 96:25:@55953.4 package.scala 96:25:@55954.4]
  assign _T_11847 = _T_11795 ? Mem1D_12_io_output : _T_11846; // @[Mux.scala 31:69:@56071.4]
  assign _T_11792 = RetimeWrapper_325_io_out; // @[package.scala 96:25:@55945.4 package.scala 96:25:@55946.4]
  assign _T_11848 = _T_11792 ? Mem1D_10_io_output : _T_11847; // @[Mux.scala 31:69:@56072.4]
  assign _T_11789 = RetimeWrapper_324_io_out; // @[package.scala 96:25:@55937.4 package.scala 96:25:@55938.4]
  assign _T_11849 = _T_11789 ? Mem1D_8_io_output : _T_11848; // @[Mux.scala 31:69:@56073.4]
  assign _T_11786 = RetimeWrapper_323_io_out; // @[package.scala 96:25:@55929.4 package.scala 96:25:@55930.4]
  assign _T_11850 = _T_11786 ? Mem1D_6_io_output : _T_11849; // @[Mux.scala 31:69:@56074.4]
  assign _T_11783 = RetimeWrapper_322_io_out; // @[package.scala 96:25:@55921.4 package.scala 96:25:@55922.4]
  assign _T_11851 = _T_11783 ? Mem1D_4_io_output : _T_11850; // @[Mux.scala 31:69:@56075.4]
  assign _T_11780 = RetimeWrapper_321_io_out; // @[package.scala 96:25:@55913.4 package.scala 96:25:@55914.4]
  assign _T_11852 = _T_11780 ? Mem1D_2_io_output : _T_11851; // @[Mux.scala 31:69:@56076.4]
  assign _T_11777 = RetimeWrapper_320_io_out; // @[package.scala 96:25:@55905.4 package.scala 96:25:@55906.4]
  assign _T_12010 = RetimeWrapper_358_io_out; // @[package.scala 96:25:@56289.4 package.scala 96:25:@56290.4]
  assign _T_12014 = _T_12010 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@56299.4]
  assign _T_12007 = RetimeWrapper_357_io_out; // @[package.scala 96:25:@56281.4 package.scala 96:25:@56282.4]
  assign _T_12015 = _T_12007 ? Mem1D_34_io_output : _T_12014; // @[Mux.scala 31:69:@56300.4]
  assign _T_12004 = RetimeWrapper_356_io_out; // @[package.scala 96:25:@56273.4 package.scala 96:25:@56274.4]
  assign _T_12016 = _T_12004 ? Mem1D_32_io_output : _T_12015; // @[Mux.scala 31:69:@56301.4]
  assign _T_12001 = RetimeWrapper_355_io_out; // @[package.scala 96:25:@56265.4 package.scala 96:25:@56266.4]
  assign _T_12017 = _T_12001 ? Mem1D_30_io_output : _T_12016; // @[Mux.scala 31:69:@56302.4]
  assign _T_11998 = RetimeWrapper_354_io_out; // @[package.scala 96:25:@56257.4 package.scala 96:25:@56258.4]
  assign _T_12018 = _T_11998 ? Mem1D_28_io_output : _T_12017; // @[Mux.scala 31:69:@56303.4]
  assign _T_11995 = RetimeWrapper_353_io_out; // @[package.scala 96:25:@56249.4 package.scala 96:25:@56250.4]
  assign _T_12019 = _T_11995 ? Mem1D_26_io_output : _T_12018; // @[Mux.scala 31:69:@56304.4]
  assign _T_11992 = RetimeWrapper_352_io_out; // @[package.scala 96:25:@56241.4 package.scala 96:25:@56242.4]
  assign _T_12020 = _T_11992 ? Mem1D_24_io_output : _T_12019; // @[Mux.scala 31:69:@56305.4]
  assign _T_11989 = RetimeWrapper_351_io_out; // @[package.scala 96:25:@56233.4 package.scala 96:25:@56234.4]
  assign _T_12021 = _T_11989 ? Mem1D_22_io_output : _T_12020; // @[Mux.scala 31:69:@56306.4]
  assign _T_11986 = RetimeWrapper_350_io_out; // @[package.scala 96:25:@56225.4 package.scala 96:25:@56226.4]
  assign _T_12022 = _T_11986 ? Mem1D_20_io_output : _T_12021; // @[Mux.scala 31:69:@56307.4]
  assign _T_11983 = RetimeWrapper_349_io_out; // @[package.scala 96:25:@56217.4 package.scala 96:25:@56218.4]
  assign _T_12023 = _T_11983 ? Mem1D_18_io_output : _T_12022; // @[Mux.scala 31:69:@56308.4]
  assign _T_11980 = RetimeWrapper_348_io_out; // @[package.scala 96:25:@56209.4 package.scala 96:25:@56210.4]
  assign _T_12024 = _T_11980 ? Mem1D_16_io_output : _T_12023; // @[Mux.scala 31:69:@56309.4]
  assign _T_11977 = RetimeWrapper_347_io_out; // @[package.scala 96:25:@56201.4 package.scala 96:25:@56202.4]
  assign _T_12025 = _T_11977 ? Mem1D_14_io_output : _T_12024; // @[Mux.scala 31:69:@56310.4]
  assign _T_11974 = RetimeWrapper_346_io_out; // @[package.scala 96:25:@56193.4 package.scala 96:25:@56194.4]
  assign _T_12026 = _T_11974 ? Mem1D_12_io_output : _T_12025; // @[Mux.scala 31:69:@56311.4]
  assign _T_11971 = RetimeWrapper_345_io_out; // @[package.scala 96:25:@56185.4 package.scala 96:25:@56186.4]
  assign _T_12027 = _T_11971 ? Mem1D_10_io_output : _T_12026; // @[Mux.scala 31:69:@56312.4]
  assign _T_11968 = RetimeWrapper_344_io_out; // @[package.scala 96:25:@56177.4 package.scala 96:25:@56178.4]
  assign _T_12028 = _T_11968 ? Mem1D_8_io_output : _T_12027; // @[Mux.scala 31:69:@56313.4]
  assign _T_11965 = RetimeWrapper_343_io_out; // @[package.scala 96:25:@56169.4 package.scala 96:25:@56170.4]
  assign _T_12029 = _T_11965 ? Mem1D_6_io_output : _T_12028; // @[Mux.scala 31:69:@56314.4]
  assign _T_11962 = RetimeWrapper_342_io_out; // @[package.scala 96:25:@56161.4 package.scala 96:25:@56162.4]
  assign _T_12030 = _T_11962 ? Mem1D_4_io_output : _T_12029; // @[Mux.scala 31:69:@56315.4]
  assign _T_11959 = RetimeWrapper_341_io_out; // @[package.scala 96:25:@56153.4 package.scala 96:25:@56154.4]
  assign _T_12031 = _T_11959 ? Mem1D_2_io_output : _T_12030; // @[Mux.scala 31:69:@56316.4]
  assign _T_11956 = RetimeWrapper_340_io_out; // @[package.scala 96:25:@56145.4 package.scala 96:25:@56146.4]
  assign _T_12189 = RetimeWrapper_378_io_out; // @[package.scala 96:25:@56529.4 package.scala 96:25:@56530.4]
  assign _T_12193 = _T_12189 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@56539.4]
  assign _T_12186 = RetimeWrapper_377_io_out; // @[package.scala 96:25:@56521.4 package.scala 96:25:@56522.4]
  assign _T_12194 = _T_12186 ? Mem1D_35_io_output : _T_12193; // @[Mux.scala 31:69:@56540.4]
  assign _T_12183 = RetimeWrapper_376_io_out; // @[package.scala 96:25:@56513.4 package.scala 96:25:@56514.4]
  assign _T_12195 = _T_12183 ? Mem1D_33_io_output : _T_12194; // @[Mux.scala 31:69:@56541.4]
  assign _T_12180 = RetimeWrapper_375_io_out; // @[package.scala 96:25:@56505.4 package.scala 96:25:@56506.4]
  assign _T_12196 = _T_12180 ? Mem1D_31_io_output : _T_12195; // @[Mux.scala 31:69:@56542.4]
  assign _T_12177 = RetimeWrapper_374_io_out; // @[package.scala 96:25:@56497.4 package.scala 96:25:@56498.4]
  assign _T_12197 = _T_12177 ? Mem1D_29_io_output : _T_12196; // @[Mux.scala 31:69:@56543.4]
  assign _T_12174 = RetimeWrapper_373_io_out; // @[package.scala 96:25:@56489.4 package.scala 96:25:@56490.4]
  assign _T_12198 = _T_12174 ? Mem1D_27_io_output : _T_12197; // @[Mux.scala 31:69:@56544.4]
  assign _T_12171 = RetimeWrapper_372_io_out; // @[package.scala 96:25:@56481.4 package.scala 96:25:@56482.4]
  assign _T_12199 = _T_12171 ? Mem1D_25_io_output : _T_12198; // @[Mux.scala 31:69:@56545.4]
  assign _T_12168 = RetimeWrapper_371_io_out; // @[package.scala 96:25:@56473.4 package.scala 96:25:@56474.4]
  assign _T_12200 = _T_12168 ? Mem1D_23_io_output : _T_12199; // @[Mux.scala 31:69:@56546.4]
  assign _T_12165 = RetimeWrapper_370_io_out; // @[package.scala 96:25:@56465.4 package.scala 96:25:@56466.4]
  assign _T_12201 = _T_12165 ? Mem1D_21_io_output : _T_12200; // @[Mux.scala 31:69:@56547.4]
  assign _T_12162 = RetimeWrapper_369_io_out; // @[package.scala 96:25:@56457.4 package.scala 96:25:@56458.4]
  assign _T_12202 = _T_12162 ? Mem1D_19_io_output : _T_12201; // @[Mux.scala 31:69:@56548.4]
  assign _T_12159 = RetimeWrapper_368_io_out; // @[package.scala 96:25:@56449.4 package.scala 96:25:@56450.4]
  assign _T_12203 = _T_12159 ? Mem1D_17_io_output : _T_12202; // @[Mux.scala 31:69:@56549.4]
  assign _T_12156 = RetimeWrapper_367_io_out; // @[package.scala 96:25:@56441.4 package.scala 96:25:@56442.4]
  assign _T_12204 = _T_12156 ? Mem1D_15_io_output : _T_12203; // @[Mux.scala 31:69:@56550.4]
  assign _T_12153 = RetimeWrapper_366_io_out; // @[package.scala 96:25:@56433.4 package.scala 96:25:@56434.4]
  assign _T_12205 = _T_12153 ? Mem1D_13_io_output : _T_12204; // @[Mux.scala 31:69:@56551.4]
  assign _T_12150 = RetimeWrapper_365_io_out; // @[package.scala 96:25:@56425.4 package.scala 96:25:@56426.4]
  assign _T_12206 = _T_12150 ? Mem1D_11_io_output : _T_12205; // @[Mux.scala 31:69:@56552.4]
  assign _T_12147 = RetimeWrapper_364_io_out; // @[package.scala 96:25:@56417.4 package.scala 96:25:@56418.4]
  assign _T_12207 = _T_12147 ? Mem1D_9_io_output : _T_12206; // @[Mux.scala 31:69:@56553.4]
  assign _T_12144 = RetimeWrapper_363_io_out; // @[package.scala 96:25:@56409.4 package.scala 96:25:@56410.4]
  assign _T_12208 = _T_12144 ? Mem1D_7_io_output : _T_12207; // @[Mux.scala 31:69:@56554.4]
  assign _T_12141 = RetimeWrapper_362_io_out; // @[package.scala 96:25:@56401.4 package.scala 96:25:@56402.4]
  assign _T_12209 = _T_12141 ? Mem1D_5_io_output : _T_12208; // @[Mux.scala 31:69:@56555.4]
  assign _T_12138 = RetimeWrapper_361_io_out; // @[package.scala 96:25:@56393.4 package.scala 96:25:@56394.4]
  assign _T_12210 = _T_12138 ? Mem1D_3_io_output : _T_12209; // @[Mux.scala 31:69:@56556.4]
  assign _T_12135 = RetimeWrapper_360_io_out; // @[package.scala 96:25:@56385.4 package.scala 96:25:@56386.4]
  assign _T_12368 = RetimeWrapper_398_io_out; // @[package.scala 96:25:@56769.4 package.scala 96:25:@56770.4]
  assign _T_12372 = _T_12368 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@56779.4]
  assign _T_12365 = RetimeWrapper_397_io_out; // @[package.scala 96:25:@56761.4 package.scala 96:25:@56762.4]
  assign _T_12373 = _T_12365 ? Mem1D_34_io_output : _T_12372; // @[Mux.scala 31:69:@56780.4]
  assign _T_12362 = RetimeWrapper_396_io_out; // @[package.scala 96:25:@56753.4 package.scala 96:25:@56754.4]
  assign _T_12374 = _T_12362 ? Mem1D_32_io_output : _T_12373; // @[Mux.scala 31:69:@56781.4]
  assign _T_12359 = RetimeWrapper_395_io_out; // @[package.scala 96:25:@56745.4 package.scala 96:25:@56746.4]
  assign _T_12375 = _T_12359 ? Mem1D_30_io_output : _T_12374; // @[Mux.scala 31:69:@56782.4]
  assign _T_12356 = RetimeWrapper_394_io_out; // @[package.scala 96:25:@56737.4 package.scala 96:25:@56738.4]
  assign _T_12376 = _T_12356 ? Mem1D_28_io_output : _T_12375; // @[Mux.scala 31:69:@56783.4]
  assign _T_12353 = RetimeWrapper_393_io_out; // @[package.scala 96:25:@56729.4 package.scala 96:25:@56730.4]
  assign _T_12377 = _T_12353 ? Mem1D_26_io_output : _T_12376; // @[Mux.scala 31:69:@56784.4]
  assign _T_12350 = RetimeWrapper_392_io_out; // @[package.scala 96:25:@56721.4 package.scala 96:25:@56722.4]
  assign _T_12378 = _T_12350 ? Mem1D_24_io_output : _T_12377; // @[Mux.scala 31:69:@56785.4]
  assign _T_12347 = RetimeWrapper_391_io_out; // @[package.scala 96:25:@56713.4 package.scala 96:25:@56714.4]
  assign _T_12379 = _T_12347 ? Mem1D_22_io_output : _T_12378; // @[Mux.scala 31:69:@56786.4]
  assign _T_12344 = RetimeWrapper_390_io_out; // @[package.scala 96:25:@56705.4 package.scala 96:25:@56706.4]
  assign _T_12380 = _T_12344 ? Mem1D_20_io_output : _T_12379; // @[Mux.scala 31:69:@56787.4]
  assign _T_12341 = RetimeWrapper_389_io_out; // @[package.scala 96:25:@56697.4 package.scala 96:25:@56698.4]
  assign _T_12381 = _T_12341 ? Mem1D_18_io_output : _T_12380; // @[Mux.scala 31:69:@56788.4]
  assign _T_12338 = RetimeWrapper_388_io_out; // @[package.scala 96:25:@56689.4 package.scala 96:25:@56690.4]
  assign _T_12382 = _T_12338 ? Mem1D_16_io_output : _T_12381; // @[Mux.scala 31:69:@56789.4]
  assign _T_12335 = RetimeWrapper_387_io_out; // @[package.scala 96:25:@56681.4 package.scala 96:25:@56682.4]
  assign _T_12383 = _T_12335 ? Mem1D_14_io_output : _T_12382; // @[Mux.scala 31:69:@56790.4]
  assign _T_12332 = RetimeWrapper_386_io_out; // @[package.scala 96:25:@56673.4 package.scala 96:25:@56674.4]
  assign _T_12384 = _T_12332 ? Mem1D_12_io_output : _T_12383; // @[Mux.scala 31:69:@56791.4]
  assign _T_12329 = RetimeWrapper_385_io_out; // @[package.scala 96:25:@56665.4 package.scala 96:25:@56666.4]
  assign _T_12385 = _T_12329 ? Mem1D_10_io_output : _T_12384; // @[Mux.scala 31:69:@56792.4]
  assign _T_12326 = RetimeWrapper_384_io_out; // @[package.scala 96:25:@56657.4 package.scala 96:25:@56658.4]
  assign _T_12386 = _T_12326 ? Mem1D_8_io_output : _T_12385; // @[Mux.scala 31:69:@56793.4]
  assign _T_12323 = RetimeWrapper_383_io_out; // @[package.scala 96:25:@56649.4 package.scala 96:25:@56650.4]
  assign _T_12387 = _T_12323 ? Mem1D_6_io_output : _T_12386; // @[Mux.scala 31:69:@56794.4]
  assign _T_12320 = RetimeWrapper_382_io_out; // @[package.scala 96:25:@56641.4 package.scala 96:25:@56642.4]
  assign _T_12388 = _T_12320 ? Mem1D_4_io_output : _T_12387; // @[Mux.scala 31:69:@56795.4]
  assign _T_12317 = RetimeWrapper_381_io_out; // @[package.scala 96:25:@56633.4 package.scala 96:25:@56634.4]
  assign _T_12389 = _T_12317 ? Mem1D_2_io_output : _T_12388; // @[Mux.scala 31:69:@56796.4]
  assign _T_12314 = RetimeWrapper_380_io_out; // @[package.scala 96:25:@56625.4 package.scala 96:25:@56626.4]
  assign _T_12547 = RetimeWrapper_418_io_out; // @[package.scala 96:25:@57009.4 package.scala 96:25:@57010.4]
  assign _T_12551 = _T_12547 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@57019.4]
  assign _T_12544 = RetimeWrapper_417_io_out; // @[package.scala 96:25:@57001.4 package.scala 96:25:@57002.4]
  assign _T_12552 = _T_12544 ? Mem1D_35_io_output : _T_12551; // @[Mux.scala 31:69:@57020.4]
  assign _T_12541 = RetimeWrapper_416_io_out; // @[package.scala 96:25:@56993.4 package.scala 96:25:@56994.4]
  assign _T_12553 = _T_12541 ? Mem1D_33_io_output : _T_12552; // @[Mux.scala 31:69:@57021.4]
  assign _T_12538 = RetimeWrapper_415_io_out; // @[package.scala 96:25:@56985.4 package.scala 96:25:@56986.4]
  assign _T_12554 = _T_12538 ? Mem1D_31_io_output : _T_12553; // @[Mux.scala 31:69:@57022.4]
  assign _T_12535 = RetimeWrapper_414_io_out; // @[package.scala 96:25:@56977.4 package.scala 96:25:@56978.4]
  assign _T_12555 = _T_12535 ? Mem1D_29_io_output : _T_12554; // @[Mux.scala 31:69:@57023.4]
  assign _T_12532 = RetimeWrapper_413_io_out; // @[package.scala 96:25:@56969.4 package.scala 96:25:@56970.4]
  assign _T_12556 = _T_12532 ? Mem1D_27_io_output : _T_12555; // @[Mux.scala 31:69:@57024.4]
  assign _T_12529 = RetimeWrapper_412_io_out; // @[package.scala 96:25:@56961.4 package.scala 96:25:@56962.4]
  assign _T_12557 = _T_12529 ? Mem1D_25_io_output : _T_12556; // @[Mux.scala 31:69:@57025.4]
  assign _T_12526 = RetimeWrapper_411_io_out; // @[package.scala 96:25:@56953.4 package.scala 96:25:@56954.4]
  assign _T_12558 = _T_12526 ? Mem1D_23_io_output : _T_12557; // @[Mux.scala 31:69:@57026.4]
  assign _T_12523 = RetimeWrapper_410_io_out; // @[package.scala 96:25:@56945.4 package.scala 96:25:@56946.4]
  assign _T_12559 = _T_12523 ? Mem1D_21_io_output : _T_12558; // @[Mux.scala 31:69:@57027.4]
  assign _T_12520 = RetimeWrapper_409_io_out; // @[package.scala 96:25:@56937.4 package.scala 96:25:@56938.4]
  assign _T_12560 = _T_12520 ? Mem1D_19_io_output : _T_12559; // @[Mux.scala 31:69:@57028.4]
  assign _T_12517 = RetimeWrapper_408_io_out; // @[package.scala 96:25:@56929.4 package.scala 96:25:@56930.4]
  assign _T_12561 = _T_12517 ? Mem1D_17_io_output : _T_12560; // @[Mux.scala 31:69:@57029.4]
  assign _T_12514 = RetimeWrapper_407_io_out; // @[package.scala 96:25:@56921.4 package.scala 96:25:@56922.4]
  assign _T_12562 = _T_12514 ? Mem1D_15_io_output : _T_12561; // @[Mux.scala 31:69:@57030.4]
  assign _T_12511 = RetimeWrapper_406_io_out; // @[package.scala 96:25:@56913.4 package.scala 96:25:@56914.4]
  assign _T_12563 = _T_12511 ? Mem1D_13_io_output : _T_12562; // @[Mux.scala 31:69:@57031.4]
  assign _T_12508 = RetimeWrapper_405_io_out; // @[package.scala 96:25:@56905.4 package.scala 96:25:@56906.4]
  assign _T_12564 = _T_12508 ? Mem1D_11_io_output : _T_12563; // @[Mux.scala 31:69:@57032.4]
  assign _T_12505 = RetimeWrapper_404_io_out; // @[package.scala 96:25:@56897.4 package.scala 96:25:@56898.4]
  assign _T_12565 = _T_12505 ? Mem1D_9_io_output : _T_12564; // @[Mux.scala 31:69:@57033.4]
  assign _T_12502 = RetimeWrapper_403_io_out; // @[package.scala 96:25:@56889.4 package.scala 96:25:@56890.4]
  assign _T_12566 = _T_12502 ? Mem1D_7_io_output : _T_12565; // @[Mux.scala 31:69:@57034.4]
  assign _T_12499 = RetimeWrapper_402_io_out; // @[package.scala 96:25:@56881.4 package.scala 96:25:@56882.4]
  assign _T_12567 = _T_12499 ? Mem1D_5_io_output : _T_12566; // @[Mux.scala 31:69:@57035.4]
  assign _T_12496 = RetimeWrapper_401_io_out; // @[package.scala 96:25:@56873.4 package.scala 96:25:@56874.4]
  assign _T_12568 = _T_12496 ? Mem1D_3_io_output : _T_12567; // @[Mux.scala 31:69:@57036.4]
  assign _T_12493 = RetimeWrapper_400_io_out; // @[package.scala 96:25:@56865.4 package.scala 96:25:@56866.4]
  assign _T_12726 = RetimeWrapper_438_io_out; // @[package.scala 96:25:@57249.4 package.scala 96:25:@57250.4]
  assign _T_12730 = _T_12726 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@57259.4]
  assign _T_12723 = RetimeWrapper_437_io_out; // @[package.scala 96:25:@57241.4 package.scala 96:25:@57242.4]
  assign _T_12731 = _T_12723 ? Mem1D_35_io_output : _T_12730; // @[Mux.scala 31:69:@57260.4]
  assign _T_12720 = RetimeWrapper_436_io_out; // @[package.scala 96:25:@57233.4 package.scala 96:25:@57234.4]
  assign _T_12732 = _T_12720 ? Mem1D_33_io_output : _T_12731; // @[Mux.scala 31:69:@57261.4]
  assign _T_12717 = RetimeWrapper_435_io_out; // @[package.scala 96:25:@57225.4 package.scala 96:25:@57226.4]
  assign _T_12733 = _T_12717 ? Mem1D_31_io_output : _T_12732; // @[Mux.scala 31:69:@57262.4]
  assign _T_12714 = RetimeWrapper_434_io_out; // @[package.scala 96:25:@57217.4 package.scala 96:25:@57218.4]
  assign _T_12734 = _T_12714 ? Mem1D_29_io_output : _T_12733; // @[Mux.scala 31:69:@57263.4]
  assign _T_12711 = RetimeWrapper_433_io_out; // @[package.scala 96:25:@57209.4 package.scala 96:25:@57210.4]
  assign _T_12735 = _T_12711 ? Mem1D_27_io_output : _T_12734; // @[Mux.scala 31:69:@57264.4]
  assign _T_12708 = RetimeWrapper_432_io_out; // @[package.scala 96:25:@57201.4 package.scala 96:25:@57202.4]
  assign _T_12736 = _T_12708 ? Mem1D_25_io_output : _T_12735; // @[Mux.scala 31:69:@57265.4]
  assign _T_12705 = RetimeWrapper_431_io_out; // @[package.scala 96:25:@57193.4 package.scala 96:25:@57194.4]
  assign _T_12737 = _T_12705 ? Mem1D_23_io_output : _T_12736; // @[Mux.scala 31:69:@57266.4]
  assign _T_12702 = RetimeWrapper_430_io_out; // @[package.scala 96:25:@57185.4 package.scala 96:25:@57186.4]
  assign _T_12738 = _T_12702 ? Mem1D_21_io_output : _T_12737; // @[Mux.scala 31:69:@57267.4]
  assign _T_12699 = RetimeWrapper_429_io_out; // @[package.scala 96:25:@57177.4 package.scala 96:25:@57178.4]
  assign _T_12739 = _T_12699 ? Mem1D_19_io_output : _T_12738; // @[Mux.scala 31:69:@57268.4]
  assign _T_12696 = RetimeWrapper_428_io_out; // @[package.scala 96:25:@57169.4 package.scala 96:25:@57170.4]
  assign _T_12740 = _T_12696 ? Mem1D_17_io_output : _T_12739; // @[Mux.scala 31:69:@57269.4]
  assign _T_12693 = RetimeWrapper_427_io_out; // @[package.scala 96:25:@57161.4 package.scala 96:25:@57162.4]
  assign _T_12741 = _T_12693 ? Mem1D_15_io_output : _T_12740; // @[Mux.scala 31:69:@57270.4]
  assign _T_12690 = RetimeWrapper_426_io_out; // @[package.scala 96:25:@57153.4 package.scala 96:25:@57154.4]
  assign _T_12742 = _T_12690 ? Mem1D_13_io_output : _T_12741; // @[Mux.scala 31:69:@57271.4]
  assign _T_12687 = RetimeWrapper_425_io_out; // @[package.scala 96:25:@57145.4 package.scala 96:25:@57146.4]
  assign _T_12743 = _T_12687 ? Mem1D_11_io_output : _T_12742; // @[Mux.scala 31:69:@57272.4]
  assign _T_12684 = RetimeWrapper_424_io_out; // @[package.scala 96:25:@57137.4 package.scala 96:25:@57138.4]
  assign _T_12744 = _T_12684 ? Mem1D_9_io_output : _T_12743; // @[Mux.scala 31:69:@57273.4]
  assign _T_12681 = RetimeWrapper_423_io_out; // @[package.scala 96:25:@57129.4 package.scala 96:25:@57130.4]
  assign _T_12745 = _T_12681 ? Mem1D_7_io_output : _T_12744; // @[Mux.scala 31:69:@57274.4]
  assign _T_12678 = RetimeWrapper_422_io_out; // @[package.scala 96:25:@57121.4 package.scala 96:25:@57122.4]
  assign _T_12746 = _T_12678 ? Mem1D_5_io_output : _T_12745; // @[Mux.scala 31:69:@57275.4]
  assign _T_12675 = RetimeWrapper_421_io_out; // @[package.scala 96:25:@57113.4 package.scala 96:25:@57114.4]
  assign _T_12747 = _T_12675 ? Mem1D_3_io_output : _T_12746; // @[Mux.scala 31:69:@57276.4]
  assign _T_12672 = RetimeWrapper_420_io_out; // @[package.scala 96:25:@57105.4 package.scala 96:25:@57106.4]
  assign _T_12905 = RetimeWrapper_458_io_out; // @[package.scala 96:25:@57489.4 package.scala 96:25:@57490.4]
  assign _T_12909 = _T_12905 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@57499.4]
  assign _T_12902 = RetimeWrapper_457_io_out; // @[package.scala 96:25:@57481.4 package.scala 96:25:@57482.4]
  assign _T_12910 = _T_12902 ? Mem1D_34_io_output : _T_12909; // @[Mux.scala 31:69:@57500.4]
  assign _T_12899 = RetimeWrapper_456_io_out; // @[package.scala 96:25:@57473.4 package.scala 96:25:@57474.4]
  assign _T_12911 = _T_12899 ? Mem1D_32_io_output : _T_12910; // @[Mux.scala 31:69:@57501.4]
  assign _T_12896 = RetimeWrapper_455_io_out; // @[package.scala 96:25:@57465.4 package.scala 96:25:@57466.4]
  assign _T_12912 = _T_12896 ? Mem1D_30_io_output : _T_12911; // @[Mux.scala 31:69:@57502.4]
  assign _T_12893 = RetimeWrapper_454_io_out; // @[package.scala 96:25:@57457.4 package.scala 96:25:@57458.4]
  assign _T_12913 = _T_12893 ? Mem1D_28_io_output : _T_12912; // @[Mux.scala 31:69:@57503.4]
  assign _T_12890 = RetimeWrapper_453_io_out; // @[package.scala 96:25:@57449.4 package.scala 96:25:@57450.4]
  assign _T_12914 = _T_12890 ? Mem1D_26_io_output : _T_12913; // @[Mux.scala 31:69:@57504.4]
  assign _T_12887 = RetimeWrapper_452_io_out; // @[package.scala 96:25:@57441.4 package.scala 96:25:@57442.4]
  assign _T_12915 = _T_12887 ? Mem1D_24_io_output : _T_12914; // @[Mux.scala 31:69:@57505.4]
  assign _T_12884 = RetimeWrapper_451_io_out; // @[package.scala 96:25:@57433.4 package.scala 96:25:@57434.4]
  assign _T_12916 = _T_12884 ? Mem1D_22_io_output : _T_12915; // @[Mux.scala 31:69:@57506.4]
  assign _T_12881 = RetimeWrapper_450_io_out; // @[package.scala 96:25:@57425.4 package.scala 96:25:@57426.4]
  assign _T_12917 = _T_12881 ? Mem1D_20_io_output : _T_12916; // @[Mux.scala 31:69:@57507.4]
  assign _T_12878 = RetimeWrapper_449_io_out; // @[package.scala 96:25:@57417.4 package.scala 96:25:@57418.4]
  assign _T_12918 = _T_12878 ? Mem1D_18_io_output : _T_12917; // @[Mux.scala 31:69:@57508.4]
  assign _T_12875 = RetimeWrapper_448_io_out; // @[package.scala 96:25:@57409.4 package.scala 96:25:@57410.4]
  assign _T_12919 = _T_12875 ? Mem1D_16_io_output : _T_12918; // @[Mux.scala 31:69:@57509.4]
  assign _T_12872 = RetimeWrapper_447_io_out; // @[package.scala 96:25:@57401.4 package.scala 96:25:@57402.4]
  assign _T_12920 = _T_12872 ? Mem1D_14_io_output : _T_12919; // @[Mux.scala 31:69:@57510.4]
  assign _T_12869 = RetimeWrapper_446_io_out; // @[package.scala 96:25:@57393.4 package.scala 96:25:@57394.4]
  assign _T_12921 = _T_12869 ? Mem1D_12_io_output : _T_12920; // @[Mux.scala 31:69:@57511.4]
  assign _T_12866 = RetimeWrapper_445_io_out; // @[package.scala 96:25:@57385.4 package.scala 96:25:@57386.4]
  assign _T_12922 = _T_12866 ? Mem1D_10_io_output : _T_12921; // @[Mux.scala 31:69:@57512.4]
  assign _T_12863 = RetimeWrapper_444_io_out; // @[package.scala 96:25:@57377.4 package.scala 96:25:@57378.4]
  assign _T_12923 = _T_12863 ? Mem1D_8_io_output : _T_12922; // @[Mux.scala 31:69:@57513.4]
  assign _T_12860 = RetimeWrapper_443_io_out; // @[package.scala 96:25:@57369.4 package.scala 96:25:@57370.4]
  assign _T_12924 = _T_12860 ? Mem1D_6_io_output : _T_12923; // @[Mux.scala 31:69:@57514.4]
  assign _T_12857 = RetimeWrapper_442_io_out; // @[package.scala 96:25:@57361.4 package.scala 96:25:@57362.4]
  assign _T_12925 = _T_12857 ? Mem1D_4_io_output : _T_12924; // @[Mux.scala 31:69:@57515.4]
  assign _T_12854 = RetimeWrapper_441_io_out; // @[package.scala 96:25:@57353.4 package.scala 96:25:@57354.4]
  assign _T_12926 = _T_12854 ? Mem1D_2_io_output : _T_12925; // @[Mux.scala 31:69:@57516.4]
  assign _T_12851 = RetimeWrapper_440_io_out; // @[package.scala 96:25:@57345.4 package.scala 96:25:@57346.4]
  assign _T_13084 = RetimeWrapper_478_io_out; // @[package.scala 96:25:@57729.4 package.scala 96:25:@57730.4]
  assign _T_13088 = _T_13084 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@57739.4]
  assign _T_13081 = RetimeWrapper_477_io_out; // @[package.scala 96:25:@57721.4 package.scala 96:25:@57722.4]
  assign _T_13089 = _T_13081 ? Mem1D_35_io_output : _T_13088; // @[Mux.scala 31:69:@57740.4]
  assign _T_13078 = RetimeWrapper_476_io_out; // @[package.scala 96:25:@57713.4 package.scala 96:25:@57714.4]
  assign _T_13090 = _T_13078 ? Mem1D_33_io_output : _T_13089; // @[Mux.scala 31:69:@57741.4]
  assign _T_13075 = RetimeWrapper_475_io_out; // @[package.scala 96:25:@57705.4 package.scala 96:25:@57706.4]
  assign _T_13091 = _T_13075 ? Mem1D_31_io_output : _T_13090; // @[Mux.scala 31:69:@57742.4]
  assign _T_13072 = RetimeWrapper_474_io_out; // @[package.scala 96:25:@57697.4 package.scala 96:25:@57698.4]
  assign _T_13092 = _T_13072 ? Mem1D_29_io_output : _T_13091; // @[Mux.scala 31:69:@57743.4]
  assign _T_13069 = RetimeWrapper_473_io_out; // @[package.scala 96:25:@57689.4 package.scala 96:25:@57690.4]
  assign _T_13093 = _T_13069 ? Mem1D_27_io_output : _T_13092; // @[Mux.scala 31:69:@57744.4]
  assign _T_13066 = RetimeWrapper_472_io_out; // @[package.scala 96:25:@57681.4 package.scala 96:25:@57682.4]
  assign _T_13094 = _T_13066 ? Mem1D_25_io_output : _T_13093; // @[Mux.scala 31:69:@57745.4]
  assign _T_13063 = RetimeWrapper_471_io_out; // @[package.scala 96:25:@57673.4 package.scala 96:25:@57674.4]
  assign _T_13095 = _T_13063 ? Mem1D_23_io_output : _T_13094; // @[Mux.scala 31:69:@57746.4]
  assign _T_13060 = RetimeWrapper_470_io_out; // @[package.scala 96:25:@57665.4 package.scala 96:25:@57666.4]
  assign _T_13096 = _T_13060 ? Mem1D_21_io_output : _T_13095; // @[Mux.scala 31:69:@57747.4]
  assign _T_13057 = RetimeWrapper_469_io_out; // @[package.scala 96:25:@57657.4 package.scala 96:25:@57658.4]
  assign _T_13097 = _T_13057 ? Mem1D_19_io_output : _T_13096; // @[Mux.scala 31:69:@57748.4]
  assign _T_13054 = RetimeWrapper_468_io_out; // @[package.scala 96:25:@57649.4 package.scala 96:25:@57650.4]
  assign _T_13098 = _T_13054 ? Mem1D_17_io_output : _T_13097; // @[Mux.scala 31:69:@57749.4]
  assign _T_13051 = RetimeWrapper_467_io_out; // @[package.scala 96:25:@57641.4 package.scala 96:25:@57642.4]
  assign _T_13099 = _T_13051 ? Mem1D_15_io_output : _T_13098; // @[Mux.scala 31:69:@57750.4]
  assign _T_13048 = RetimeWrapper_466_io_out; // @[package.scala 96:25:@57633.4 package.scala 96:25:@57634.4]
  assign _T_13100 = _T_13048 ? Mem1D_13_io_output : _T_13099; // @[Mux.scala 31:69:@57751.4]
  assign _T_13045 = RetimeWrapper_465_io_out; // @[package.scala 96:25:@57625.4 package.scala 96:25:@57626.4]
  assign _T_13101 = _T_13045 ? Mem1D_11_io_output : _T_13100; // @[Mux.scala 31:69:@57752.4]
  assign _T_13042 = RetimeWrapper_464_io_out; // @[package.scala 96:25:@57617.4 package.scala 96:25:@57618.4]
  assign _T_13102 = _T_13042 ? Mem1D_9_io_output : _T_13101; // @[Mux.scala 31:69:@57753.4]
  assign _T_13039 = RetimeWrapper_463_io_out; // @[package.scala 96:25:@57609.4 package.scala 96:25:@57610.4]
  assign _T_13103 = _T_13039 ? Mem1D_7_io_output : _T_13102; // @[Mux.scala 31:69:@57754.4]
  assign _T_13036 = RetimeWrapper_462_io_out; // @[package.scala 96:25:@57601.4 package.scala 96:25:@57602.4]
  assign _T_13104 = _T_13036 ? Mem1D_5_io_output : _T_13103; // @[Mux.scala 31:69:@57755.4]
  assign _T_13033 = RetimeWrapper_461_io_out; // @[package.scala 96:25:@57593.4 package.scala 96:25:@57594.4]
  assign _T_13105 = _T_13033 ? Mem1D_3_io_output : _T_13104; // @[Mux.scala 31:69:@57756.4]
  assign _T_13030 = RetimeWrapper_460_io_out; // @[package.scala 96:25:@57585.4 package.scala 96:25:@57586.4]
  assign _T_13263 = RetimeWrapper_498_io_out; // @[package.scala 96:25:@57969.4 package.scala 96:25:@57970.4]
  assign _T_13267 = _T_13263 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@57979.4]
  assign _T_13260 = RetimeWrapper_497_io_out; // @[package.scala 96:25:@57961.4 package.scala 96:25:@57962.4]
  assign _T_13268 = _T_13260 ? Mem1D_35_io_output : _T_13267; // @[Mux.scala 31:69:@57980.4]
  assign _T_13257 = RetimeWrapper_496_io_out; // @[package.scala 96:25:@57953.4 package.scala 96:25:@57954.4]
  assign _T_13269 = _T_13257 ? Mem1D_33_io_output : _T_13268; // @[Mux.scala 31:69:@57981.4]
  assign _T_13254 = RetimeWrapper_495_io_out; // @[package.scala 96:25:@57945.4 package.scala 96:25:@57946.4]
  assign _T_13270 = _T_13254 ? Mem1D_31_io_output : _T_13269; // @[Mux.scala 31:69:@57982.4]
  assign _T_13251 = RetimeWrapper_494_io_out; // @[package.scala 96:25:@57937.4 package.scala 96:25:@57938.4]
  assign _T_13271 = _T_13251 ? Mem1D_29_io_output : _T_13270; // @[Mux.scala 31:69:@57983.4]
  assign _T_13248 = RetimeWrapper_493_io_out; // @[package.scala 96:25:@57929.4 package.scala 96:25:@57930.4]
  assign _T_13272 = _T_13248 ? Mem1D_27_io_output : _T_13271; // @[Mux.scala 31:69:@57984.4]
  assign _T_13245 = RetimeWrapper_492_io_out; // @[package.scala 96:25:@57921.4 package.scala 96:25:@57922.4]
  assign _T_13273 = _T_13245 ? Mem1D_25_io_output : _T_13272; // @[Mux.scala 31:69:@57985.4]
  assign _T_13242 = RetimeWrapper_491_io_out; // @[package.scala 96:25:@57913.4 package.scala 96:25:@57914.4]
  assign _T_13274 = _T_13242 ? Mem1D_23_io_output : _T_13273; // @[Mux.scala 31:69:@57986.4]
  assign _T_13239 = RetimeWrapper_490_io_out; // @[package.scala 96:25:@57905.4 package.scala 96:25:@57906.4]
  assign _T_13275 = _T_13239 ? Mem1D_21_io_output : _T_13274; // @[Mux.scala 31:69:@57987.4]
  assign _T_13236 = RetimeWrapper_489_io_out; // @[package.scala 96:25:@57897.4 package.scala 96:25:@57898.4]
  assign _T_13276 = _T_13236 ? Mem1D_19_io_output : _T_13275; // @[Mux.scala 31:69:@57988.4]
  assign _T_13233 = RetimeWrapper_488_io_out; // @[package.scala 96:25:@57889.4 package.scala 96:25:@57890.4]
  assign _T_13277 = _T_13233 ? Mem1D_17_io_output : _T_13276; // @[Mux.scala 31:69:@57989.4]
  assign _T_13230 = RetimeWrapper_487_io_out; // @[package.scala 96:25:@57881.4 package.scala 96:25:@57882.4]
  assign _T_13278 = _T_13230 ? Mem1D_15_io_output : _T_13277; // @[Mux.scala 31:69:@57990.4]
  assign _T_13227 = RetimeWrapper_486_io_out; // @[package.scala 96:25:@57873.4 package.scala 96:25:@57874.4]
  assign _T_13279 = _T_13227 ? Mem1D_13_io_output : _T_13278; // @[Mux.scala 31:69:@57991.4]
  assign _T_13224 = RetimeWrapper_485_io_out; // @[package.scala 96:25:@57865.4 package.scala 96:25:@57866.4]
  assign _T_13280 = _T_13224 ? Mem1D_11_io_output : _T_13279; // @[Mux.scala 31:69:@57992.4]
  assign _T_13221 = RetimeWrapper_484_io_out; // @[package.scala 96:25:@57857.4 package.scala 96:25:@57858.4]
  assign _T_13281 = _T_13221 ? Mem1D_9_io_output : _T_13280; // @[Mux.scala 31:69:@57993.4]
  assign _T_13218 = RetimeWrapper_483_io_out; // @[package.scala 96:25:@57849.4 package.scala 96:25:@57850.4]
  assign _T_13282 = _T_13218 ? Mem1D_7_io_output : _T_13281; // @[Mux.scala 31:69:@57994.4]
  assign _T_13215 = RetimeWrapper_482_io_out; // @[package.scala 96:25:@57841.4 package.scala 96:25:@57842.4]
  assign _T_13283 = _T_13215 ? Mem1D_5_io_output : _T_13282; // @[Mux.scala 31:69:@57995.4]
  assign _T_13212 = RetimeWrapper_481_io_out; // @[package.scala 96:25:@57833.4 package.scala 96:25:@57834.4]
  assign _T_13284 = _T_13212 ? Mem1D_3_io_output : _T_13283; // @[Mux.scala 31:69:@57996.4]
  assign _T_13209 = RetimeWrapper_480_io_out; // @[package.scala 96:25:@57825.4 package.scala 96:25:@57826.4]
  assign _T_13442 = RetimeWrapper_518_io_out; // @[package.scala 96:25:@58209.4 package.scala 96:25:@58210.4]
  assign _T_13446 = _T_13442 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@58219.4]
  assign _T_13439 = RetimeWrapper_517_io_out; // @[package.scala 96:25:@58201.4 package.scala 96:25:@58202.4]
  assign _T_13447 = _T_13439 ? Mem1D_35_io_output : _T_13446; // @[Mux.scala 31:69:@58220.4]
  assign _T_13436 = RetimeWrapper_516_io_out; // @[package.scala 96:25:@58193.4 package.scala 96:25:@58194.4]
  assign _T_13448 = _T_13436 ? Mem1D_33_io_output : _T_13447; // @[Mux.scala 31:69:@58221.4]
  assign _T_13433 = RetimeWrapper_515_io_out; // @[package.scala 96:25:@58185.4 package.scala 96:25:@58186.4]
  assign _T_13449 = _T_13433 ? Mem1D_31_io_output : _T_13448; // @[Mux.scala 31:69:@58222.4]
  assign _T_13430 = RetimeWrapper_514_io_out; // @[package.scala 96:25:@58177.4 package.scala 96:25:@58178.4]
  assign _T_13450 = _T_13430 ? Mem1D_29_io_output : _T_13449; // @[Mux.scala 31:69:@58223.4]
  assign _T_13427 = RetimeWrapper_513_io_out; // @[package.scala 96:25:@58169.4 package.scala 96:25:@58170.4]
  assign _T_13451 = _T_13427 ? Mem1D_27_io_output : _T_13450; // @[Mux.scala 31:69:@58224.4]
  assign _T_13424 = RetimeWrapper_512_io_out; // @[package.scala 96:25:@58161.4 package.scala 96:25:@58162.4]
  assign _T_13452 = _T_13424 ? Mem1D_25_io_output : _T_13451; // @[Mux.scala 31:69:@58225.4]
  assign _T_13421 = RetimeWrapper_511_io_out; // @[package.scala 96:25:@58153.4 package.scala 96:25:@58154.4]
  assign _T_13453 = _T_13421 ? Mem1D_23_io_output : _T_13452; // @[Mux.scala 31:69:@58226.4]
  assign _T_13418 = RetimeWrapper_510_io_out; // @[package.scala 96:25:@58145.4 package.scala 96:25:@58146.4]
  assign _T_13454 = _T_13418 ? Mem1D_21_io_output : _T_13453; // @[Mux.scala 31:69:@58227.4]
  assign _T_13415 = RetimeWrapper_509_io_out; // @[package.scala 96:25:@58137.4 package.scala 96:25:@58138.4]
  assign _T_13455 = _T_13415 ? Mem1D_19_io_output : _T_13454; // @[Mux.scala 31:69:@58228.4]
  assign _T_13412 = RetimeWrapper_508_io_out; // @[package.scala 96:25:@58129.4 package.scala 96:25:@58130.4]
  assign _T_13456 = _T_13412 ? Mem1D_17_io_output : _T_13455; // @[Mux.scala 31:69:@58229.4]
  assign _T_13409 = RetimeWrapper_507_io_out; // @[package.scala 96:25:@58121.4 package.scala 96:25:@58122.4]
  assign _T_13457 = _T_13409 ? Mem1D_15_io_output : _T_13456; // @[Mux.scala 31:69:@58230.4]
  assign _T_13406 = RetimeWrapper_506_io_out; // @[package.scala 96:25:@58113.4 package.scala 96:25:@58114.4]
  assign _T_13458 = _T_13406 ? Mem1D_13_io_output : _T_13457; // @[Mux.scala 31:69:@58231.4]
  assign _T_13403 = RetimeWrapper_505_io_out; // @[package.scala 96:25:@58105.4 package.scala 96:25:@58106.4]
  assign _T_13459 = _T_13403 ? Mem1D_11_io_output : _T_13458; // @[Mux.scala 31:69:@58232.4]
  assign _T_13400 = RetimeWrapper_504_io_out; // @[package.scala 96:25:@58097.4 package.scala 96:25:@58098.4]
  assign _T_13460 = _T_13400 ? Mem1D_9_io_output : _T_13459; // @[Mux.scala 31:69:@58233.4]
  assign _T_13397 = RetimeWrapper_503_io_out; // @[package.scala 96:25:@58089.4 package.scala 96:25:@58090.4]
  assign _T_13461 = _T_13397 ? Mem1D_7_io_output : _T_13460; // @[Mux.scala 31:69:@58234.4]
  assign _T_13394 = RetimeWrapper_502_io_out; // @[package.scala 96:25:@58081.4 package.scala 96:25:@58082.4]
  assign _T_13462 = _T_13394 ? Mem1D_5_io_output : _T_13461; // @[Mux.scala 31:69:@58235.4]
  assign _T_13391 = RetimeWrapper_501_io_out; // @[package.scala 96:25:@58073.4 package.scala 96:25:@58074.4]
  assign _T_13463 = _T_13391 ? Mem1D_3_io_output : _T_13462; // @[Mux.scala 31:69:@58236.4]
  assign _T_13388 = RetimeWrapper_500_io_out; // @[package.scala 96:25:@58065.4 package.scala 96:25:@58066.4]
  assign _T_13621 = RetimeWrapper_538_io_out; // @[package.scala 96:25:@58449.4 package.scala 96:25:@58450.4]
  assign _T_13625 = _T_13621 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@58459.4]
  assign _T_13618 = RetimeWrapper_537_io_out; // @[package.scala 96:25:@58441.4 package.scala 96:25:@58442.4]
  assign _T_13626 = _T_13618 ? Mem1D_34_io_output : _T_13625; // @[Mux.scala 31:69:@58460.4]
  assign _T_13615 = RetimeWrapper_536_io_out; // @[package.scala 96:25:@58433.4 package.scala 96:25:@58434.4]
  assign _T_13627 = _T_13615 ? Mem1D_32_io_output : _T_13626; // @[Mux.scala 31:69:@58461.4]
  assign _T_13612 = RetimeWrapper_535_io_out; // @[package.scala 96:25:@58425.4 package.scala 96:25:@58426.4]
  assign _T_13628 = _T_13612 ? Mem1D_30_io_output : _T_13627; // @[Mux.scala 31:69:@58462.4]
  assign _T_13609 = RetimeWrapper_534_io_out; // @[package.scala 96:25:@58417.4 package.scala 96:25:@58418.4]
  assign _T_13629 = _T_13609 ? Mem1D_28_io_output : _T_13628; // @[Mux.scala 31:69:@58463.4]
  assign _T_13606 = RetimeWrapper_533_io_out; // @[package.scala 96:25:@58409.4 package.scala 96:25:@58410.4]
  assign _T_13630 = _T_13606 ? Mem1D_26_io_output : _T_13629; // @[Mux.scala 31:69:@58464.4]
  assign _T_13603 = RetimeWrapper_532_io_out; // @[package.scala 96:25:@58401.4 package.scala 96:25:@58402.4]
  assign _T_13631 = _T_13603 ? Mem1D_24_io_output : _T_13630; // @[Mux.scala 31:69:@58465.4]
  assign _T_13600 = RetimeWrapper_531_io_out; // @[package.scala 96:25:@58393.4 package.scala 96:25:@58394.4]
  assign _T_13632 = _T_13600 ? Mem1D_22_io_output : _T_13631; // @[Mux.scala 31:69:@58466.4]
  assign _T_13597 = RetimeWrapper_530_io_out; // @[package.scala 96:25:@58385.4 package.scala 96:25:@58386.4]
  assign _T_13633 = _T_13597 ? Mem1D_20_io_output : _T_13632; // @[Mux.scala 31:69:@58467.4]
  assign _T_13594 = RetimeWrapper_529_io_out; // @[package.scala 96:25:@58377.4 package.scala 96:25:@58378.4]
  assign _T_13634 = _T_13594 ? Mem1D_18_io_output : _T_13633; // @[Mux.scala 31:69:@58468.4]
  assign _T_13591 = RetimeWrapper_528_io_out; // @[package.scala 96:25:@58369.4 package.scala 96:25:@58370.4]
  assign _T_13635 = _T_13591 ? Mem1D_16_io_output : _T_13634; // @[Mux.scala 31:69:@58469.4]
  assign _T_13588 = RetimeWrapper_527_io_out; // @[package.scala 96:25:@58361.4 package.scala 96:25:@58362.4]
  assign _T_13636 = _T_13588 ? Mem1D_14_io_output : _T_13635; // @[Mux.scala 31:69:@58470.4]
  assign _T_13585 = RetimeWrapper_526_io_out; // @[package.scala 96:25:@58353.4 package.scala 96:25:@58354.4]
  assign _T_13637 = _T_13585 ? Mem1D_12_io_output : _T_13636; // @[Mux.scala 31:69:@58471.4]
  assign _T_13582 = RetimeWrapper_525_io_out; // @[package.scala 96:25:@58345.4 package.scala 96:25:@58346.4]
  assign _T_13638 = _T_13582 ? Mem1D_10_io_output : _T_13637; // @[Mux.scala 31:69:@58472.4]
  assign _T_13579 = RetimeWrapper_524_io_out; // @[package.scala 96:25:@58337.4 package.scala 96:25:@58338.4]
  assign _T_13639 = _T_13579 ? Mem1D_8_io_output : _T_13638; // @[Mux.scala 31:69:@58473.4]
  assign _T_13576 = RetimeWrapper_523_io_out; // @[package.scala 96:25:@58329.4 package.scala 96:25:@58330.4]
  assign _T_13640 = _T_13576 ? Mem1D_6_io_output : _T_13639; // @[Mux.scala 31:69:@58474.4]
  assign _T_13573 = RetimeWrapper_522_io_out; // @[package.scala 96:25:@58321.4 package.scala 96:25:@58322.4]
  assign _T_13641 = _T_13573 ? Mem1D_4_io_output : _T_13640; // @[Mux.scala 31:69:@58475.4]
  assign _T_13570 = RetimeWrapper_521_io_out; // @[package.scala 96:25:@58313.4 package.scala 96:25:@58314.4]
  assign _T_13642 = _T_13570 ? Mem1D_2_io_output : _T_13641; // @[Mux.scala 31:69:@58476.4]
  assign _T_13567 = RetimeWrapper_520_io_out; // @[package.scala 96:25:@58305.4 package.scala 96:25:@58306.4]
  assign _T_13800 = RetimeWrapper_558_io_out; // @[package.scala 96:25:@58689.4 package.scala 96:25:@58690.4]
  assign _T_13804 = _T_13800 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@58699.4]
  assign _T_13797 = RetimeWrapper_557_io_out; // @[package.scala 96:25:@58681.4 package.scala 96:25:@58682.4]
  assign _T_13805 = _T_13797 ? Mem1D_35_io_output : _T_13804; // @[Mux.scala 31:69:@58700.4]
  assign _T_13794 = RetimeWrapper_556_io_out; // @[package.scala 96:25:@58673.4 package.scala 96:25:@58674.4]
  assign _T_13806 = _T_13794 ? Mem1D_33_io_output : _T_13805; // @[Mux.scala 31:69:@58701.4]
  assign _T_13791 = RetimeWrapper_555_io_out; // @[package.scala 96:25:@58665.4 package.scala 96:25:@58666.4]
  assign _T_13807 = _T_13791 ? Mem1D_31_io_output : _T_13806; // @[Mux.scala 31:69:@58702.4]
  assign _T_13788 = RetimeWrapper_554_io_out; // @[package.scala 96:25:@58657.4 package.scala 96:25:@58658.4]
  assign _T_13808 = _T_13788 ? Mem1D_29_io_output : _T_13807; // @[Mux.scala 31:69:@58703.4]
  assign _T_13785 = RetimeWrapper_553_io_out; // @[package.scala 96:25:@58649.4 package.scala 96:25:@58650.4]
  assign _T_13809 = _T_13785 ? Mem1D_27_io_output : _T_13808; // @[Mux.scala 31:69:@58704.4]
  assign _T_13782 = RetimeWrapper_552_io_out; // @[package.scala 96:25:@58641.4 package.scala 96:25:@58642.4]
  assign _T_13810 = _T_13782 ? Mem1D_25_io_output : _T_13809; // @[Mux.scala 31:69:@58705.4]
  assign _T_13779 = RetimeWrapper_551_io_out; // @[package.scala 96:25:@58633.4 package.scala 96:25:@58634.4]
  assign _T_13811 = _T_13779 ? Mem1D_23_io_output : _T_13810; // @[Mux.scala 31:69:@58706.4]
  assign _T_13776 = RetimeWrapper_550_io_out; // @[package.scala 96:25:@58625.4 package.scala 96:25:@58626.4]
  assign _T_13812 = _T_13776 ? Mem1D_21_io_output : _T_13811; // @[Mux.scala 31:69:@58707.4]
  assign _T_13773 = RetimeWrapper_549_io_out; // @[package.scala 96:25:@58617.4 package.scala 96:25:@58618.4]
  assign _T_13813 = _T_13773 ? Mem1D_19_io_output : _T_13812; // @[Mux.scala 31:69:@58708.4]
  assign _T_13770 = RetimeWrapper_548_io_out; // @[package.scala 96:25:@58609.4 package.scala 96:25:@58610.4]
  assign _T_13814 = _T_13770 ? Mem1D_17_io_output : _T_13813; // @[Mux.scala 31:69:@58709.4]
  assign _T_13767 = RetimeWrapper_547_io_out; // @[package.scala 96:25:@58601.4 package.scala 96:25:@58602.4]
  assign _T_13815 = _T_13767 ? Mem1D_15_io_output : _T_13814; // @[Mux.scala 31:69:@58710.4]
  assign _T_13764 = RetimeWrapper_546_io_out; // @[package.scala 96:25:@58593.4 package.scala 96:25:@58594.4]
  assign _T_13816 = _T_13764 ? Mem1D_13_io_output : _T_13815; // @[Mux.scala 31:69:@58711.4]
  assign _T_13761 = RetimeWrapper_545_io_out; // @[package.scala 96:25:@58585.4 package.scala 96:25:@58586.4]
  assign _T_13817 = _T_13761 ? Mem1D_11_io_output : _T_13816; // @[Mux.scala 31:69:@58712.4]
  assign _T_13758 = RetimeWrapper_544_io_out; // @[package.scala 96:25:@58577.4 package.scala 96:25:@58578.4]
  assign _T_13818 = _T_13758 ? Mem1D_9_io_output : _T_13817; // @[Mux.scala 31:69:@58713.4]
  assign _T_13755 = RetimeWrapper_543_io_out; // @[package.scala 96:25:@58569.4 package.scala 96:25:@58570.4]
  assign _T_13819 = _T_13755 ? Mem1D_7_io_output : _T_13818; // @[Mux.scala 31:69:@58714.4]
  assign _T_13752 = RetimeWrapper_542_io_out; // @[package.scala 96:25:@58561.4 package.scala 96:25:@58562.4]
  assign _T_13820 = _T_13752 ? Mem1D_5_io_output : _T_13819; // @[Mux.scala 31:69:@58715.4]
  assign _T_13749 = RetimeWrapper_541_io_out; // @[package.scala 96:25:@58553.4 package.scala 96:25:@58554.4]
  assign _T_13821 = _T_13749 ? Mem1D_3_io_output : _T_13820; // @[Mux.scala 31:69:@58716.4]
  assign _T_13746 = RetimeWrapper_540_io_out; // @[package.scala 96:25:@58545.4 package.scala 96:25:@58546.4]
  assign _T_13979 = RetimeWrapper_578_io_out; // @[package.scala 96:25:@58929.4 package.scala 96:25:@58930.4]
  assign _T_13983 = _T_13979 ? Mem1D_37_io_output : Mem1D_39_io_output; // @[Mux.scala 31:69:@58939.4]
  assign _T_13976 = RetimeWrapper_577_io_out; // @[package.scala 96:25:@58921.4 package.scala 96:25:@58922.4]
  assign _T_13984 = _T_13976 ? Mem1D_35_io_output : _T_13983; // @[Mux.scala 31:69:@58940.4]
  assign _T_13973 = RetimeWrapper_576_io_out; // @[package.scala 96:25:@58913.4 package.scala 96:25:@58914.4]
  assign _T_13985 = _T_13973 ? Mem1D_33_io_output : _T_13984; // @[Mux.scala 31:69:@58941.4]
  assign _T_13970 = RetimeWrapper_575_io_out; // @[package.scala 96:25:@58905.4 package.scala 96:25:@58906.4]
  assign _T_13986 = _T_13970 ? Mem1D_31_io_output : _T_13985; // @[Mux.scala 31:69:@58942.4]
  assign _T_13967 = RetimeWrapper_574_io_out; // @[package.scala 96:25:@58897.4 package.scala 96:25:@58898.4]
  assign _T_13987 = _T_13967 ? Mem1D_29_io_output : _T_13986; // @[Mux.scala 31:69:@58943.4]
  assign _T_13964 = RetimeWrapper_573_io_out; // @[package.scala 96:25:@58889.4 package.scala 96:25:@58890.4]
  assign _T_13988 = _T_13964 ? Mem1D_27_io_output : _T_13987; // @[Mux.scala 31:69:@58944.4]
  assign _T_13961 = RetimeWrapper_572_io_out; // @[package.scala 96:25:@58881.4 package.scala 96:25:@58882.4]
  assign _T_13989 = _T_13961 ? Mem1D_25_io_output : _T_13988; // @[Mux.scala 31:69:@58945.4]
  assign _T_13958 = RetimeWrapper_571_io_out; // @[package.scala 96:25:@58873.4 package.scala 96:25:@58874.4]
  assign _T_13990 = _T_13958 ? Mem1D_23_io_output : _T_13989; // @[Mux.scala 31:69:@58946.4]
  assign _T_13955 = RetimeWrapper_570_io_out; // @[package.scala 96:25:@58865.4 package.scala 96:25:@58866.4]
  assign _T_13991 = _T_13955 ? Mem1D_21_io_output : _T_13990; // @[Mux.scala 31:69:@58947.4]
  assign _T_13952 = RetimeWrapper_569_io_out; // @[package.scala 96:25:@58857.4 package.scala 96:25:@58858.4]
  assign _T_13992 = _T_13952 ? Mem1D_19_io_output : _T_13991; // @[Mux.scala 31:69:@58948.4]
  assign _T_13949 = RetimeWrapper_568_io_out; // @[package.scala 96:25:@58849.4 package.scala 96:25:@58850.4]
  assign _T_13993 = _T_13949 ? Mem1D_17_io_output : _T_13992; // @[Mux.scala 31:69:@58949.4]
  assign _T_13946 = RetimeWrapper_567_io_out; // @[package.scala 96:25:@58841.4 package.scala 96:25:@58842.4]
  assign _T_13994 = _T_13946 ? Mem1D_15_io_output : _T_13993; // @[Mux.scala 31:69:@58950.4]
  assign _T_13943 = RetimeWrapper_566_io_out; // @[package.scala 96:25:@58833.4 package.scala 96:25:@58834.4]
  assign _T_13995 = _T_13943 ? Mem1D_13_io_output : _T_13994; // @[Mux.scala 31:69:@58951.4]
  assign _T_13940 = RetimeWrapper_565_io_out; // @[package.scala 96:25:@58825.4 package.scala 96:25:@58826.4]
  assign _T_13996 = _T_13940 ? Mem1D_11_io_output : _T_13995; // @[Mux.scala 31:69:@58952.4]
  assign _T_13937 = RetimeWrapper_564_io_out; // @[package.scala 96:25:@58817.4 package.scala 96:25:@58818.4]
  assign _T_13997 = _T_13937 ? Mem1D_9_io_output : _T_13996; // @[Mux.scala 31:69:@58953.4]
  assign _T_13934 = RetimeWrapper_563_io_out; // @[package.scala 96:25:@58809.4 package.scala 96:25:@58810.4]
  assign _T_13998 = _T_13934 ? Mem1D_7_io_output : _T_13997; // @[Mux.scala 31:69:@58954.4]
  assign _T_13931 = RetimeWrapper_562_io_out; // @[package.scala 96:25:@58801.4 package.scala 96:25:@58802.4]
  assign _T_13999 = _T_13931 ? Mem1D_5_io_output : _T_13998; // @[Mux.scala 31:69:@58955.4]
  assign _T_13928 = RetimeWrapper_561_io_out; // @[package.scala 96:25:@58793.4 package.scala 96:25:@58794.4]
  assign _T_14000 = _T_13928 ? Mem1D_3_io_output : _T_13999; // @[Mux.scala 31:69:@58956.4]
  assign _T_13925 = RetimeWrapper_560_io_out; // @[package.scala 96:25:@58785.4 package.scala 96:25:@58786.4]
  assign _T_14158 = RetimeWrapper_598_io_out; // @[package.scala 96:25:@59169.4 package.scala 96:25:@59170.4]
  assign _T_14162 = _T_14158 ? Mem1D_36_io_output : Mem1D_38_io_output; // @[Mux.scala 31:69:@59179.4]
  assign _T_14155 = RetimeWrapper_597_io_out; // @[package.scala 96:25:@59161.4 package.scala 96:25:@59162.4]
  assign _T_14163 = _T_14155 ? Mem1D_34_io_output : _T_14162; // @[Mux.scala 31:69:@59180.4]
  assign _T_14152 = RetimeWrapper_596_io_out; // @[package.scala 96:25:@59153.4 package.scala 96:25:@59154.4]
  assign _T_14164 = _T_14152 ? Mem1D_32_io_output : _T_14163; // @[Mux.scala 31:69:@59181.4]
  assign _T_14149 = RetimeWrapper_595_io_out; // @[package.scala 96:25:@59145.4 package.scala 96:25:@59146.4]
  assign _T_14165 = _T_14149 ? Mem1D_30_io_output : _T_14164; // @[Mux.scala 31:69:@59182.4]
  assign _T_14146 = RetimeWrapper_594_io_out; // @[package.scala 96:25:@59137.4 package.scala 96:25:@59138.4]
  assign _T_14166 = _T_14146 ? Mem1D_28_io_output : _T_14165; // @[Mux.scala 31:69:@59183.4]
  assign _T_14143 = RetimeWrapper_593_io_out; // @[package.scala 96:25:@59129.4 package.scala 96:25:@59130.4]
  assign _T_14167 = _T_14143 ? Mem1D_26_io_output : _T_14166; // @[Mux.scala 31:69:@59184.4]
  assign _T_14140 = RetimeWrapper_592_io_out; // @[package.scala 96:25:@59121.4 package.scala 96:25:@59122.4]
  assign _T_14168 = _T_14140 ? Mem1D_24_io_output : _T_14167; // @[Mux.scala 31:69:@59185.4]
  assign _T_14137 = RetimeWrapper_591_io_out; // @[package.scala 96:25:@59113.4 package.scala 96:25:@59114.4]
  assign _T_14169 = _T_14137 ? Mem1D_22_io_output : _T_14168; // @[Mux.scala 31:69:@59186.4]
  assign _T_14134 = RetimeWrapper_590_io_out; // @[package.scala 96:25:@59105.4 package.scala 96:25:@59106.4]
  assign _T_14170 = _T_14134 ? Mem1D_20_io_output : _T_14169; // @[Mux.scala 31:69:@59187.4]
  assign _T_14131 = RetimeWrapper_589_io_out; // @[package.scala 96:25:@59097.4 package.scala 96:25:@59098.4]
  assign _T_14171 = _T_14131 ? Mem1D_18_io_output : _T_14170; // @[Mux.scala 31:69:@59188.4]
  assign _T_14128 = RetimeWrapper_588_io_out; // @[package.scala 96:25:@59089.4 package.scala 96:25:@59090.4]
  assign _T_14172 = _T_14128 ? Mem1D_16_io_output : _T_14171; // @[Mux.scala 31:69:@59189.4]
  assign _T_14125 = RetimeWrapper_587_io_out; // @[package.scala 96:25:@59081.4 package.scala 96:25:@59082.4]
  assign _T_14173 = _T_14125 ? Mem1D_14_io_output : _T_14172; // @[Mux.scala 31:69:@59190.4]
  assign _T_14122 = RetimeWrapper_586_io_out; // @[package.scala 96:25:@59073.4 package.scala 96:25:@59074.4]
  assign _T_14174 = _T_14122 ? Mem1D_12_io_output : _T_14173; // @[Mux.scala 31:69:@59191.4]
  assign _T_14119 = RetimeWrapper_585_io_out; // @[package.scala 96:25:@59065.4 package.scala 96:25:@59066.4]
  assign _T_14175 = _T_14119 ? Mem1D_10_io_output : _T_14174; // @[Mux.scala 31:69:@59192.4]
  assign _T_14116 = RetimeWrapper_584_io_out; // @[package.scala 96:25:@59057.4 package.scala 96:25:@59058.4]
  assign _T_14176 = _T_14116 ? Mem1D_8_io_output : _T_14175; // @[Mux.scala 31:69:@59193.4]
  assign _T_14113 = RetimeWrapper_583_io_out; // @[package.scala 96:25:@59049.4 package.scala 96:25:@59050.4]
  assign _T_14177 = _T_14113 ? Mem1D_6_io_output : _T_14176; // @[Mux.scala 31:69:@59194.4]
  assign _T_14110 = RetimeWrapper_582_io_out; // @[package.scala 96:25:@59041.4 package.scala 96:25:@59042.4]
  assign _T_14178 = _T_14110 ? Mem1D_4_io_output : _T_14177; // @[Mux.scala 31:69:@59195.4]
  assign _T_14107 = RetimeWrapper_581_io_out; // @[package.scala 96:25:@59033.4 package.scala 96:25:@59034.4]
  assign _T_14179 = _T_14107 ? Mem1D_2_io_output : _T_14178; // @[Mux.scala 31:69:@59196.4]
  assign _T_14104 = RetimeWrapper_580_io_out; // @[package.scala 96:25:@59025.4 package.scala 96:25:@59026.4]
  assign io_rPort_29_output_0 = _T_14104 ? Mem1D_io_output : _T_14179; // @[MemPrimitives.scala 148:13:@59198.4]
  assign io_rPort_28_output_0 = _T_13925 ? Mem1D_1_io_output : _T_14000; // @[MemPrimitives.scala 148:13:@58958.4]
  assign io_rPort_27_output_0 = _T_13746 ? Mem1D_1_io_output : _T_13821; // @[MemPrimitives.scala 148:13:@58718.4]
  assign io_rPort_26_output_0 = _T_13567 ? Mem1D_io_output : _T_13642; // @[MemPrimitives.scala 148:13:@58478.4]
  assign io_rPort_25_output_0 = _T_13388 ? Mem1D_1_io_output : _T_13463; // @[MemPrimitives.scala 148:13:@58238.4]
  assign io_rPort_24_output_0 = _T_13209 ? Mem1D_1_io_output : _T_13284; // @[MemPrimitives.scala 148:13:@57998.4]
  assign io_rPort_23_output_0 = _T_13030 ? Mem1D_1_io_output : _T_13105; // @[MemPrimitives.scala 148:13:@57758.4]
  assign io_rPort_22_output_0 = _T_12851 ? Mem1D_io_output : _T_12926; // @[MemPrimitives.scala 148:13:@57518.4]
  assign io_rPort_21_output_0 = _T_12672 ? Mem1D_1_io_output : _T_12747; // @[MemPrimitives.scala 148:13:@57278.4]
  assign io_rPort_20_output_0 = _T_12493 ? Mem1D_1_io_output : _T_12568; // @[MemPrimitives.scala 148:13:@57038.4]
  assign io_rPort_19_output_0 = _T_12314 ? Mem1D_io_output : _T_12389; // @[MemPrimitives.scala 148:13:@56798.4]
  assign io_rPort_18_output_0 = _T_12135 ? Mem1D_1_io_output : _T_12210; // @[MemPrimitives.scala 148:13:@56558.4]
  assign io_rPort_17_output_0 = _T_11956 ? Mem1D_io_output : _T_12031; // @[MemPrimitives.scala 148:13:@56318.4]
  assign io_rPort_16_output_0 = _T_11777 ? Mem1D_io_output : _T_11852; // @[MemPrimitives.scala 148:13:@56078.4]
  assign io_rPort_15_output_0 = _T_11598 ? Mem1D_io_output : _T_11673; // @[MemPrimitives.scala 148:13:@55838.4]
  assign io_rPort_14_output_0 = _T_11419 ? Mem1D_1_io_output : _T_11494; // @[MemPrimitives.scala 148:13:@55598.4]
  assign io_rPort_13_output_0 = _T_11240 ? Mem1D_io_output : _T_11315; // @[MemPrimitives.scala 148:13:@55358.4]
  assign io_rPort_12_output_0 = _T_11061 ? Mem1D_1_io_output : _T_11136; // @[MemPrimitives.scala 148:13:@55118.4]
  assign io_rPort_11_output_0 = _T_10882 ? Mem1D_1_io_output : _T_10957; // @[MemPrimitives.scala 148:13:@54878.4]
  assign io_rPort_10_output_0 = _T_10703 ? Mem1D_io_output : _T_10778; // @[MemPrimitives.scala 148:13:@54638.4]
  assign io_rPort_9_output_0 = _T_10524 ? Mem1D_io_output : _T_10599; // @[MemPrimitives.scala 148:13:@54398.4]
  assign io_rPort_8_output_0 = _T_10345 ? Mem1D_1_io_output : _T_10420; // @[MemPrimitives.scala 148:13:@54158.4]
  assign io_rPort_7_output_0 = _T_10166 ? Mem1D_1_io_output : _T_10241; // @[MemPrimitives.scala 148:13:@53918.4]
  assign io_rPort_6_output_0 = _T_9987 ? Mem1D_1_io_output : _T_10062; // @[MemPrimitives.scala 148:13:@53678.4]
  assign io_rPort_5_output_0 = _T_9808 ? Mem1D_io_output : _T_9883; // @[MemPrimitives.scala 148:13:@53438.4]
  assign io_rPort_4_output_0 = _T_9629 ? Mem1D_io_output : _T_9704; // @[MemPrimitives.scala 148:13:@53198.4]
  assign io_rPort_3_output_0 = _T_9450 ? Mem1D_io_output : _T_9525; // @[MemPrimitives.scala 148:13:@52958.4]
  assign io_rPort_2_output_0 = _T_9271 ? Mem1D_1_io_output : _T_9346; // @[MemPrimitives.scala 148:13:@52718.4]
  assign io_rPort_1_output_0 = _T_9092 ? Mem1D_io_output : _T_9167; // @[MemPrimitives.scala 148:13:@52478.4]
  assign io_rPort_0_output_0 = _T_8913 ? Mem1D_io_output : _T_8988; // @[MemPrimitives.scala 148:13:@52238.4]
  assign Mem1D_clock = clock; // @[:@44320.4]
  assign Mem1D_reset = reset; // @[:@44321.4]
  assign Mem1D_io_r_ofs_0 = _T_2879[7:0]; // @[MemPrimitives.scala 127:28:@46419.4]
  assign Mem1D_io_r_backpressure = _T_2879[8]; // @[MemPrimitives.scala 128:32:@46420.4]
  assign Mem1D_io_w_ofs_0 = _T_1245[7:0]; // @[MemPrimitives.scala 94:28:@44989.4]
  assign Mem1D_io_w_data_0 = _T_1245[15:8]; // @[MemPrimitives.scala 95:29:@44990.4]
  assign Mem1D_io_w_en_0 = _T_1245[16]; // @[MemPrimitives.scala 96:27:@44991.4]
  assign Mem1D_1_clock = clock; // @[:@44336.4]
  assign Mem1D_1_reset = reset; // @[:@44337.4]
  assign Mem1D_1_io_r_ofs_0 = _T_3031[7:0]; // @[MemPrimitives.scala 127:28:@46562.4]
  assign Mem1D_1_io_r_backpressure = _T_3031[8]; // @[MemPrimitives.scala 128:32:@46563.4]
  assign Mem1D_1_io_w_ofs_0 = _T_1283[7:0]; // @[MemPrimitives.scala 94:28:@45022.4]
  assign Mem1D_1_io_w_data_0 = _T_1283[15:8]; // @[MemPrimitives.scala 95:29:@45023.4]
  assign Mem1D_1_io_w_en_0 = _T_1283[16]; // @[MemPrimitives.scala 96:27:@45024.4]
  assign Mem1D_2_clock = clock; // @[:@44352.4]
  assign Mem1D_2_reset = reset; // @[:@44353.4]
  assign Mem1D_2_io_r_ofs_0 = _T_3183[7:0]; // @[MemPrimitives.scala 127:28:@46705.4]
  assign Mem1D_2_io_r_backpressure = _T_3183[8]; // @[MemPrimitives.scala 128:32:@46706.4]
  assign Mem1D_2_io_w_ofs_0 = _T_1321[7:0]; // @[MemPrimitives.scala 94:28:@45055.4]
  assign Mem1D_2_io_w_data_0 = _T_1321[15:8]; // @[MemPrimitives.scala 95:29:@45056.4]
  assign Mem1D_2_io_w_en_0 = _T_1321[16]; // @[MemPrimitives.scala 96:27:@45057.4]
  assign Mem1D_3_clock = clock; // @[:@44368.4]
  assign Mem1D_3_reset = reset; // @[:@44369.4]
  assign Mem1D_3_io_r_ofs_0 = _T_3335[7:0]; // @[MemPrimitives.scala 127:28:@46848.4]
  assign Mem1D_3_io_r_backpressure = _T_3335[8]; // @[MemPrimitives.scala 128:32:@46849.4]
  assign Mem1D_3_io_w_ofs_0 = _T_1359[7:0]; // @[MemPrimitives.scala 94:28:@45088.4]
  assign Mem1D_3_io_w_data_0 = _T_1359[15:8]; // @[MemPrimitives.scala 95:29:@45089.4]
  assign Mem1D_3_io_w_en_0 = _T_1359[16]; // @[MemPrimitives.scala 96:27:@45090.4]
  assign Mem1D_4_clock = clock; // @[:@44384.4]
  assign Mem1D_4_reset = reset; // @[:@44385.4]
  assign Mem1D_4_io_r_ofs_0 = _T_3487[7:0]; // @[MemPrimitives.scala 127:28:@46991.4]
  assign Mem1D_4_io_r_backpressure = _T_3487[8]; // @[MemPrimitives.scala 128:32:@46992.4]
  assign Mem1D_4_io_w_ofs_0 = _T_1397[7:0]; // @[MemPrimitives.scala 94:28:@45121.4]
  assign Mem1D_4_io_w_data_0 = _T_1397[15:8]; // @[MemPrimitives.scala 95:29:@45122.4]
  assign Mem1D_4_io_w_en_0 = _T_1397[16]; // @[MemPrimitives.scala 96:27:@45123.4]
  assign Mem1D_5_clock = clock; // @[:@44400.4]
  assign Mem1D_5_reset = reset; // @[:@44401.4]
  assign Mem1D_5_io_r_ofs_0 = _T_3639[7:0]; // @[MemPrimitives.scala 127:28:@47134.4]
  assign Mem1D_5_io_r_backpressure = _T_3639[8]; // @[MemPrimitives.scala 128:32:@47135.4]
  assign Mem1D_5_io_w_ofs_0 = _T_1435[7:0]; // @[MemPrimitives.scala 94:28:@45154.4]
  assign Mem1D_5_io_w_data_0 = _T_1435[15:8]; // @[MemPrimitives.scala 95:29:@45155.4]
  assign Mem1D_5_io_w_en_0 = _T_1435[16]; // @[MemPrimitives.scala 96:27:@45156.4]
  assign Mem1D_6_clock = clock; // @[:@44416.4]
  assign Mem1D_6_reset = reset; // @[:@44417.4]
  assign Mem1D_6_io_r_ofs_0 = _T_3791[7:0]; // @[MemPrimitives.scala 127:28:@47277.4]
  assign Mem1D_6_io_r_backpressure = _T_3791[8]; // @[MemPrimitives.scala 128:32:@47278.4]
  assign Mem1D_6_io_w_ofs_0 = _T_1473[7:0]; // @[MemPrimitives.scala 94:28:@45187.4]
  assign Mem1D_6_io_w_data_0 = _T_1473[15:8]; // @[MemPrimitives.scala 95:29:@45188.4]
  assign Mem1D_6_io_w_en_0 = _T_1473[16]; // @[MemPrimitives.scala 96:27:@45189.4]
  assign Mem1D_7_clock = clock; // @[:@44432.4]
  assign Mem1D_7_reset = reset; // @[:@44433.4]
  assign Mem1D_7_io_r_ofs_0 = _T_3943[7:0]; // @[MemPrimitives.scala 127:28:@47420.4]
  assign Mem1D_7_io_r_backpressure = _T_3943[8]; // @[MemPrimitives.scala 128:32:@47421.4]
  assign Mem1D_7_io_w_ofs_0 = _T_1511[7:0]; // @[MemPrimitives.scala 94:28:@45220.4]
  assign Mem1D_7_io_w_data_0 = _T_1511[15:8]; // @[MemPrimitives.scala 95:29:@45221.4]
  assign Mem1D_7_io_w_en_0 = _T_1511[16]; // @[MemPrimitives.scala 96:27:@45222.4]
  assign Mem1D_8_clock = clock; // @[:@44448.4]
  assign Mem1D_8_reset = reset; // @[:@44449.4]
  assign Mem1D_8_io_r_ofs_0 = _T_4095[7:0]; // @[MemPrimitives.scala 127:28:@47563.4]
  assign Mem1D_8_io_r_backpressure = _T_4095[8]; // @[MemPrimitives.scala 128:32:@47564.4]
  assign Mem1D_8_io_w_ofs_0 = _T_1549[7:0]; // @[MemPrimitives.scala 94:28:@45253.4]
  assign Mem1D_8_io_w_data_0 = _T_1549[15:8]; // @[MemPrimitives.scala 95:29:@45254.4]
  assign Mem1D_8_io_w_en_0 = _T_1549[16]; // @[MemPrimitives.scala 96:27:@45255.4]
  assign Mem1D_9_clock = clock; // @[:@44464.4]
  assign Mem1D_9_reset = reset; // @[:@44465.4]
  assign Mem1D_9_io_r_ofs_0 = _T_4247[7:0]; // @[MemPrimitives.scala 127:28:@47706.4]
  assign Mem1D_9_io_r_backpressure = _T_4247[8]; // @[MemPrimitives.scala 128:32:@47707.4]
  assign Mem1D_9_io_w_ofs_0 = _T_1587[7:0]; // @[MemPrimitives.scala 94:28:@45286.4]
  assign Mem1D_9_io_w_data_0 = _T_1587[15:8]; // @[MemPrimitives.scala 95:29:@45287.4]
  assign Mem1D_9_io_w_en_0 = _T_1587[16]; // @[MemPrimitives.scala 96:27:@45288.4]
  assign Mem1D_10_clock = clock; // @[:@44480.4]
  assign Mem1D_10_reset = reset; // @[:@44481.4]
  assign Mem1D_10_io_r_ofs_0 = _T_4399[7:0]; // @[MemPrimitives.scala 127:28:@47849.4]
  assign Mem1D_10_io_r_backpressure = _T_4399[8]; // @[MemPrimitives.scala 128:32:@47850.4]
  assign Mem1D_10_io_w_ofs_0 = _T_1625[7:0]; // @[MemPrimitives.scala 94:28:@45319.4]
  assign Mem1D_10_io_w_data_0 = _T_1625[15:8]; // @[MemPrimitives.scala 95:29:@45320.4]
  assign Mem1D_10_io_w_en_0 = _T_1625[16]; // @[MemPrimitives.scala 96:27:@45321.4]
  assign Mem1D_11_clock = clock; // @[:@44496.4]
  assign Mem1D_11_reset = reset; // @[:@44497.4]
  assign Mem1D_11_io_r_ofs_0 = _T_4551[7:0]; // @[MemPrimitives.scala 127:28:@47992.4]
  assign Mem1D_11_io_r_backpressure = _T_4551[8]; // @[MemPrimitives.scala 128:32:@47993.4]
  assign Mem1D_11_io_w_ofs_0 = _T_1663[7:0]; // @[MemPrimitives.scala 94:28:@45352.4]
  assign Mem1D_11_io_w_data_0 = _T_1663[15:8]; // @[MemPrimitives.scala 95:29:@45353.4]
  assign Mem1D_11_io_w_en_0 = _T_1663[16]; // @[MemPrimitives.scala 96:27:@45354.4]
  assign Mem1D_12_clock = clock; // @[:@44512.4]
  assign Mem1D_12_reset = reset; // @[:@44513.4]
  assign Mem1D_12_io_r_ofs_0 = _T_4703[7:0]; // @[MemPrimitives.scala 127:28:@48135.4]
  assign Mem1D_12_io_r_backpressure = _T_4703[8]; // @[MemPrimitives.scala 128:32:@48136.4]
  assign Mem1D_12_io_w_ofs_0 = _T_1701[7:0]; // @[MemPrimitives.scala 94:28:@45385.4]
  assign Mem1D_12_io_w_data_0 = _T_1701[15:8]; // @[MemPrimitives.scala 95:29:@45386.4]
  assign Mem1D_12_io_w_en_0 = _T_1701[16]; // @[MemPrimitives.scala 96:27:@45387.4]
  assign Mem1D_13_clock = clock; // @[:@44528.4]
  assign Mem1D_13_reset = reset; // @[:@44529.4]
  assign Mem1D_13_io_r_ofs_0 = _T_4855[7:0]; // @[MemPrimitives.scala 127:28:@48278.4]
  assign Mem1D_13_io_r_backpressure = _T_4855[8]; // @[MemPrimitives.scala 128:32:@48279.4]
  assign Mem1D_13_io_w_ofs_0 = _T_1739[7:0]; // @[MemPrimitives.scala 94:28:@45418.4]
  assign Mem1D_13_io_w_data_0 = _T_1739[15:8]; // @[MemPrimitives.scala 95:29:@45419.4]
  assign Mem1D_13_io_w_en_0 = _T_1739[16]; // @[MemPrimitives.scala 96:27:@45420.4]
  assign Mem1D_14_clock = clock; // @[:@44544.4]
  assign Mem1D_14_reset = reset; // @[:@44545.4]
  assign Mem1D_14_io_r_ofs_0 = _T_5007[7:0]; // @[MemPrimitives.scala 127:28:@48421.4]
  assign Mem1D_14_io_r_backpressure = _T_5007[8]; // @[MemPrimitives.scala 128:32:@48422.4]
  assign Mem1D_14_io_w_ofs_0 = _T_1777[7:0]; // @[MemPrimitives.scala 94:28:@45451.4]
  assign Mem1D_14_io_w_data_0 = _T_1777[15:8]; // @[MemPrimitives.scala 95:29:@45452.4]
  assign Mem1D_14_io_w_en_0 = _T_1777[16]; // @[MemPrimitives.scala 96:27:@45453.4]
  assign Mem1D_15_clock = clock; // @[:@44560.4]
  assign Mem1D_15_reset = reset; // @[:@44561.4]
  assign Mem1D_15_io_r_ofs_0 = _T_5159[7:0]; // @[MemPrimitives.scala 127:28:@48564.4]
  assign Mem1D_15_io_r_backpressure = _T_5159[8]; // @[MemPrimitives.scala 128:32:@48565.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1815[7:0]; // @[MemPrimitives.scala 94:28:@45484.4]
  assign Mem1D_15_io_w_data_0 = _T_1815[15:8]; // @[MemPrimitives.scala 95:29:@45485.4]
  assign Mem1D_15_io_w_en_0 = _T_1815[16]; // @[MemPrimitives.scala 96:27:@45486.4]
  assign Mem1D_16_clock = clock; // @[:@44576.4]
  assign Mem1D_16_reset = reset; // @[:@44577.4]
  assign Mem1D_16_io_r_ofs_0 = _T_5311[7:0]; // @[MemPrimitives.scala 127:28:@48707.4]
  assign Mem1D_16_io_r_backpressure = _T_5311[8]; // @[MemPrimitives.scala 128:32:@48708.4]
  assign Mem1D_16_io_w_ofs_0 = _T_1853[7:0]; // @[MemPrimitives.scala 94:28:@45517.4]
  assign Mem1D_16_io_w_data_0 = _T_1853[15:8]; // @[MemPrimitives.scala 95:29:@45518.4]
  assign Mem1D_16_io_w_en_0 = _T_1853[16]; // @[MemPrimitives.scala 96:27:@45519.4]
  assign Mem1D_17_clock = clock; // @[:@44592.4]
  assign Mem1D_17_reset = reset; // @[:@44593.4]
  assign Mem1D_17_io_r_ofs_0 = _T_5463[7:0]; // @[MemPrimitives.scala 127:28:@48850.4]
  assign Mem1D_17_io_r_backpressure = _T_5463[8]; // @[MemPrimitives.scala 128:32:@48851.4]
  assign Mem1D_17_io_w_ofs_0 = _T_1891[7:0]; // @[MemPrimitives.scala 94:28:@45550.4]
  assign Mem1D_17_io_w_data_0 = _T_1891[15:8]; // @[MemPrimitives.scala 95:29:@45551.4]
  assign Mem1D_17_io_w_en_0 = _T_1891[16]; // @[MemPrimitives.scala 96:27:@45552.4]
  assign Mem1D_18_clock = clock; // @[:@44608.4]
  assign Mem1D_18_reset = reset; // @[:@44609.4]
  assign Mem1D_18_io_r_ofs_0 = _T_5615[7:0]; // @[MemPrimitives.scala 127:28:@48993.4]
  assign Mem1D_18_io_r_backpressure = _T_5615[8]; // @[MemPrimitives.scala 128:32:@48994.4]
  assign Mem1D_18_io_w_ofs_0 = _T_1929[7:0]; // @[MemPrimitives.scala 94:28:@45583.4]
  assign Mem1D_18_io_w_data_0 = _T_1929[15:8]; // @[MemPrimitives.scala 95:29:@45584.4]
  assign Mem1D_18_io_w_en_0 = _T_1929[16]; // @[MemPrimitives.scala 96:27:@45585.4]
  assign Mem1D_19_clock = clock; // @[:@44624.4]
  assign Mem1D_19_reset = reset; // @[:@44625.4]
  assign Mem1D_19_io_r_ofs_0 = _T_5767[7:0]; // @[MemPrimitives.scala 127:28:@49136.4]
  assign Mem1D_19_io_r_backpressure = _T_5767[8]; // @[MemPrimitives.scala 128:32:@49137.4]
  assign Mem1D_19_io_w_ofs_0 = _T_1967[7:0]; // @[MemPrimitives.scala 94:28:@45616.4]
  assign Mem1D_19_io_w_data_0 = _T_1967[15:8]; // @[MemPrimitives.scala 95:29:@45617.4]
  assign Mem1D_19_io_w_en_0 = _T_1967[16]; // @[MemPrimitives.scala 96:27:@45618.4]
  assign Mem1D_20_clock = clock; // @[:@44640.4]
  assign Mem1D_20_reset = reset; // @[:@44641.4]
  assign Mem1D_20_io_r_ofs_0 = _T_5919[7:0]; // @[MemPrimitives.scala 127:28:@49279.4]
  assign Mem1D_20_io_r_backpressure = _T_5919[8]; // @[MemPrimitives.scala 128:32:@49280.4]
  assign Mem1D_20_io_w_ofs_0 = _T_2005[7:0]; // @[MemPrimitives.scala 94:28:@45649.4]
  assign Mem1D_20_io_w_data_0 = _T_2005[15:8]; // @[MemPrimitives.scala 95:29:@45650.4]
  assign Mem1D_20_io_w_en_0 = _T_2005[16]; // @[MemPrimitives.scala 96:27:@45651.4]
  assign Mem1D_21_clock = clock; // @[:@44656.4]
  assign Mem1D_21_reset = reset; // @[:@44657.4]
  assign Mem1D_21_io_r_ofs_0 = _T_6071[7:0]; // @[MemPrimitives.scala 127:28:@49422.4]
  assign Mem1D_21_io_r_backpressure = _T_6071[8]; // @[MemPrimitives.scala 128:32:@49423.4]
  assign Mem1D_21_io_w_ofs_0 = _T_2043[7:0]; // @[MemPrimitives.scala 94:28:@45682.4]
  assign Mem1D_21_io_w_data_0 = _T_2043[15:8]; // @[MemPrimitives.scala 95:29:@45683.4]
  assign Mem1D_21_io_w_en_0 = _T_2043[16]; // @[MemPrimitives.scala 96:27:@45684.4]
  assign Mem1D_22_clock = clock; // @[:@44672.4]
  assign Mem1D_22_reset = reset; // @[:@44673.4]
  assign Mem1D_22_io_r_ofs_0 = _T_6223[7:0]; // @[MemPrimitives.scala 127:28:@49565.4]
  assign Mem1D_22_io_r_backpressure = _T_6223[8]; // @[MemPrimitives.scala 128:32:@49566.4]
  assign Mem1D_22_io_w_ofs_0 = _T_2081[7:0]; // @[MemPrimitives.scala 94:28:@45715.4]
  assign Mem1D_22_io_w_data_0 = _T_2081[15:8]; // @[MemPrimitives.scala 95:29:@45716.4]
  assign Mem1D_22_io_w_en_0 = _T_2081[16]; // @[MemPrimitives.scala 96:27:@45717.4]
  assign Mem1D_23_clock = clock; // @[:@44688.4]
  assign Mem1D_23_reset = reset; // @[:@44689.4]
  assign Mem1D_23_io_r_ofs_0 = _T_6375[7:0]; // @[MemPrimitives.scala 127:28:@49708.4]
  assign Mem1D_23_io_r_backpressure = _T_6375[8]; // @[MemPrimitives.scala 128:32:@49709.4]
  assign Mem1D_23_io_w_ofs_0 = _T_2119[7:0]; // @[MemPrimitives.scala 94:28:@45748.4]
  assign Mem1D_23_io_w_data_0 = _T_2119[15:8]; // @[MemPrimitives.scala 95:29:@45749.4]
  assign Mem1D_23_io_w_en_0 = _T_2119[16]; // @[MemPrimitives.scala 96:27:@45750.4]
  assign Mem1D_24_clock = clock; // @[:@44704.4]
  assign Mem1D_24_reset = reset; // @[:@44705.4]
  assign Mem1D_24_io_r_ofs_0 = _T_6527[7:0]; // @[MemPrimitives.scala 127:28:@49851.4]
  assign Mem1D_24_io_r_backpressure = _T_6527[8]; // @[MemPrimitives.scala 128:32:@49852.4]
  assign Mem1D_24_io_w_ofs_0 = _T_2157[7:0]; // @[MemPrimitives.scala 94:28:@45781.4]
  assign Mem1D_24_io_w_data_0 = _T_2157[15:8]; // @[MemPrimitives.scala 95:29:@45782.4]
  assign Mem1D_24_io_w_en_0 = _T_2157[16]; // @[MemPrimitives.scala 96:27:@45783.4]
  assign Mem1D_25_clock = clock; // @[:@44720.4]
  assign Mem1D_25_reset = reset; // @[:@44721.4]
  assign Mem1D_25_io_r_ofs_0 = _T_6679[7:0]; // @[MemPrimitives.scala 127:28:@49994.4]
  assign Mem1D_25_io_r_backpressure = _T_6679[8]; // @[MemPrimitives.scala 128:32:@49995.4]
  assign Mem1D_25_io_w_ofs_0 = _T_2195[7:0]; // @[MemPrimitives.scala 94:28:@45814.4]
  assign Mem1D_25_io_w_data_0 = _T_2195[15:8]; // @[MemPrimitives.scala 95:29:@45815.4]
  assign Mem1D_25_io_w_en_0 = _T_2195[16]; // @[MemPrimitives.scala 96:27:@45816.4]
  assign Mem1D_26_clock = clock; // @[:@44736.4]
  assign Mem1D_26_reset = reset; // @[:@44737.4]
  assign Mem1D_26_io_r_ofs_0 = _T_6831[7:0]; // @[MemPrimitives.scala 127:28:@50137.4]
  assign Mem1D_26_io_r_backpressure = _T_6831[8]; // @[MemPrimitives.scala 128:32:@50138.4]
  assign Mem1D_26_io_w_ofs_0 = _T_2233[7:0]; // @[MemPrimitives.scala 94:28:@45847.4]
  assign Mem1D_26_io_w_data_0 = _T_2233[15:8]; // @[MemPrimitives.scala 95:29:@45848.4]
  assign Mem1D_26_io_w_en_0 = _T_2233[16]; // @[MemPrimitives.scala 96:27:@45849.4]
  assign Mem1D_27_clock = clock; // @[:@44752.4]
  assign Mem1D_27_reset = reset; // @[:@44753.4]
  assign Mem1D_27_io_r_ofs_0 = _T_6983[7:0]; // @[MemPrimitives.scala 127:28:@50280.4]
  assign Mem1D_27_io_r_backpressure = _T_6983[8]; // @[MemPrimitives.scala 128:32:@50281.4]
  assign Mem1D_27_io_w_ofs_0 = _T_2271[7:0]; // @[MemPrimitives.scala 94:28:@45880.4]
  assign Mem1D_27_io_w_data_0 = _T_2271[15:8]; // @[MemPrimitives.scala 95:29:@45881.4]
  assign Mem1D_27_io_w_en_0 = _T_2271[16]; // @[MemPrimitives.scala 96:27:@45882.4]
  assign Mem1D_28_clock = clock; // @[:@44768.4]
  assign Mem1D_28_reset = reset; // @[:@44769.4]
  assign Mem1D_28_io_r_ofs_0 = _T_7135[7:0]; // @[MemPrimitives.scala 127:28:@50423.4]
  assign Mem1D_28_io_r_backpressure = _T_7135[8]; // @[MemPrimitives.scala 128:32:@50424.4]
  assign Mem1D_28_io_w_ofs_0 = _T_2309[7:0]; // @[MemPrimitives.scala 94:28:@45913.4]
  assign Mem1D_28_io_w_data_0 = _T_2309[15:8]; // @[MemPrimitives.scala 95:29:@45914.4]
  assign Mem1D_28_io_w_en_0 = _T_2309[16]; // @[MemPrimitives.scala 96:27:@45915.4]
  assign Mem1D_29_clock = clock; // @[:@44784.4]
  assign Mem1D_29_reset = reset; // @[:@44785.4]
  assign Mem1D_29_io_r_ofs_0 = _T_7287[7:0]; // @[MemPrimitives.scala 127:28:@50566.4]
  assign Mem1D_29_io_r_backpressure = _T_7287[8]; // @[MemPrimitives.scala 128:32:@50567.4]
  assign Mem1D_29_io_w_ofs_0 = _T_2347[7:0]; // @[MemPrimitives.scala 94:28:@45946.4]
  assign Mem1D_29_io_w_data_0 = _T_2347[15:8]; // @[MemPrimitives.scala 95:29:@45947.4]
  assign Mem1D_29_io_w_en_0 = _T_2347[16]; // @[MemPrimitives.scala 96:27:@45948.4]
  assign Mem1D_30_clock = clock; // @[:@44800.4]
  assign Mem1D_30_reset = reset; // @[:@44801.4]
  assign Mem1D_30_io_r_ofs_0 = _T_7439[7:0]; // @[MemPrimitives.scala 127:28:@50709.4]
  assign Mem1D_30_io_r_backpressure = _T_7439[8]; // @[MemPrimitives.scala 128:32:@50710.4]
  assign Mem1D_30_io_w_ofs_0 = _T_2385[7:0]; // @[MemPrimitives.scala 94:28:@45979.4]
  assign Mem1D_30_io_w_data_0 = _T_2385[15:8]; // @[MemPrimitives.scala 95:29:@45980.4]
  assign Mem1D_30_io_w_en_0 = _T_2385[16]; // @[MemPrimitives.scala 96:27:@45981.4]
  assign Mem1D_31_clock = clock; // @[:@44816.4]
  assign Mem1D_31_reset = reset; // @[:@44817.4]
  assign Mem1D_31_io_r_ofs_0 = _T_7591[7:0]; // @[MemPrimitives.scala 127:28:@50852.4]
  assign Mem1D_31_io_r_backpressure = _T_7591[8]; // @[MemPrimitives.scala 128:32:@50853.4]
  assign Mem1D_31_io_w_ofs_0 = _T_2423[7:0]; // @[MemPrimitives.scala 94:28:@46012.4]
  assign Mem1D_31_io_w_data_0 = _T_2423[15:8]; // @[MemPrimitives.scala 95:29:@46013.4]
  assign Mem1D_31_io_w_en_0 = _T_2423[16]; // @[MemPrimitives.scala 96:27:@46014.4]
  assign Mem1D_32_clock = clock; // @[:@44832.4]
  assign Mem1D_32_reset = reset; // @[:@44833.4]
  assign Mem1D_32_io_r_ofs_0 = _T_7743[7:0]; // @[MemPrimitives.scala 127:28:@50995.4]
  assign Mem1D_32_io_r_backpressure = _T_7743[8]; // @[MemPrimitives.scala 128:32:@50996.4]
  assign Mem1D_32_io_w_ofs_0 = _T_2461[7:0]; // @[MemPrimitives.scala 94:28:@46045.4]
  assign Mem1D_32_io_w_data_0 = _T_2461[15:8]; // @[MemPrimitives.scala 95:29:@46046.4]
  assign Mem1D_32_io_w_en_0 = _T_2461[16]; // @[MemPrimitives.scala 96:27:@46047.4]
  assign Mem1D_33_clock = clock; // @[:@44848.4]
  assign Mem1D_33_reset = reset; // @[:@44849.4]
  assign Mem1D_33_io_r_ofs_0 = _T_7895[7:0]; // @[MemPrimitives.scala 127:28:@51138.4]
  assign Mem1D_33_io_r_backpressure = _T_7895[8]; // @[MemPrimitives.scala 128:32:@51139.4]
  assign Mem1D_33_io_w_ofs_0 = _T_2499[7:0]; // @[MemPrimitives.scala 94:28:@46078.4]
  assign Mem1D_33_io_w_data_0 = _T_2499[15:8]; // @[MemPrimitives.scala 95:29:@46079.4]
  assign Mem1D_33_io_w_en_0 = _T_2499[16]; // @[MemPrimitives.scala 96:27:@46080.4]
  assign Mem1D_34_clock = clock; // @[:@44864.4]
  assign Mem1D_34_reset = reset; // @[:@44865.4]
  assign Mem1D_34_io_r_ofs_0 = _T_8047[7:0]; // @[MemPrimitives.scala 127:28:@51281.4]
  assign Mem1D_34_io_r_backpressure = _T_8047[8]; // @[MemPrimitives.scala 128:32:@51282.4]
  assign Mem1D_34_io_w_ofs_0 = _T_2537[7:0]; // @[MemPrimitives.scala 94:28:@46111.4]
  assign Mem1D_34_io_w_data_0 = _T_2537[15:8]; // @[MemPrimitives.scala 95:29:@46112.4]
  assign Mem1D_34_io_w_en_0 = _T_2537[16]; // @[MemPrimitives.scala 96:27:@46113.4]
  assign Mem1D_35_clock = clock; // @[:@44880.4]
  assign Mem1D_35_reset = reset; // @[:@44881.4]
  assign Mem1D_35_io_r_ofs_0 = _T_8199[7:0]; // @[MemPrimitives.scala 127:28:@51424.4]
  assign Mem1D_35_io_r_backpressure = _T_8199[8]; // @[MemPrimitives.scala 128:32:@51425.4]
  assign Mem1D_35_io_w_ofs_0 = _T_2575[7:0]; // @[MemPrimitives.scala 94:28:@46144.4]
  assign Mem1D_35_io_w_data_0 = _T_2575[15:8]; // @[MemPrimitives.scala 95:29:@46145.4]
  assign Mem1D_35_io_w_en_0 = _T_2575[16]; // @[MemPrimitives.scala 96:27:@46146.4]
  assign Mem1D_36_clock = clock; // @[:@44896.4]
  assign Mem1D_36_reset = reset; // @[:@44897.4]
  assign Mem1D_36_io_r_ofs_0 = _T_8351[7:0]; // @[MemPrimitives.scala 127:28:@51567.4]
  assign Mem1D_36_io_r_backpressure = _T_8351[8]; // @[MemPrimitives.scala 128:32:@51568.4]
  assign Mem1D_36_io_w_ofs_0 = _T_2613[7:0]; // @[MemPrimitives.scala 94:28:@46177.4]
  assign Mem1D_36_io_w_data_0 = _T_2613[15:8]; // @[MemPrimitives.scala 95:29:@46178.4]
  assign Mem1D_36_io_w_en_0 = _T_2613[16]; // @[MemPrimitives.scala 96:27:@46179.4]
  assign Mem1D_37_clock = clock; // @[:@44912.4]
  assign Mem1D_37_reset = reset; // @[:@44913.4]
  assign Mem1D_37_io_r_ofs_0 = _T_8503[7:0]; // @[MemPrimitives.scala 127:28:@51710.4]
  assign Mem1D_37_io_r_backpressure = _T_8503[8]; // @[MemPrimitives.scala 128:32:@51711.4]
  assign Mem1D_37_io_w_ofs_0 = _T_2651[7:0]; // @[MemPrimitives.scala 94:28:@46210.4]
  assign Mem1D_37_io_w_data_0 = _T_2651[15:8]; // @[MemPrimitives.scala 95:29:@46211.4]
  assign Mem1D_37_io_w_en_0 = _T_2651[16]; // @[MemPrimitives.scala 96:27:@46212.4]
  assign Mem1D_38_clock = clock; // @[:@44928.4]
  assign Mem1D_38_reset = reset; // @[:@44929.4]
  assign Mem1D_38_io_r_ofs_0 = _T_8655[7:0]; // @[MemPrimitives.scala 127:28:@51853.4]
  assign Mem1D_38_io_r_backpressure = _T_8655[8]; // @[MemPrimitives.scala 128:32:@51854.4]
  assign Mem1D_38_io_w_ofs_0 = _T_2689[7:0]; // @[MemPrimitives.scala 94:28:@46243.4]
  assign Mem1D_38_io_w_data_0 = _T_2689[15:8]; // @[MemPrimitives.scala 95:29:@46244.4]
  assign Mem1D_38_io_w_en_0 = _T_2689[16]; // @[MemPrimitives.scala 96:27:@46245.4]
  assign Mem1D_39_clock = clock; // @[:@44944.4]
  assign Mem1D_39_reset = reset; // @[:@44945.4]
  assign Mem1D_39_io_r_ofs_0 = _T_8807[7:0]; // @[MemPrimitives.scala 127:28:@51996.4]
  assign Mem1D_39_io_r_backpressure = _T_8807[8]; // @[MemPrimitives.scala 128:32:@51997.4]
  assign Mem1D_39_io_w_ofs_0 = _T_2727[7:0]; // @[MemPrimitives.scala 94:28:@46276.4]
  assign Mem1D_39_io_w_data_0 = _T_2727[15:8]; // @[MemPrimitives.scala 95:29:@46277.4]
  assign Mem1D_39_io_w_en_0 = _T_2727[16]; // @[MemPrimitives.scala 96:27:@46278.4]
  assign StickySelects_clock = clock; // @[:@46340.4]
  assign StickySelects_reset = reset; // @[:@46341.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_2735; // @[MemPrimitives.scala 122:60:@46342.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_2741; // @[MemPrimitives.scala 122:60:@46343.4]
  assign StickySelects_io_ins_2 = io_rPort_3_en_0 & _T_2747; // @[MemPrimitives.scala 122:60:@46344.4]
  assign StickySelects_io_ins_3 = io_rPort_4_en_0 & _T_2753; // @[MemPrimitives.scala 122:60:@46345.4]
  assign StickySelects_io_ins_4 = io_rPort_5_en_0 & _T_2759; // @[MemPrimitives.scala 122:60:@46346.4]
  assign StickySelects_io_ins_5 = io_rPort_9_en_0 & _T_2765; // @[MemPrimitives.scala 122:60:@46347.4]
  assign StickySelects_io_ins_6 = io_rPort_10_en_0 & _T_2771; // @[MemPrimitives.scala 122:60:@46348.4]
  assign StickySelects_io_ins_7 = io_rPort_13_en_0 & _T_2777; // @[MemPrimitives.scala 122:60:@46349.4]
  assign StickySelects_io_ins_8 = io_rPort_15_en_0 & _T_2783; // @[MemPrimitives.scala 122:60:@46350.4]
  assign StickySelects_io_ins_9 = io_rPort_16_en_0 & _T_2789; // @[MemPrimitives.scala 122:60:@46351.4]
  assign StickySelects_io_ins_10 = io_rPort_17_en_0 & _T_2795; // @[MemPrimitives.scala 122:60:@46352.4]
  assign StickySelects_io_ins_11 = io_rPort_19_en_0 & _T_2801; // @[MemPrimitives.scala 122:60:@46353.4]
  assign StickySelects_io_ins_12 = io_rPort_22_en_0 & _T_2807; // @[MemPrimitives.scala 122:60:@46354.4]
  assign StickySelects_io_ins_13 = io_rPort_26_en_0 & _T_2813; // @[MemPrimitives.scala 122:60:@46355.4]
  assign StickySelects_io_ins_14 = io_rPort_29_en_0 & _T_2819; // @[MemPrimitives.scala 122:60:@46356.4]
  assign StickySelects_1_clock = clock; // @[:@46483.4]
  assign StickySelects_1_reset = reset; // @[:@46484.4]
  assign StickySelects_1_io_ins_0 = io_rPort_2_en_0 & _T_2887; // @[MemPrimitives.scala 122:60:@46485.4]
  assign StickySelects_1_io_ins_1 = io_rPort_6_en_0 & _T_2893; // @[MemPrimitives.scala 122:60:@46486.4]
  assign StickySelects_1_io_ins_2 = io_rPort_7_en_0 & _T_2899; // @[MemPrimitives.scala 122:60:@46487.4]
  assign StickySelects_1_io_ins_3 = io_rPort_8_en_0 & _T_2905; // @[MemPrimitives.scala 122:60:@46488.4]
  assign StickySelects_1_io_ins_4 = io_rPort_11_en_0 & _T_2911; // @[MemPrimitives.scala 122:60:@46489.4]
  assign StickySelects_1_io_ins_5 = io_rPort_12_en_0 & _T_2917; // @[MemPrimitives.scala 122:60:@46490.4]
  assign StickySelects_1_io_ins_6 = io_rPort_14_en_0 & _T_2923; // @[MemPrimitives.scala 122:60:@46491.4]
  assign StickySelects_1_io_ins_7 = io_rPort_18_en_0 & _T_2929; // @[MemPrimitives.scala 122:60:@46492.4]
  assign StickySelects_1_io_ins_8 = io_rPort_20_en_0 & _T_2935; // @[MemPrimitives.scala 122:60:@46493.4]
  assign StickySelects_1_io_ins_9 = io_rPort_21_en_0 & _T_2941; // @[MemPrimitives.scala 122:60:@46494.4]
  assign StickySelects_1_io_ins_10 = io_rPort_23_en_0 & _T_2947; // @[MemPrimitives.scala 122:60:@46495.4]
  assign StickySelects_1_io_ins_11 = io_rPort_24_en_0 & _T_2953; // @[MemPrimitives.scala 122:60:@46496.4]
  assign StickySelects_1_io_ins_12 = io_rPort_25_en_0 & _T_2959; // @[MemPrimitives.scala 122:60:@46497.4]
  assign StickySelects_1_io_ins_13 = io_rPort_27_en_0 & _T_2965; // @[MemPrimitives.scala 122:60:@46498.4]
  assign StickySelects_1_io_ins_14 = io_rPort_28_en_0 & _T_2971; // @[MemPrimitives.scala 122:60:@46499.4]
  assign StickySelects_2_clock = clock; // @[:@46626.4]
  assign StickySelects_2_reset = reset; // @[:@46627.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_3039; // @[MemPrimitives.scala 122:60:@46628.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_3045; // @[MemPrimitives.scala 122:60:@46629.4]
  assign StickySelects_2_io_ins_2 = io_rPort_3_en_0 & _T_3051; // @[MemPrimitives.scala 122:60:@46630.4]
  assign StickySelects_2_io_ins_3 = io_rPort_4_en_0 & _T_3057; // @[MemPrimitives.scala 122:60:@46631.4]
  assign StickySelects_2_io_ins_4 = io_rPort_5_en_0 & _T_3063; // @[MemPrimitives.scala 122:60:@46632.4]
  assign StickySelects_2_io_ins_5 = io_rPort_9_en_0 & _T_3069; // @[MemPrimitives.scala 122:60:@46633.4]
  assign StickySelects_2_io_ins_6 = io_rPort_10_en_0 & _T_3075; // @[MemPrimitives.scala 122:60:@46634.4]
  assign StickySelects_2_io_ins_7 = io_rPort_13_en_0 & _T_3081; // @[MemPrimitives.scala 122:60:@46635.4]
  assign StickySelects_2_io_ins_8 = io_rPort_15_en_0 & _T_3087; // @[MemPrimitives.scala 122:60:@46636.4]
  assign StickySelects_2_io_ins_9 = io_rPort_16_en_0 & _T_3093; // @[MemPrimitives.scala 122:60:@46637.4]
  assign StickySelects_2_io_ins_10 = io_rPort_17_en_0 & _T_3099; // @[MemPrimitives.scala 122:60:@46638.4]
  assign StickySelects_2_io_ins_11 = io_rPort_19_en_0 & _T_3105; // @[MemPrimitives.scala 122:60:@46639.4]
  assign StickySelects_2_io_ins_12 = io_rPort_22_en_0 & _T_3111; // @[MemPrimitives.scala 122:60:@46640.4]
  assign StickySelects_2_io_ins_13 = io_rPort_26_en_0 & _T_3117; // @[MemPrimitives.scala 122:60:@46641.4]
  assign StickySelects_2_io_ins_14 = io_rPort_29_en_0 & _T_3123; // @[MemPrimitives.scala 122:60:@46642.4]
  assign StickySelects_3_clock = clock; // @[:@46769.4]
  assign StickySelects_3_reset = reset; // @[:@46770.4]
  assign StickySelects_3_io_ins_0 = io_rPort_2_en_0 & _T_3191; // @[MemPrimitives.scala 122:60:@46771.4]
  assign StickySelects_3_io_ins_1 = io_rPort_6_en_0 & _T_3197; // @[MemPrimitives.scala 122:60:@46772.4]
  assign StickySelects_3_io_ins_2 = io_rPort_7_en_0 & _T_3203; // @[MemPrimitives.scala 122:60:@46773.4]
  assign StickySelects_3_io_ins_3 = io_rPort_8_en_0 & _T_3209; // @[MemPrimitives.scala 122:60:@46774.4]
  assign StickySelects_3_io_ins_4 = io_rPort_11_en_0 & _T_3215; // @[MemPrimitives.scala 122:60:@46775.4]
  assign StickySelects_3_io_ins_5 = io_rPort_12_en_0 & _T_3221; // @[MemPrimitives.scala 122:60:@46776.4]
  assign StickySelects_3_io_ins_6 = io_rPort_14_en_0 & _T_3227; // @[MemPrimitives.scala 122:60:@46777.4]
  assign StickySelects_3_io_ins_7 = io_rPort_18_en_0 & _T_3233; // @[MemPrimitives.scala 122:60:@46778.4]
  assign StickySelects_3_io_ins_8 = io_rPort_20_en_0 & _T_3239; // @[MemPrimitives.scala 122:60:@46779.4]
  assign StickySelects_3_io_ins_9 = io_rPort_21_en_0 & _T_3245; // @[MemPrimitives.scala 122:60:@46780.4]
  assign StickySelects_3_io_ins_10 = io_rPort_23_en_0 & _T_3251; // @[MemPrimitives.scala 122:60:@46781.4]
  assign StickySelects_3_io_ins_11 = io_rPort_24_en_0 & _T_3257; // @[MemPrimitives.scala 122:60:@46782.4]
  assign StickySelects_3_io_ins_12 = io_rPort_25_en_0 & _T_3263; // @[MemPrimitives.scala 122:60:@46783.4]
  assign StickySelects_3_io_ins_13 = io_rPort_27_en_0 & _T_3269; // @[MemPrimitives.scala 122:60:@46784.4]
  assign StickySelects_3_io_ins_14 = io_rPort_28_en_0 & _T_3275; // @[MemPrimitives.scala 122:60:@46785.4]
  assign StickySelects_4_clock = clock; // @[:@46912.4]
  assign StickySelects_4_reset = reset; // @[:@46913.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_3343; // @[MemPrimitives.scala 122:60:@46914.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_3349; // @[MemPrimitives.scala 122:60:@46915.4]
  assign StickySelects_4_io_ins_2 = io_rPort_3_en_0 & _T_3355; // @[MemPrimitives.scala 122:60:@46916.4]
  assign StickySelects_4_io_ins_3 = io_rPort_4_en_0 & _T_3361; // @[MemPrimitives.scala 122:60:@46917.4]
  assign StickySelects_4_io_ins_4 = io_rPort_5_en_0 & _T_3367; // @[MemPrimitives.scala 122:60:@46918.4]
  assign StickySelects_4_io_ins_5 = io_rPort_9_en_0 & _T_3373; // @[MemPrimitives.scala 122:60:@46919.4]
  assign StickySelects_4_io_ins_6 = io_rPort_10_en_0 & _T_3379; // @[MemPrimitives.scala 122:60:@46920.4]
  assign StickySelects_4_io_ins_7 = io_rPort_13_en_0 & _T_3385; // @[MemPrimitives.scala 122:60:@46921.4]
  assign StickySelects_4_io_ins_8 = io_rPort_15_en_0 & _T_3391; // @[MemPrimitives.scala 122:60:@46922.4]
  assign StickySelects_4_io_ins_9 = io_rPort_16_en_0 & _T_3397; // @[MemPrimitives.scala 122:60:@46923.4]
  assign StickySelects_4_io_ins_10 = io_rPort_17_en_0 & _T_3403; // @[MemPrimitives.scala 122:60:@46924.4]
  assign StickySelects_4_io_ins_11 = io_rPort_19_en_0 & _T_3409; // @[MemPrimitives.scala 122:60:@46925.4]
  assign StickySelects_4_io_ins_12 = io_rPort_22_en_0 & _T_3415; // @[MemPrimitives.scala 122:60:@46926.4]
  assign StickySelects_4_io_ins_13 = io_rPort_26_en_0 & _T_3421; // @[MemPrimitives.scala 122:60:@46927.4]
  assign StickySelects_4_io_ins_14 = io_rPort_29_en_0 & _T_3427; // @[MemPrimitives.scala 122:60:@46928.4]
  assign StickySelects_5_clock = clock; // @[:@47055.4]
  assign StickySelects_5_reset = reset; // @[:@47056.4]
  assign StickySelects_5_io_ins_0 = io_rPort_2_en_0 & _T_3495; // @[MemPrimitives.scala 122:60:@47057.4]
  assign StickySelects_5_io_ins_1 = io_rPort_6_en_0 & _T_3501; // @[MemPrimitives.scala 122:60:@47058.4]
  assign StickySelects_5_io_ins_2 = io_rPort_7_en_0 & _T_3507; // @[MemPrimitives.scala 122:60:@47059.4]
  assign StickySelects_5_io_ins_3 = io_rPort_8_en_0 & _T_3513; // @[MemPrimitives.scala 122:60:@47060.4]
  assign StickySelects_5_io_ins_4 = io_rPort_11_en_0 & _T_3519; // @[MemPrimitives.scala 122:60:@47061.4]
  assign StickySelects_5_io_ins_5 = io_rPort_12_en_0 & _T_3525; // @[MemPrimitives.scala 122:60:@47062.4]
  assign StickySelects_5_io_ins_6 = io_rPort_14_en_0 & _T_3531; // @[MemPrimitives.scala 122:60:@47063.4]
  assign StickySelects_5_io_ins_7 = io_rPort_18_en_0 & _T_3537; // @[MemPrimitives.scala 122:60:@47064.4]
  assign StickySelects_5_io_ins_8 = io_rPort_20_en_0 & _T_3543; // @[MemPrimitives.scala 122:60:@47065.4]
  assign StickySelects_5_io_ins_9 = io_rPort_21_en_0 & _T_3549; // @[MemPrimitives.scala 122:60:@47066.4]
  assign StickySelects_5_io_ins_10 = io_rPort_23_en_0 & _T_3555; // @[MemPrimitives.scala 122:60:@47067.4]
  assign StickySelects_5_io_ins_11 = io_rPort_24_en_0 & _T_3561; // @[MemPrimitives.scala 122:60:@47068.4]
  assign StickySelects_5_io_ins_12 = io_rPort_25_en_0 & _T_3567; // @[MemPrimitives.scala 122:60:@47069.4]
  assign StickySelects_5_io_ins_13 = io_rPort_27_en_0 & _T_3573; // @[MemPrimitives.scala 122:60:@47070.4]
  assign StickySelects_5_io_ins_14 = io_rPort_28_en_0 & _T_3579; // @[MemPrimitives.scala 122:60:@47071.4]
  assign StickySelects_6_clock = clock; // @[:@47198.4]
  assign StickySelects_6_reset = reset; // @[:@47199.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_3647; // @[MemPrimitives.scala 122:60:@47200.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_3653; // @[MemPrimitives.scala 122:60:@47201.4]
  assign StickySelects_6_io_ins_2 = io_rPort_3_en_0 & _T_3659; // @[MemPrimitives.scala 122:60:@47202.4]
  assign StickySelects_6_io_ins_3 = io_rPort_4_en_0 & _T_3665; // @[MemPrimitives.scala 122:60:@47203.4]
  assign StickySelects_6_io_ins_4 = io_rPort_5_en_0 & _T_3671; // @[MemPrimitives.scala 122:60:@47204.4]
  assign StickySelects_6_io_ins_5 = io_rPort_9_en_0 & _T_3677; // @[MemPrimitives.scala 122:60:@47205.4]
  assign StickySelects_6_io_ins_6 = io_rPort_10_en_0 & _T_3683; // @[MemPrimitives.scala 122:60:@47206.4]
  assign StickySelects_6_io_ins_7 = io_rPort_13_en_0 & _T_3689; // @[MemPrimitives.scala 122:60:@47207.4]
  assign StickySelects_6_io_ins_8 = io_rPort_15_en_0 & _T_3695; // @[MemPrimitives.scala 122:60:@47208.4]
  assign StickySelects_6_io_ins_9 = io_rPort_16_en_0 & _T_3701; // @[MemPrimitives.scala 122:60:@47209.4]
  assign StickySelects_6_io_ins_10 = io_rPort_17_en_0 & _T_3707; // @[MemPrimitives.scala 122:60:@47210.4]
  assign StickySelects_6_io_ins_11 = io_rPort_19_en_0 & _T_3713; // @[MemPrimitives.scala 122:60:@47211.4]
  assign StickySelects_6_io_ins_12 = io_rPort_22_en_0 & _T_3719; // @[MemPrimitives.scala 122:60:@47212.4]
  assign StickySelects_6_io_ins_13 = io_rPort_26_en_0 & _T_3725; // @[MemPrimitives.scala 122:60:@47213.4]
  assign StickySelects_6_io_ins_14 = io_rPort_29_en_0 & _T_3731; // @[MemPrimitives.scala 122:60:@47214.4]
  assign StickySelects_7_clock = clock; // @[:@47341.4]
  assign StickySelects_7_reset = reset; // @[:@47342.4]
  assign StickySelects_7_io_ins_0 = io_rPort_2_en_0 & _T_3799; // @[MemPrimitives.scala 122:60:@47343.4]
  assign StickySelects_7_io_ins_1 = io_rPort_6_en_0 & _T_3805; // @[MemPrimitives.scala 122:60:@47344.4]
  assign StickySelects_7_io_ins_2 = io_rPort_7_en_0 & _T_3811; // @[MemPrimitives.scala 122:60:@47345.4]
  assign StickySelects_7_io_ins_3 = io_rPort_8_en_0 & _T_3817; // @[MemPrimitives.scala 122:60:@47346.4]
  assign StickySelects_7_io_ins_4 = io_rPort_11_en_0 & _T_3823; // @[MemPrimitives.scala 122:60:@47347.4]
  assign StickySelects_7_io_ins_5 = io_rPort_12_en_0 & _T_3829; // @[MemPrimitives.scala 122:60:@47348.4]
  assign StickySelects_7_io_ins_6 = io_rPort_14_en_0 & _T_3835; // @[MemPrimitives.scala 122:60:@47349.4]
  assign StickySelects_7_io_ins_7 = io_rPort_18_en_0 & _T_3841; // @[MemPrimitives.scala 122:60:@47350.4]
  assign StickySelects_7_io_ins_8 = io_rPort_20_en_0 & _T_3847; // @[MemPrimitives.scala 122:60:@47351.4]
  assign StickySelects_7_io_ins_9 = io_rPort_21_en_0 & _T_3853; // @[MemPrimitives.scala 122:60:@47352.4]
  assign StickySelects_7_io_ins_10 = io_rPort_23_en_0 & _T_3859; // @[MemPrimitives.scala 122:60:@47353.4]
  assign StickySelects_7_io_ins_11 = io_rPort_24_en_0 & _T_3865; // @[MemPrimitives.scala 122:60:@47354.4]
  assign StickySelects_7_io_ins_12 = io_rPort_25_en_0 & _T_3871; // @[MemPrimitives.scala 122:60:@47355.4]
  assign StickySelects_7_io_ins_13 = io_rPort_27_en_0 & _T_3877; // @[MemPrimitives.scala 122:60:@47356.4]
  assign StickySelects_7_io_ins_14 = io_rPort_28_en_0 & _T_3883; // @[MemPrimitives.scala 122:60:@47357.4]
  assign StickySelects_8_clock = clock; // @[:@47484.4]
  assign StickySelects_8_reset = reset; // @[:@47485.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_3951; // @[MemPrimitives.scala 122:60:@47486.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_3957; // @[MemPrimitives.scala 122:60:@47487.4]
  assign StickySelects_8_io_ins_2 = io_rPort_3_en_0 & _T_3963; // @[MemPrimitives.scala 122:60:@47488.4]
  assign StickySelects_8_io_ins_3 = io_rPort_4_en_0 & _T_3969; // @[MemPrimitives.scala 122:60:@47489.4]
  assign StickySelects_8_io_ins_4 = io_rPort_5_en_0 & _T_3975; // @[MemPrimitives.scala 122:60:@47490.4]
  assign StickySelects_8_io_ins_5 = io_rPort_9_en_0 & _T_3981; // @[MemPrimitives.scala 122:60:@47491.4]
  assign StickySelects_8_io_ins_6 = io_rPort_10_en_0 & _T_3987; // @[MemPrimitives.scala 122:60:@47492.4]
  assign StickySelects_8_io_ins_7 = io_rPort_13_en_0 & _T_3993; // @[MemPrimitives.scala 122:60:@47493.4]
  assign StickySelects_8_io_ins_8 = io_rPort_15_en_0 & _T_3999; // @[MemPrimitives.scala 122:60:@47494.4]
  assign StickySelects_8_io_ins_9 = io_rPort_16_en_0 & _T_4005; // @[MemPrimitives.scala 122:60:@47495.4]
  assign StickySelects_8_io_ins_10 = io_rPort_17_en_0 & _T_4011; // @[MemPrimitives.scala 122:60:@47496.4]
  assign StickySelects_8_io_ins_11 = io_rPort_19_en_0 & _T_4017; // @[MemPrimitives.scala 122:60:@47497.4]
  assign StickySelects_8_io_ins_12 = io_rPort_22_en_0 & _T_4023; // @[MemPrimitives.scala 122:60:@47498.4]
  assign StickySelects_8_io_ins_13 = io_rPort_26_en_0 & _T_4029; // @[MemPrimitives.scala 122:60:@47499.4]
  assign StickySelects_8_io_ins_14 = io_rPort_29_en_0 & _T_4035; // @[MemPrimitives.scala 122:60:@47500.4]
  assign StickySelects_9_clock = clock; // @[:@47627.4]
  assign StickySelects_9_reset = reset; // @[:@47628.4]
  assign StickySelects_9_io_ins_0 = io_rPort_2_en_0 & _T_4103; // @[MemPrimitives.scala 122:60:@47629.4]
  assign StickySelects_9_io_ins_1 = io_rPort_6_en_0 & _T_4109; // @[MemPrimitives.scala 122:60:@47630.4]
  assign StickySelects_9_io_ins_2 = io_rPort_7_en_0 & _T_4115; // @[MemPrimitives.scala 122:60:@47631.4]
  assign StickySelects_9_io_ins_3 = io_rPort_8_en_0 & _T_4121; // @[MemPrimitives.scala 122:60:@47632.4]
  assign StickySelects_9_io_ins_4 = io_rPort_11_en_0 & _T_4127; // @[MemPrimitives.scala 122:60:@47633.4]
  assign StickySelects_9_io_ins_5 = io_rPort_12_en_0 & _T_4133; // @[MemPrimitives.scala 122:60:@47634.4]
  assign StickySelects_9_io_ins_6 = io_rPort_14_en_0 & _T_4139; // @[MemPrimitives.scala 122:60:@47635.4]
  assign StickySelects_9_io_ins_7 = io_rPort_18_en_0 & _T_4145; // @[MemPrimitives.scala 122:60:@47636.4]
  assign StickySelects_9_io_ins_8 = io_rPort_20_en_0 & _T_4151; // @[MemPrimitives.scala 122:60:@47637.4]
  assign StickySelects_9_io_ins_9 = io_rPort_21_en_0 & _T_4157; // @[MemPrimitives.scala 122:60:@47638.4]
  assign StickySelects_9_io_ins_10 = io_rPort_23_en_0 & _T_4163; // @[MemPrimitives.scala 122:60:@47639.4]
  assign StickySelects_9_io_ins_11 = io_rPort_24_en_0 & _T_4169; // @[MemPrimitives.scala 122:60:@47640.4]
  assign StickySelects_9_io_ins_12 = io_rPort_25_en_0 & _T_4175; // @[MemPrimitives.scala 122:60:@47641.4]
  assign StickySelects_9_io_ins_13 = io_rPort_27_en_0 & _T_4181; // @[MemPrimitives.scala 122:60:@47642.4]
  assign StickySelects_9_io_ins_14 = io_rPort_28_en_0 & _T_4187; // @[MemPrimitives.scala 122:60:@47643.4]
  assign StickySelects_10_clock = clock; // @[:@47770.4]
  assign StickySelects_10_reset = reset; // @[:@47771.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_4255; // @[MemPrimitives.scala 122:60:@47772.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_4261; // @[MemPrimitives.scala 122:60:@47773.4]
  assign StickySelects_10_io_ins_2 = io_rPort_3_en_0 & _T_4267; // @[MemPrimitives.scala 122:60:@47774.4]
  assign StickySelects_10_io_ins_3 = io_rPort_4_en_0 & _T_4273; // @[MemPrimitives.scala 122:60:@47775.4]
  assign StickySelects_10_io_ins_4 = io_rPort_5_en_0 & _T_4279; // @[MemPrimitives.scala 122:60:@47776.4]
  assign StickySelects_10_io_ins_5 = io_rPort_9_en_0 & _T_4285; // @[MemPrimitives.scala 122:60:@47777.4]
  assign StickySelects_10_io_ins_6 = io_rPort_10_en_0 & _T_4291; // @[MemPrimitives.scala 122:60:@47778.4]
  assign StickySelects_10_io_ins_7 = io_rPort_13_en_0 & _T_4297; // @[MemPrimitives.scala 122:60:@47779.4]
  assign StickySelects_10_io_ins_8 = io_rPort_15_en_0 & _T_4303; // @[MemPrimitives.scala 122:60:@47780.4]
  assign StickySelects_10_io_ins_9 = io_rPort_16_en_0 & _T_4309; // @[MemPrimitives.scala 122:60:@47781.4]
  assign StickySelects_10_io_ins_10 = io_rPort_17_en_0 & _T_4315; // @[MemPrimitives.scala 122:60:@47782.4]
  assign StickySelects_10_io_ins_11 = io_rPort_19_en_0 & _T_4321; // @[MemPrimitives.scala 122:60:@47783.4]
  assign StickySelects_10_io_ins_12 = io_rPort_22_en_0 & _T_4327; // @[MemPrimitives.scala 122:60:@47784.4]
  assign StickySelects_10_io_ins_13 = io_rPort_26_en_0 & _T_4333; // @[MemPrimitives.scala 122:60:@47785.4]
  assign StickySelects_10_io_ins_14 = io_rPort_29_en_0 & _T_4339; // @[MemPrimitives.scala 122:60:@47786.4]
  assign StickySelects_11_clock = clock; // @[:@47913.4]
  assign StickySelects_11_reset = reset; // @[:@47914.4]
  assign StickySelects_11_io_ins_0 = io_rPort_2_en_0 & _T_4407; // @[MemPrimitives.scala 122:60:@47915.4]
  assign StickySelects_11_io_ins_1 = io_rPort_6_en_0 & _T_4413; // @[MemPrimitives.scala 122:60:@47916.4]
  assign StickySelects_11_io_ins_2 = io_rPort_7_en_0 & _T_4419; // @[MemPrimitives.scala 122:60:@47917.4]
  assign StickySelects_11_io_ins_3 = io_rPort_8_en_0 & _T_4425; // @[MemPrimitives.scala 122:60:@47918.4]
  assign StickySelects_11_io_ins_4 = io_rPort_11_en_0 & _T_4431; // @[MemPrimitives.scala 122:60:@47919.4]
  assign StickySelects_11_io_ins_5 = io_rPort_12_en_0 & _T_4437; // @[MemPrimitives.scala 122:60:@47920.4]
  assign StickySelects_11_io_ins_6 = io_rPort_14_en_0 & _T_4443; // @[MemPrimitives.scala 122:60:@47921.4]
  assign StickySelects_11_io_ins_7 = io_rPort_18_en_0 & _T_4449; // @[MemPrimitives.scala 122:60:@47922.4]
  assign StickySelects_11_io_ins_8 = io_rPort_20_en_0 & _T_4455; // @[MemPrimitives.scala 122:60:@47923.4]
  assign StickySelects_11_io_ins_9 = io_rPort_21_en_0 & _T_4461; // @[MemPrimitives.scala 122:60:@47924.4]
  assign StickySelects_11_io_ins_10 = io_rPort_23_en_0 & _T_4467; // @[MemPrimitives.scala 122:60:@47925.4]
  assign StickySelects_11_io_ins_11 = io_rPort_24_en_0 & _T_4473; // @[MemPrimitives.scala 122:60:@47926.4]
  assign StickySelects_11_io_ins_12 = io_rPort_25_en_0 & _T_4479; // @[MemPrimitives.scala 122:60:@47927.4]
  assign StickySelects_11_io_ins_13 = io_rPort_27_en_0 & _T_4485; // @[MemPrimitives.scala 122:60:@47928.4]
  assign StickySelects_11_io_ins_14 = io_rPort_28_en_0 & _T_4491; // @[MemPrimitives.scala 122:60:@47929.4]
  assign StickySelects_12_clock = clock; // @[:@48056.4]
  assign StickySelects_12_reset = reset; // @[:@48057.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_4559; // @[MemPrimitives.scala 122:60:@48058.4]
  assign StickySelects_12_io_ins_1 = io_rPort_1_en_0 & _T_4565; // @[MemPrimitives.scala 122:60:@48059.4]
  assign StickySelects_12_io_ins_2 = io_rPort_3_en_0 & _T_4571; // @[MemPrimitives.scala 122:60:@48060.4]
  assign StickySelects_12_io_ins_3 = io_rPort_4_en_0 & _T_4577; // @[MemPrimitives.scala 122:60:@48061.4]
  assign StickySelects_12_io_ins_4 = io_rPort_5_en_0 & _T_4583; // @[MemPrimitives.scala 122:60:@48062.4]
  assign StickySelects_12_io_ins_5 = io_rPort_9_en_0 & _T_4589; // @[MemPrimitives.scala 122:60:@48063.4]
  assign StickySelects_12_io_ins_6 = io_rPort_10_en_0 & _T_4595; // @[MemPrimitives.scala 122:60:@48064.4]
  assign StickySelects_12_io_ins_7 = io_rPort_13_en_0 & _T_4601; // @[MemPrimitives.scala 122:60:@48065.4]
  assign StickySelects_12_io_ins_8 = io_rPort_15_en_0 & _T_4607; // @[MemPrimitives.scala 122:60:@48066.4]
  assign StickySelects_12_io_ins_9 = io_rPort_16_en_0 & _T_4613; // @[MemPrimitives.scala 122:60:@48067.4]
  assign StickySelects_12_io_ins_10 = io_rPort_17_en_0 & _T_4619; // @[MemPrimitives.scala 122:60:@48068.4]
  assign StickySelects_12_io_ins_11 = io_rPort_19_en_0 & _T_4625; // @[MemPrimitives.scala 122:60:@48069.4]
  assign StickySelects_12_io_ins_12 = io_rPort_22_en_0 & _T_4631; // @[MemPrimitives.scala 122:60:@48070.4]
  assign StickySelects_12_io_ins_13 = io_rPort_26_en_0 & _T_4637; // @[MemPrimitives.scala 122:60:@48071.4]
  assign StickySelects_12_io_ins_14 = io_rPort_29_en_0 & _T_4643; // @[MemPrimitives.scala 122:60:@48072.4]
  assign StickySelects_13_clock = clock; // @[:@48199.4]
  assign StickySelects_13_reset = reset; // @[:@48200.4]
  assign StickySelects_13_io_ins_0 = io_rPort_2_en_0 & _T_4711; // @[MemPrimitives.scala 122:60:@48201.4]
  assign StickySelects_13_io_ins_1 = io_rPort_6_en_0 & _T_4717; // @[MemPrimitives.scala 122:60:@48202.4]
  assign StickySelects_13_io_ins_2 = io_rPort_7_en_0 & _T_4723; // @[MemPrimitives.scala 122:60:@48203.4]
  assign StickySelects_13_io_ins_3 = io_rPort_8_en_0 & _T_4729; // @[MemPrimitives.scala 122:60:@48204.4]
  assign StickySelects_13_io_ins_4 = io_rPort_11_en_0 & _T_4735; // @[MemPrimitives.scala 122:60:@48205.4]
  assign StickySelects_13_io_ins_5 = io_rPort_12_en_0 & _T_4741; // @[MemPrimitives.scala 122:60:@48206.4]
  assign StickySelects_13_io_ins_6 = io_rPort_14_en_0 & _T_4747; // @[MemPrimitives.scala 122:60:@48207.4]
  assign StickySelects_13_io_ins_7 = io_rPort_18_en_0 & _T_4753; // @[MemPrimitives.scala 122:60:@48208.4]
  assign StickySelects_13_io_ins_8 = io_rPort_20_en_0 & _T_4759; // @[MemPrimitives.scala 122:60:@48209.4]
  assign StickySelects_13_io_ins_9 = io_rPort_21_en_0 & _T_4765; // @[MemPrimitives.scala 122:60:@48210.4]
  assign StickySelects_13_io_ins_10 = io_rPort_23_en_0 & _T_4771; // @[MemPrimitives.scala 122:60:@48211.4]
  assign StickySelects_13_io_ins_11 = io_rPort_24_en_0 & _T_4777; // @[MemPrimitives.scala 122:60:@48212.4]
  assign StickySelects_13_io_ins_12 = io_rPort_25_en_0 & _T_4783; // @[MemPrimitives.scala 122:60:@48213.4]
  assign StickySelects_13_io_ins_13 = io_rPort_27_en_0 & _T_4789; // @[MemPrimitives.scala 122:60:@48214.4]
  assign StickySelects_13_io_ins_14 = io_rPort_28_en_0 & _T_4795; // @[MemPrimitives.scala 122:60:@48215.4]
  assign StickySelects_14_clock = clock; // @[:@48342.4]
  assign StickySelects_14_reset = reset; // @[:@48343.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_4863; // @[MemPrimitives.scala 122:60:@48344.4]
  assign StickySelects_14_io_ins_1 = io_rPort_1_en_0 & _T_4869; // @[MemPrimitives.scala 122:60:@48345.4]
  assign StickySelects_14_io_ins_2 = io_rPort_3_en_0 & _T_4875; // @[MemPrimitives.scala 122:60:@48346.4]
  assign StickySelects_14_io_ins_3 = io_rPort_4_en_0 & _T_4881; // @[MemPrimitives.scala 122:60:@48347.4]
  assign StickySelects_14_io_ins_4 = io_rPort_5_en_0 & _T_4887; // @[MemPrimitives.scala 122:60:@48348.4]
  assign StickySelects_14_io_ins_5 = io_rPort_9_en_0 & _T_4893; // @[MemPrimitives.scala 122:60:@48349.4]
  assign StickySelects_14_io_ins_6 = io_rPort_10_en_0 & _T_4899; // @[MemPrimitives.scala 122:60:@48350.4]
  assign StickySelects_14_io_ins_7 = io_rPort_13_en_0 & _T_4905; // @[MemPrimitives.scala 122:60:@48351.4]
  assign StickySelects_14_io_ins_8 = io_rPort_15_en_0 & _T_4911; // @[MemPrimitives.scala 122:60:@48352.4]
  assign StickySelects_14_io_ins_9 = io_rPort_16_en_0 & _T_4917; // @[MemPrimitives.scala 122:60:@48353.4]
  assign StickySelects_14_io_ins_10 = io_rPort_17_en_0 & _T_4923; // @[MemPrimitives.scala 122:60:@48354.4]
  assign StickySelects_14_io_ins_11 = io_rPort_19_en_0 & _T_4929; // @[MemPrimitives.scala 122:60:@48355.4]
  assign StickySelects_14_io_ins_12 = io_rPort_22_en_0 & _T_4935; // @[MemPrimitives.scala 122:60:@48356.4]
  assign StickySelects_14_io_ins_13 = io_rPort_26_en_0 & _T_4941; // @[MemPrimitives.scala 122:60:@48357.4]
  assign StickySelects_14_io_ins_14 = io_rPort_29_en_0 & _T_4947; // @[MemPrimitives.scala 122:60:@48358.4]
  assign StickySelects_15_clock = clock; // @[:@48485.4]
  assign StickySelects_15_reset = reset; // @[:@48486.4]
  assign StickySelects_15_io_ins_0 = io_rPort_2_en_0 & _T_5015; // @[MemPrimitives.scala 122:60:@48487.4]
  assign StickySelects_15_io_ins_1 = io_rPort_6_en_0 & _T_5021; // @[MemPrimitives.scala 122:60:@48488.4]
  assign StickySelects_15_io_ins_2 = io_rPort_7_en_0 & _T_5027; // @[MemPrimitives.scala 122:60:@48489.4]
  assign StickySelects_15_io_ins_3 = io_rPort_8_en_0 & _T_5033; // @[MemPrimitives.scala 122:60:@48490.4]
  assign StickySelects_15_io_ins_4 = io_rPort_11_en_0 & _T_5039; // @[MemPrimitives.scala 122:60:@48491.4]
  assign StickySelects_15_io_ins_5 = io_rPort_12_en_0 & _T_5045; // @[MemPrimitives.scala 122:60:@48492.4]
  assign StickySelects_15_io_ins_6 = io_rPort_14_en_0 & _T_5051; // @[MemPrimitives.scala 122:60:@48493.4]
  assign StickySelects_15_io_ins_7 = io_rPort_18_en_0 & _T_5057; // @[MemPrimitives.scala 122:60:@48494.4]
  assign StickySelects_15_io_ins_8 = io_rPort_20_en_0 & _T_5063; // @[MemPrimitives.scala 122:60:@48495.4]
  assign StickySelects_15_io_ins_9 = io_rPort_21_en_0 & _T_5069; // @[MemPrimitives.scala 122:60:@48496.4]
  assign StickySelects_15_io_ins_10 = io_rPort_23_en_0 & _T_5075; // @[MemPrimitives.scala 122:60:@48497.4]
  assign StickySelects_15_io_ins_11 = io_rPort_24_en_0 & _T_5081; // @[MemPrimitives.scala 122:60:@48498.4]
  assign StickySelects_15_io_ins_12 = io_rPort_25_en_0 & _T_5087; // @[MemPrimitives.scala 122:60:@48499.4]
  assign StickySelects_15_io_ins_13 = io_rPort_27_en_0 & _T_5093; // @[MemPrimitives.scala 122:60:@48500.4]
  assign StickySelects_15_io_ins_14 = io_rPort_28_en_0 & _T_5099; // @[MemPrimitives.scala 122:60:@48501.4]
  assign StickySelects_16_clock = clock; // @[:@48628.4]
  assign StickySelects_16_reset = reset; // @[:@48629.4]
  assign StickySelects_16_io_ins_0 = io_rPort_0_en_0 & _T_5167; // @[MemPrimitives.scala 122:60:@48630.4]
  assign StickySelects_16_io_ins_1 = io_rPort_1_en_0 & _T_5173; // @[MemPrimitives.scala 122:60:@48631.4]
  assign StickySelects_16_io_ins_2 = io_rPort_3_en_0 & _T_5179; // @[MemPrimitives.scala 122:60:@48632.4]
  assign StickySelects_16_io_ins_3 = io_rPort_4_en_0 & _T_5185; // @[MemPrimitives.scala 122:60:@48633.4]
  assign StickySelects_16_io_ins_4 = io_rPort_5_en_0 & _T_5191; // @[MemPrimitives.scala 122:60:@48634.4]
  assign StickySelects_16_io_ins_5 = io_rPort_9_en_0 & _T_5197; // @[MemPrimitives.scala 122:60:@48635.4]
  assign StickySelects_16_io_ins_6 = io_rPort_10_en_0 & _T_5203; // @[MemPrimitives.scala 122:60:@48636.4]
  assign StickySelects_16_io_ins_7 = io_rPort_13_en_0 & _T_5209; // @[MemPrimitives.scala 122:60:@48637.4]
  assign StickySelects_16_io_ins_8 = io_rPort_15_en_0 & _T_5215; // @[MemPrimitives.scala 122:60:@48638.4]
  assign StickySelects_16_io_ins_9 = io_rPort_16_en_0 & _T_5221; // @[MemPrimitives.scala 122:60:@48639.4]
  assign StickySelects_16_io_ins_10 = io_rPort_17_en_0 & _T_5227; // @[MemPrimitives.scala 122:60:@48640.4]
  assign StickySelects_16_io_ins_11 = io_rPort_19_en_0 & _T_5233; // @[MemPrimitives.scala 122:60:@48641.4]
  assign StickySelects_16_io_ins_12 = io_rPort_22_en_0 & _T_5239; // @[MemPrimitives.scala 122:60:@48642.4]
  assign StickySelects_16_io_ins_13 = io_rPort_26_en_0 & _T_5245; // @[MemPrimitives.scala 122:60:@48643.4]
  assign StickySelects_16_io_ins_14 = io_rPort_29_en_0 & _T_5251; // @[MemPrimitives.scala 122:60:@48644.4]
  assign StickySelects_17_clock = clock; // @[:@48771.4]
  assign StickySelects_17_reset = reset; // @[:@48772.4]
  assign StickySelects_17_io_ins_0 = io_rPort_2_en_0 & _T_5319; // @[MemPrimitives.scala 122:60:@48773.4]
  assign StickySelects_17_io_ins_1 = io_rPort_6_en_0 & _T_5325; // @[MemPrimitives.scala 122:60:@48774.4]
  assign StickySelects_17_io_ins_2 = io_rPort_7_en_0 & _T_5331; // @[MemPrimitives.scala 122:60:@48775.4]
  assign StickySelects_17_io_ins_3 = io_rPort_8_en_0 & _T_5337; // @[MemPrimitives.scala 122:60:@48776.4]
  assign StickySelects_17_io_ins_4 = io_rPort_11_en_0 & _T_5343; // @[MemPrimitives.scala 122:60:@48777.4]
  assign StickySelects_17_io_ins_5 = io_rPort_12_en_0 & _T_5349; // @[MemPrimitives.scala 122:60:@48778.4]
  assign StickySelects_17_io_ins_6 = io_rPort_14_en_0 & _T_5355; // @[MemPrimitives.scala 122:60:@48779.4]
  assign StickySelects_17_io_ins_7 = io_rPort_18_en_0 & _T_5361; // @[MemPrimitives.scala 122:60:@48780.4]
  assign StickySelects_17_io_ins_8 = io_rPort_20_en_0 & _T_5367; // @[MemPrimitives.scala 122:60:@48781.4]
  assign StickySelects_17_io_ins_9 = io_rPort_21_en_0 & _T_5373; // @[MemPrimitives.scala 122:60:@48782.4]
  assign StickySelects_17_io_ins_10 = io_rPort_23_en_0 & _T_5379; // @[MemPrimitives.scala 122:60:@48783.4]
  assign StickySelects_17_io_ins_11 = io_rPort_24_en_0 & _T_5385; // @[MemPrimitives.scala 122:60:@48784.4]
  assign StickySelects_17_io_ins_12 = io_rPort_25_en_0 & _T_5391; // @[MemPrimitives.scala 122:60:@48785.4]
  assign StickySelects_17_io_ins_13 = io_rPort_27_en_0 & _T_5397; // @[MemPrimitives.scala 122:60:@48786.4]
  assign StickySelects_17_io_ins_14 = io_rPort_28_en_0 & _T_5403; // @[MemPrimitives.scala 122:60:@48787.4]
  assign StickySelects_18_clock = clock; // @[:@48914.4]
  assign StickySelects_18_reset = reset; // @[:@48915.4]
  assign StickySelects_18_io_ins_0 = io_rPort_0_en_0 & _T_5471; // @[MemPrimitives.scala 122:60:@48916.4]
  assign StickySelects_18_io_ins_1 = io_rPort_1_en_0 & _T_5477; // @[MemPrimitives.scala 122:60:@48917.4]
  assign StickySelects_18_io_ins_2 = io_rPort_3_en_0 & _T_5483; // @[MemPrimitives.scala 122:60:@48918.4]
  assign StickySelects_18_io_ins_3 = io_rPort_4_en_0 & _T_5489; // @[MemPrimitives.scala 122:60:@48919.4]
  assign StickySelects_18_io_ins_4 = io_rPort_5_en_0 & _T_5495; // @[MemPrimitives.scala 122:60:@48920.4]
  assign StickySelects_18_io_ins_5 = io_rPort_9_en_0 & _T_5501; // @[MemPrimitives.scala 122:60:@48921.4]
  assign StickySelects_18_io_ins_6 = io_rPort_10_en_0 & _T_5507; // @[MemPrimitives.scala 122:60:@48922.4]
  assign StickySelects_18_io_ins_7 = io_rPort_13_en_0 & _T_5513; // @[MemPrimitives.scala 122:60:@48923.4]
  assign StickySelects_18_io_ins_8 = io_rPort_15_en_0 & _T_5519; // @[MemPrimitives.scala 122:60:@48924.4]
  assign StickySelects_18_io_ins_9 = io_rPort_16_en_0 & _T_5525; // @[MemPrimitives.scala 122:60:@48925.4]
  assign StickySelects_18_io_ins_10 = io_rPort_17_en_0 & _T_5531; // @[MemPrimitives.scala 122:60:@48926.4]
  assign StickySelects_18_io_ins_11 = io_rPort_19_en_0 & _T_5537; // @[MemPrimitives.scala 122:60:@48927.4]
  assign StickySelects_18_io_ins_12 = io_rPort_22_en_0 & _T_5543; // @[MemPrimitives.scala 122:60:@48928.4]
  assign StickySelects_18_io_ins_13 = io_rPort_26_en_0 & _T_5549; // @[MemPrimitives.scala 122:60:@48929.4]
  assign StickySelects_18_io_ins_14 = io_rPort_29_en_0 & _T_5555; // @[MemPrimitives.scala 122:60:@48930.4]
  assign StickySelects_19_clock = clock; // @[:@49057.4]
  assign StickySelects_19_reset = reset; // @[:@49058.4]
  assign StickySelects_19_io_ins_0 = io_rPort_2_en_0 & _T_5623; // @[MemPrimitives.scala 122:60:@49059.4]
  assign StickySelects_19_io_ins_1 = io_rPort_6_en_0 & _T_5629; // @[MemPrimitives.scala 122:60:@49060.4]
  assign StickySelects_19_io_ins_2 = io_rPort_7_en_0 & _T_5635; // @[MemPrimitives.scala 122:60:@49061.4]
  assign StickySelects_19_io_ins_3 = io_rPort_8_en_0 & _T_5641; // @[MemPrimitives.scala 122:60:@49062.4]
  assign StickySelects_19_io_ins_4 = io_rPort_11_en_0 & _T_5647; // @[MemPrimitives.scala 122:60:@49063.4]
  assign StickySelects_19_io_ins_5 = io_rPort_12_en_0 & _T_5653; // @[MemPrimitives.scala 122:60:@49064.4]
  assign StickySelects_19_io_ins_6 = io_rPort_14_en_0 & _T_5659; // @[MemPrimitives.scala 122:60:@49065.4]
  assign StickySelects_19_io_ins_7 = io_rPort_18_en_0 & _T_5665; // @[MemPrimitives.scala 122:60:@49066.4]
  assign StickySelects_19_io_ins_8 = io_rPort_20_en_0 & _T_5671; // @[MemPrimitives.scala 122:60:@49067.4]
  assign StickySelects_19_io_ins_9 = io_rPort_21_en_0 & _T_5677; // @[MemPrimitives.scala 122:60:@49068.4]
  assign StickySelects_19_io_ins_10 = io_rPort_23_en_0 & _T_5683; // @[MemPrimitives.scala 122:60:@49069.4]
  assign StickySelects_19_io_ins_11 = io_rPort_24_en_0 & _T_5689; // @[MemPrimitives.scala 122:60:@49070.4]
  assign StickySelects_19_io_ins_12 = io_rPort_25_en_0 & _T_5695; // @[MemPrimitives.scala 122:60:@49071.4]
  assign StickySelects_19_io_ins_13 = io_rPort_27_en_0 & _T_5701; // @[MemPrimitives.scala 122:60:@49072.4]
  assign StickySelects_19_io_ins_14 = io_rPort_28_en_0 & _T_5707; // @[MemPrimitives.scala 122:60:@49073.4]
  assign StickySelects_20_clock = clock; // @[:@49200.4]
  assign StickySelects_20_reset = reset; // @[:@49201.4]
  assign StickySelects_20_io_ins_0 = io_rPort_0_en_0 & _T_5775; // @[MemPrimitives.scala 122:60:@49202.4]
  assign StickySelects_20_io_ins_1 = io_rPort_1_en_0 & _T_5781; // @[MemPrimitives.scala 122:60:@49203.4]
  assign StickySelects_20_io_ins_2 = io_rPort_3_en_0 & _T_5787; // @[MemPrimitives.scala 122:60:@49204.4]
  assign StickySelects_20_io_ins_3 = io_rPort_4_en_0 & _T_5793; // @[MemPrimitives.scala 122:60:@49205.4]
  assign StickySelects_20_io_ins_4 = io_rPort_5_en_0 & _T_5799; // @[MemPrimitives.scala 122:60:@49206.4]
  assign StickySelects_20_io_ins_5 = io_rPort_9_en_0 & _T_5805; // @[MemPrimitives.scala 122:60:@49207.4]
  assign StickySelects_20_io_ins_6 = io_rPort_10_en_0 & _T_5811; // @[MemPrimitives.scala 122:60:@49208.4]
  assign StickySelects_20_io_ins_7 = io_rPort_13_en_0 & _T_5817; // @[MemPrimitives.scala 122:60:@49209.4]
  assign StickySelects_20_io_ins_8 = io_rPort_15_en_0 & _T_5823; // @[MemPrimitives.scala 122:60:@49210.4]
  assign StickySelects_20_io_ins_9 = io_rPort_16_en_0 & _T_5829; // @[MemPrimitives.scala 122:60:@49211.4]
  assign StickySelects_20_io_ins_10 = io_rPort_17_en_0 & _T_5835; // @[MemPrimitives.scala 122:60:@49212.4]
  assign StickySelects_20_io_ins_11 = io_rPort_19_en_0 & _T_5841; // @[MemPrimitives.scala 122:60:@49213.4]
  assign StickySelects_20_io_ins_12 = io_rPort_22_en_0 & _T_5847; // @[MemPrimitives.scala 122:60:@49214.4]
  assign StickySelects_20_io_ins_13 = io_rPort_26_en_0 & _T_5853; // @[MemPrimitives.scala 122:60:@49215.4]
  assign StickySelects_20_io_ins_14 = io_rPort_29_en_0 & _T_5859; // @[MemPrimitives.scala 122:60:@49216.4]
  assign StickySelects_21_clock = clock; // @[:@49343.4]
  assign StickySelects_21_reset = reset; // @[:@49344.4]
  assign StickySelects_21_io_ins_0 = io_rPort_2_en_0 & _T_5927; // @[MemPrimitives.scala 122:60:@49345.4]
  assign StickySelects_21_io_ins_1 = io_rPort_6_en_0 & _T_5933; // @[MemPrimitives.scala 122:60:@49346.4]
  assign StickySelects_21_io_ins_2 = io_rPort_7_en_0 & _T_5939; // @[MemPrimitives.scala 122:60:@49347.4]
  assign StickySelects_21_io_ins_3 = io_rPort_8_en_0 & _T_5945; // @[MemPrimitives.scala 122:60:@49348.4]
  assign StickySelects_21_io_ins_4 = io_rPort_11_en_0 & _T_5951; // @[MemPrimitives.scala 122:60:@49349.4]
  assign StickySelects_21_io_ins_5 = io_rPort_12_en_0 & _T_5957; // @[MemPrimitives.scala 122:60:@49350.4]
  assign StickySelects_21_io_ins_6 = io_rPort_14_en_0 & _T_5963; // @[MemPrimitives.scala 122:60:@49351.4]
  assign StickySelects_21_io_ins_7 = io_rPort_18_en_0 & _T_5969; // @[MemPrimitives.scala 122:60:@49352.4]
  assign StickySelects_21_io_ins_8 = io_rPort_20_en_0 & _T_5975; // @[MemPrimitives.scala 122:60:@49353.4]
  assign StickySelects_21_io_ins_9 = io_rPort_21_en_0 & _T_5981; // @[MemPrimitives.scala 122:60:@49354.4]
  assign StickySelects_21_io_ins_10 = io_rPort_23_en_0 & _T_5987; // @[MemPrimitives.scala 122:60:@49355.4]
  assign StickySelects_21_io_ins_11 = io_rPort_24_en_0 & _T_5993; // @[MemPrimitives.scala 122:60:@49356.4]
  assign StickySelects_21_io_ins_12 = io_rPort_25_en_0 & _T_5999; // @[MemPrimitives.scala 122:60:@49357.4]
  assign StickySelects_21_io_ins_13 = io_rPort_27_en_0 & _T_6005; // @[MemPrimitives.scala 122:60:@49358.4]
  assign StickySelects_21_io_ins_14 = io_rPort_28_en_0 & _T_6011; // @[MemPrimitives.scala 122:60:@49359.4]
  assign StickySelects_22_clock = clock; // @[:@49486.4]
  assign StickySelects_22_reset = reset; // @[:@49487.4]
  assign StickySelects_22_io_ins_0 = io_rPort_0_en_0 & _T_6079; // @[MemPrimitives.scala 122:60:@49488.4]
  assign StickySelects_22_io_ins_1 = io_rPort_1_en_0 & _T_6085; // @[MemPrimitives.scala 122:60:@49489.4]
  assign StickySelects_22_io_ins_2 = io_rPort_3_en_0 & _T_6091; // @[MemPrimitives.scala 122:60:@49490.4]
  assign StickySelects_22_io_ins_3 = io_rPort_4_en_0 & _T_6097; // @[MemPrimitives.scala 122:60:@49491.4]
  assign StickySelects_22_io_ins_4 = io_rPort_5_en_0 & _T_6103; // @[MemPrimitives.scala 122:60:@49492.4]
  assign StickySelects_22_io_ins_5 = io_rPort_9_en_0 & _T_6109; // @[MemPrimitives.scala 122:60:@49493.4]
  assign StickySelects_22_io_ins_6 = io_rPort_10_en_0 & _T_6115; // @[MemPrimitives.scala 122:60:@49494.4]
  assign StickySelects_22_io_ins_7 = io_rPort_13_en_0 & _T_6121; // @[MemPrimitives.scala 122:60:@49495.4]
  assign StickySelects_22_io_ins_8 = io_rPort_15_en_0 & _T_6127; // @[MemPrimitives.scala 122:60:@49496.4]
  assign StickySelects_22_io_ins_9 = io_rPort_16_en_0 & _T_6133; // @[MemPrimitives.scala 122:60:@49497.4]
  assign StickySelects_22_io_ins_10 = io_rPort_17_en_0 & _T_6139; // @[MemPrimitives.scala 122:60:@49498.4]
  assign StickySelects_22_io_ins_11 = io_rPort_19_en_0 & _T_6145; // @[MemPrimitives.scala 122:60:@49499.4]
  assign StickySelects_22_io_ins_12 = io_rPort_22_en_0 & _T_6151; // @[MemPrimitives.scala 122:60:@49500.4]
  assign StickySelects_22_io_ins_13 = io_rPort_26_en_0 & _T_6157; // @[MemPrimitives.scala 122:60:@49501.4]
  assign StickySelects_22_io_ins_14 = io_rPort_29_en_0 & _T_6163; // @[MemPrimitives.scala 122:60:@49502.4]
  assign StickySelects_23_clock = clock; // @[:@49629.4]
  assign StickySelects_23_reset = reset; // @[:@49630.4]
  assign StickySelects_23_io_ins_0 = io_rPort_2_en_0 & _T_6231; // @[MemPrimitives.scala 122:60:@49631.4]
  assign StickySelects_23_io_ins_1 = io_rPort_6_en_0 & _T_6237; // @[MemPrimitives.scala 122:60:@49632.4]
  assign StickySelects_23_io_ins_2 = io_rPort_7_en_0 & _T_6243; // @[MemPrimitives.scala 122:60:@49633.4]
  assign StickySelects_23_io_ins_3 = io_rPort_8_en_0 & _T_6249; // @[MemPrimitives.scala 122:60:@49634.4]
  assign StickySelects_23_io_ins_4 = io_rPort_11_en_0 & _T_6255; // @[MemPrimitives.scala 122:60:@49635.4]
  assign StickySelects_23_io_ins_5 = io_rPort_12_en_0 & _T_6261; // @[MemPrimitives.scala 122:60:@49636.4]
  assign StickySelects_23_io_ins_6 = io_rPort_14_en_0 & _T_6267; // @[MemPrimitives.scala 122:60:@49637.4]
  assign StickySelects_23_io_ins_7 = io_rPort_18_en_0 & _T_6273; // @[MemPrimitives.scala 122:60:@49638.4]
  assign StickySelects_23_io_ins_8 = io_rPort_20_en_0 & _T_6279; // @[MemPrimitives.scala 122:60:@49639.4]
  assign StickySelects_23_io_ins_9 = io_rPort_21_en_0 & _T_6285; // @[MemPrimitives.scala 122:60:@49640.4]
  assign StickySelects_23_io_ins_10 = io_rPort_23_en_0 & _T_6291; // @[MemPrimitives.scala 122:60:@49641.4]
  assign StickySelects_23_io_ins_11 = io_rPort_24_en_0 & _T_6297; // @[MemPrimitives.scala 122:60:@49642.4]
  assign StickySelects_23_io_ins_12 = io_rPort_25_en_0 & _T_6303; // @[MemPrimitives.scala 122:60:@49643.4]
  assign StickySelects_23_io_ins_13 = io_rPort_27_en_0 & _T_6309; // @[MemPrimitives.scala 122:60:@49644.4]
  assign StickySelects_23_io_ins_14 = io_rPort_28_en_0 & _T_6315; // @[MemPrimitives.scala 122:60:@49645.4]
  assign StickySelects_24_clock = clock; // @[:@49772.4]
  assign StickySelects_24_reset = reset; // @[:@49773.4]
  assign StickySelects_24_io_ins_0 = io_rPort_0_en_0 & _T_6383; // @[MemPrimitives.scala 122:60:@49774.4]
  assign StickySelects_24_io_ins_1 = io_rPort_1_en_0 & _T_6389; // @[MemPrimitives.scala 122:60:@49775.4]
  assign StickySelects_24_io_ins_2 = io_rPort_3_en_0 & _T_6395; // @[MemPrimitives.scala 122:60:@49776.4]
  assign StickySelects_24_io_ins_3 = io_rPort_4_en_0 & _T_6401; // @[MemPrimitives.scala 122:60:@49777.4]
  assign StickySelects_24_io_ins_4 = io_rPort_5_en_0 & _T_6407; // @[MemPrimitives.scala 122:60:@49778.4]
  assign StickySelects_24_io_ins_5 = io_rPort_9_en_0 & _T_6413; // @[MemPrimitives.scala 122:60:@49779.4]
  assign StickySelects_24_io_ins_6 = io_rPort_10_en_0 & _T_6419; // @[MemPrimitives.scala 122:60:@49780.4]
  assign StickySelects_24_io_ins_7 = io_rPort_13_en_0 & _T_6425; // @[MemPrimitives.scala 122:60:@49781.4]
  assign StickySelects_24_io_ins_8 = io_rPort_15_en_0 & _T_6431; // @[MemPrimitives.scala 122:60:@49782.4]
  assign StickySelects_24_io_ins_9 = io_rPort_16_en_0 & _T_6437; // @[MemPrimitives.scala 122:60:@49783.4]
  assign StickySelects_24_io_ins_10 = io_rPort_17_en_0 & _T_6443; // @[MemPrimitives.scala 122:60:@49784.4]
  assign StickySelects_24_io_ins_11 = io_rPort_19_en_0 & _T_6449; // @[MemPrimitives.scala 122:60:@49785.4]
  assign StickySelects_24_io_ins_12 = io_rPort_22_en_0 & _T_6455; // @[MemPrimitives.scala 122:60:@49786.4]
  assign StickySelects_24_io_ins_13 = io_rPort_26_en_0 & _T_6461; // @[MemPrimitives.scala 122:60:@49787.4]
  assign StickySelects_24_io_ins_14 = io_rPort_29_en_0 & _T_6467; // @[MemPrimitives.scala 122:60:@49788.4]
  assign StickySelects_25_clock = clock; // @[:@49915.4]
  assign StickySelects_25_reset = reset; // @[:@49916.4]
  assign StickySelects_25_io_ins_0 = io_rPort_2_en_0 & _T_6535; // @[MemPrimitives.scala 122:60:@49917.4]
  assign StickySelects_25_io_ins_1 = io_rPort_6_en_0 & _T_6541; // @[MemPrimitives.scala 122:60:@49918.4]
  assign StickySelects_25_io_ins_2 = io_rPort_7_en_0 & _T_6547; // @[MemPrimitives.scala 122:60:@49919.4]
  assign StickySelects_25_io_ins_3 = io_rPort_8_en_0 & _T_6553; // @[MemPrimitives.scala 122:60:@49920.4]
  assign StickySelects_25_io_ins_4 = io_rPort_11_en_0 & _T_6559; // @[MemPrimitives.scala 122:60:@49921.4]
  assign StickySelects_25_io_ins_5 = io_rPort_12_en_0 & _T_6565; // @[MemPrimitives.scala 122:60:@49922.4]
  assign StickySelects_25_io_ins_6 = io_rPort_14_en_0 & _T_6571; // @[MemPrimitives.scala 122:60:@49923.4]
  assign StickySelects_25_io_ins_7 = io_rPort_18_en_0 & _T_6577; // @[MemPrimitives.scala 122:60:@49924.4]
  assign StickySelects_25_io_ins_8 = io_rPort_20_en_0 & _T_6583; // @[MemPrimitives.scala 122:60:@49925.4]
  assign StickySelects_25_io_ins_9 = io_rPort_21_en_0 & _T_6589; // @[MemPrimitives.scala 122:60:@49926.4]
  assign StickySelects_25_io_ins_10 = io_rPort_23_en_0 & _T_6595; // @[MemPrimitives.scala 122:60:@49927.4]
  assign StickySelects_25_io_ins_11 = io_rPort_24_en_0 & _T_6601; // @[MemPrimitives.scala 122:60:@49928.4]
  assign StickySelects_25_io_ins_12 = io_rPort_25_en_0 & _T_6607; // @[MemPrimitives.scala 122:60:@49929.4]
  assign StickySelects_25_io_ins_13 = io_rPort_27_en_0 & _T_6613; // @[MemPrimitives.scala 122:60:@49930.4]
  assign StickySelects_25_io_ins_14 = io_rPort_28_en_0 & _T_6619; // @[MemPrimitives.scala 122:60:@49931.4]
  assign StickySelects_26_clock = clock; // @[:@50058.4]
  assign StickySelects_26_reset = reset; // @[:@50059.4]
  assign StickySelects_26_io_ins_0 = io_rPort_0_en_0 & _T_6687; // @[MemPrimitives.scala 122:60:@50060.4]
  assign StickySelects_26_io_ins_1 = io_rPort_1_en_0 & _T_6693; // @[MemPrimitives.scala 122:60:@50061.4]
  assign StickySelects_26_io_ins_2 = io_rPort_3_en_0 & _T_6699; // @[MemPrimitives.scala 122:60:@50062.4]
  assign StickySelects_26_io_ins_3 = io_rPort_4_en_0 & _T_6705; // @[MemPrimitives.scala 122:60:@50063.4]
  assign StickySelects_26_io_ins_4 = io_rPort_5_en_0 & _T_6711; // @[MemPrimitives.scala 122:60:@50064.4]
  assign StickySelects_26_io_ins_5 = io_rPort_9_en_0 & _T_6717; // @[MemPrimitives.scala 122:60:@50065.4]
  assign StickySelects_26_io_ins_6 = io_rPort_10_en_0 & _T_6723; // @[MemPrimitives.scala 122:60:@50066.4]
  assign StickySelects_26_io_ins_7 = io_rPort_13_en_0 & _T_6729; // @[MemPrimitives.scala 122:60:@50067.4]
  assign StickySelects_26_io_ins_8 = io_rPort_15_en_0 & _T_6735; // @[MemPrimitives.scala 122:60:@50068.4]
  assign StickySelects_26_io_ins_9 = io_rPort_16_en_0 & _T_6741; // @[MemPrimitives.scala 122:60:@50069.4]
  assign StickySelects_26_io_ins_10 = io_rPort_17_en_0 & _T_6747; // @[MemPrimitives.scala 122:60:@50070.4]
  assign StickySelects_26_io_ins_11 = io_rPort_19_en_0 & _T_6753; // @[MemPrimitives.scala 122:60:@50071.4]
  assign StickySelects_26_io_ins_12 = io_rPort_22_en_0 & _T_6759; // @[MemPrimitives.scala 122:60:@50072.4]
  assign StickySelects_26_io_ins_13 = io_rPort_26_en_0 & _T_6765; // @[MemPrimitives.scala 122:60:@50073.4]
  assign StickySelects_26_io_ins_14 = io_rPort_29_en_0 & _T_6771; // @[MemPrimitives.scala 122:60:@50074.4]
  assign StickySelects_27_clock = clock; // @[:@50201.4]
  assign StickySelects_27_reset = reset; // @[:@50202.4]
  assign StickySelects_27_io_ins_0 = io_rPort_2_en_0 & _T_6839; // @[MemPrimitives.scala 122:60:@50203.4]
  assign StickySelects_27_io_ins_1 = io_rPort_6_en_0 & _T_6845; // @[MemPrimitives.scala 122:60:@50204.4]
  assign StickySelects_27_io_ins_2 = io_rPort_7_en_0 & _T_6851; // @[MemPrimitives.scala 122:60:@50205.4]
  assign StickySelects_27_io_ins_3 = io_rPort_8_en_0 & _T_6857; // @[MemPrimitives.scala 122:60:@50206.4]
  assign StickySelects_27_io_ins_4 = io_rPort_11_en_0 & _T_6863; // @[MemPrimitives.scala 122:60:@50207.4]
  assign StickySelects_27_io_ins_5 = io_rPort_12_en_0 & _T_6869; // @[MemPrimitives.scala 122:60:@50208.4]
  assign StickySelects_27_io_ins_6 = io_rPort_14_en_0 & _T_6875; // @[MemPrimitives.scala 122:60:@50209.4]
  assign StickySelects_27_io_ins_7 = io_rPort_18_en_0 & _T_6881; // @[MemPrimitives.scala 122:60:@50210.4]
  assign StickySelects_27_io_ins_8 = io_rPort_20_en_0 & _T_6887; // @[MemPrimitives.scala 122:60:@50211.4]
  assign StickySelects_27_io_ins_9 = io_rPort_21_en_0 & _T_6893; // @[MemPrimitives.scala 122:60:@50212.4]
  assign StickySelects_27_io_ins_10 = io_rPort_23_en_0 & _T_6899; // @[MemPrimitives.scala 122:60:@50213.4]
  assign StickySelects_27_io_ins_11 = io_rPort_24_en_0 & _T_6905; // @[MemPrimitives.scala 122:60:@50214.4]
  assign StickySelects_27_io_ins_12 = io_rPort_25_en_0 & _T_6911; // @[MemPrimitives.scala 122:60:@50215.4]
  assign StickySelects_27_io_ins_13 = io_rPort_27_en_0 & _T_6917; // @[MemPrimitives.scala 122:60:@50216.4]
  assign StickySelects_27_io_ins_14 = io_rPort_28_en_0 & _T_6923; // @[MemPrimitives.scala 122:60:@50217.4]
  assign StickySelects_28_clock = clock; // @[:@50344.4]
  assign StickySelects_28_reset = reset; // @[:@50345.4]
  assign StickySelects_28_io_ins_0 = io_rPort_0_en_0 & _T_6991; // @[MemPrimitives.scala 122:60:@50346.4]
  assign StickySelects_28_io_ins_1 = io_rPort_1_en_0 & _T_6997; // @[MemPrimitives.scala 122:60:@50347.4]
  assign StickySelects_28_io_ins_2 = io_rPort_3_en_0 & _T_7003; // @[MemPrimitives.scala 122:60:@50348.4]
  assign StickySelects_28_io_ins_3 = io_rPort_4_en_0 & _T_7009; // @[MemPrimitives.scala 122:60:@50349.4]
  assign StickySelects_28_io_ins_4 = io_rPort_5_en_0 & _T_7015; // @[MemPrimitives.scala 122:60:@50350.4]
  assign StickySelects_28_io_ins_5 = io_rPort_9_en_0 & _T_7021; // @[MemPrimitives.scala 122:60:@50351.4]
  assign StickySelects_28_io_ins_6 = io_rPort_10_en_0 & _T_7027; // @[MemPrimitives.scala 122:60:@50352.4]
  assign StickySelects_28_io_ins_7 = io_rPort_13_en_0 & _T_7033; // @[MemPrimitives.scala 122:60:@50353.4]
  assign StickySelects_28_io_ins_8 = io_rPort_15_en_0 & _T_7039; // @[MemPrimitives.scala 122:60:@50354.4]
  assign StickySelects_28_io_ins_9 = io_rPort_16_en_0 & _T_7045; // @[MemPrimitives.scala 122:60:@50355.4]
  assign StickySelects_28_io_ins_10 = io_rPort_17_en_0 & _T_7051; // @[MemPrimitives.scala 122:60:@50356.4]
  assign StickySelects_28_io_ins_11 = io_rPort_19_en_0 & _T_7057; // @[MemPrimitives.scala 122:60:@50357.4]
  assign StickySelects_28_io_ins_12 = io_rPort_22_en_0 & _T_7063; // @[MemPrimitives.scala 122:60:@50358.4]
  assign StickySelects_28_io_ins_13 = io_rPort_26_en_0 & _T_7069; // @[MemPrimitives.scala 122:60:@50359.4]
  assign StickySelects_28_io_ins_14 = io_rPort_29_en_0 & _T_7075; // @[MemPrimitives.scala 122:60:@50360.4]
  assign StickySelects_29_clock = clock; // @[:@50487.4]
  assign StickySelects_29_reset = reset; // @[:@50488.4]
  assign StickySelects_29_io_ins_0 = io_rPort_2_en_0 & _T_7143; // @[MemPrimitives.scala 122:60:@50489.4]
  assign StickySelects_29_io_ins_1 = io_rPort_6_en_0 & _T_7149; // @[MemPrimitives.scala 122:60:@50490.4]
  assign StickySelects_29_io_ins_2 = io_rPort_7_en_0 & _T_7155; // @[MemPrimitives.scala 122:60:@50491.4]
  assign StickySelects_29_io_ins_3 = io_rPort_8_en_0 & _T_7161; // @[MemPrimitives.scala 122:60:@50492.4]
  assign StickySelects_29_io_ins_4 = io_rPort_11_en_0 & _T_7167; // @[MemPrimitives.scala 122:60:@50493.4]
  assign StickySelects_29_io_ins_5 = io_rPort_12_en_0 & _T_7173; // @[MemPrimitives.scala 122:60:@50494.4]
  assign StickySelects_29_io_ins_6 = io_rPort_14_en_0 & _T_7179; // @[MemPrimitives.scala 122:60:@50495.4]
  assign StickySelects_29_io_ins_7 = io_rPort_18_en_0 & _T_7185; // @[MemPrimitives.scala 122:60:@50496.4]
  assign StickySelects_29_io_ins_8 = io_rPort_20_en_0 & _T_7191; // @[MemPrimitives.scala 122:60:@50497.4]
  assign StickySelects_29_io_ins_9 = io_rPort_21_en_0 & _T_7197; // @[MemPrimitives.scala 122:60:@50498.4]
  assign StickySelects_29_io_ins_10 = io_rPort_23_en_0 & _T_7203; // @[MemPrimitives.scala 122:60:@50499.4]
  assign StickySelects_29_io_ins_11 = io_rPort_24_en_0 & _T_7209; // @[MemPrimitives.scala 122:60:@50500.4]
  assign StickySelects_29_io_ins_12 = io_rPort_25_en_0 & _T_7215; // @[MemPrimitives.scala 122:60:@50501.4]
  assign StickySelects_29_io_ins_13 = io_rPort_27_en_0 & _T_7221; // @[MemPrimitives.scala 122:60:@50502.4]
  assign StickySelects_29_io_ins_14 = io_rPort_28_en_0 & _T_7227; // @[MemPrimitives.scala 122:60:@50503.4]
  assign StickySelects_30_clock = clock; // @[:@50630.4]
  assign StickySelects_30_reset = reset; // @[:@50631.4]
  assign StickySelects_30_io_ins_0 = io_rPort_0_en_0 & _T_7295; // @[MemPrimitives.scala 122:60:@50632.4]
  assign StickySelects_30_io_ins_1 = io_rPort_1_en_0 & _T_7301; // @[MemPrimitives.scala 122:60:@50633.4]
  assign StickySelects_30_io_ins_2 = io_rPort_3_en_0 & _T_7307; // @[MemPrimitives.scala 122:60:@50634.4]
  assign StickySelects_30_io_ins_3 = io_rPort_4_en_0 & _T_7313; // @[MemPrimitives.scala 122:60:@50635.4]
  assign StickySelects_30_io_ins_4 = io_rPort_5_en_0 & _T_7319; // @[MemPrimitives.scala 122:60:@50636.4]
  assign StickySelects_30_io_ins_5 = io_rPort_9_en_0 & _T_7325; // @[MemPrimitives.scala 122:60:@50637.4]
  assign StickySelects_30_io_ins_6 = io_rPort_10_en_0 & _T_7331; // @[MemPrimitives.scala 122:60:@50638.4]
  assign StickySelects_30_io_ins_7 = io_rPort_13_en_0 & _T_7337; // @[MemPrimitives.scala 122:60:@50639.4]
  assign StickySelects_30_io_ins_8 = io_rPort_15_en_0 & _T_7343; // @[MemPrimitives.scala 122:60:@50640.4]
  assign StickySelects_30_io_ins_9 = io_rPort_16_en_0 & _T_7349; // @[MemPrimitives.scala 122:60:@50641.4]
  assign StickySelects_30_io_ins_10 = io_rPort_17_en_0 & _T_7355; // @[MemPrimitives.scala 122:60:@50642.4]
  assign StickySelects_30_io_ins_11 = io_rPort_19_en_0 & _T_7361; // @[MemPrimitives.scala 122:60:@50643.4]
  assign StickySelects_30_io_ins_12 = io_rPort_22_en_0 & _T_7367; // @[MemPrimitives.scala 122:60:@50644.4]
  assign StickySelects_30_io_ins_13 = io_rPort_26_en_0 & _T_7373; // @[MemPrimitives.scala 122:60:@50645.4]
  assign StickySelects_30_io_ins_14 = io_rPort_29_en_0 & _T_7379; // @[MemPrimitives.scala 122:60:@50646.4]
  assign StickySelects_31_clock = clock; // @[:@50773.4]
  assign StickySelects_31_reset = reset; // @[:@50774.4]
  assign StickySelects_31_io_ins_0 = io_rPort_2_en_0 & _T_7447; // @[MemPrimitives.scala 122:60:@50775.4]
  assign StickySelects_31_io_ins_1 = io_rPort_6_en_0 & _T_7453; // @[MemPrimitives.scala 122:60:@50776.4]
  assign StickySelects_31_io_ins_2 = io_rPort_7_en_0 & _T_7459; // @[MemPrimitives.scala 122:60:@50777.4]
  assign StickySelects_31_io_ins_3 = io_rPort_8_en_0 & _T_7465; // @[MemPrimitives.scala 122:60:@50778.4]
  assign StickySelects_31_io_ins_4 = io_rPort_11_en_0 & _T_7471; // @[MemPrimitives.scala 122:60:@50779.4]
  assign StickySelects_31_io_ins_5 = io_rPort_12_en_0 & _T_7477; // @[MemPrimitives.scala 122:60:@50780.4]
  assign StickySelects_31_io_ins_6 = io_rPort_14_en_0 & _T_7483; // @[MemPrimitives.scala 122:60:@50781.4]
  assign StickySelects_31_io_ins_7 = io_rPort_18_en_0 & _T_7489; // @[MemPrimitives.scala 122:60:@50782.4]
  assign StickySelects_31_io_ins_8 = io_rPort_20_en_0 & _T_7495; // @[MemPrimitives.scala 122:60:@50783.4]
  assign StickySelects_31_io_ins_9 = io_rPort_21_en_0 & _T_7501; // @[MemPrimitives.scala 122:60:@50784.4]
  assign StickySelects_31_io_ins_10 = io_rPort_23_en_0 & _T_7507; // @[MemPrimitives.scala 122:60:@50785.4]
  assign StickySelects_31_io_ins_11 = io_rPort_24_en_0 & _T_7513; // @[MemPrimitives.scala 122:60:@50786.4]
  assign StickySelects_31_io_ins_12 = io_rPort_25_en_0 & _T_7519; // @[MemPrimitives.scala 122:60:@50787.4]
  assign StickySelects_31_io_ins_13 = io_rPort_27_en_0 & _T_7525; // @[MemPrimitives.scala 122:60:@50788.4]
  assign StickySelects_31_io_ins_14 = io_rPort_28_en_0 & _T_7531; // @[MemPrimitives.scala 122:60:@50789.4]
  assign StickySelects_32_clock = clock; // @[:@50916.4]
  assign StickySelects_32_reset = reset; // @[:@50917.4]
  assign StickySelects_32_io_ins_0 = io_rPort_0_en_0 & _T_7599; // @[MemPrimitives.scala 122:60:@50918.4]
  assign StickySelects_32_io_ins_1 = io_rPort_1_en_0 & _T_7605; // @[MemPrimitives.scala 122:60:@50919.4]
  assign StickySelects_32_io_ins_2 = io_rPort_3_en_0 & _T_7611; // @[MemPrimitives.scala 122:60:@50920.4]
  assign StickySelects_32_io_ins_3 = io_rPort_4_en_0 & _T_7617; // @[MemPrimitives.scala 122:60:@50921.4]
  assign StickySelects_32_io_ins_4 = io_rPort_5_en_0 & _T_7623; // @[MemPrimitives.scala 122:60:@50922.4]
  assign StickySelects_32_io_ins_5 = io_rPort_9_en_0 & _T_7629; // @[MemPrimitives.scala 122:60:@50923.4]
  assign StickySelects_32_io_ins_6 = io_rPort_10_en_0 & _T_7635; // @[MemPrimitives.scala 122:60:@50924.4]
  assign StickySelects_32_io_ins_7 = io_rPort_13_en_0 & _T_7641; // @[MemPrimitives.scala 122:60:@50925.4]
  assign StickySelects_32_io_ins_8 = io_rPort_15_en_0 & _T_7647; // @[MemPrimitives.scala 122:60:@50926.4]
  assign StickySelects_32_io_ins_9 = io_rPort_16_en_0 & _T_7653; // @[MemPrimitives.scala 122:60:@50927.4]
  assign StickySelects_32_io_ins_10 = io_rPort_17_en_0 & _T_7659; // @[MemPrimitives.scala 122:60:@50928.4]
  assign StickySelects_32_io_ins_11 = io_rPort_19_en_0 & _T_7665; // @[MemPrimitives.scala 122:60:@50929.4]
  assign StickySelects_32_io_ins_12 = io_rPort_22_en_0 & _T_7671; // @[MemPrimitives.scala 122:60:@50930.4]
  assign StickySelects_32_io_ins_13 = io_rPort_26_en_0 & _T_7677; // @[MemPrimitives.scala 122:60:@50931.4]
  assign StickySelects_32_io_ins_14 = io_rPort_29_en_0 & _T_7683; // @[MemPrimitives.scala 122:60:@50932.4]
  assign StickySelects_33_clock = clock; // @[:@51059.4]
  assign StickySelects_33_reset = reset; // @[:@51060.4]
  assign StickySelects_33_io_ins_0 = io_rPort_2_en_0 & _T_7751; // @[MemPrimitives.scala 122:60:@51061.4]
  assign StickySelects_33_io_ins_1 = io_rPort_6_en_0 & _T_7757; // @[MemPrimitives.scala 122:60:@51062.4]
  assign StickySelects_33_io_ins_2 = io_rPort_7_en_0 & _T_7763; // @[MemPrimitives.scala 122:60:@51063.4]
  assign StickySelects_33_io_ins_3 = io_rPort_8_en_0 & _T_7769; // @[MemPrimitives.scala 122:60:@51064.4]
  assign StickySelects_33_io_ins_4 = io_rPort_11_en_0 & _T_7775; // @[MemPrimitives.scala 122:60:@51065.4]
  assign StickySelects_33_io_ins_5 = io_rPort_12_en_0 & _T_7781; // @[MemPrimitives.scala 122:60:@51066.4]
  assign StickySelects_33_io_ins_6 = io_rPort_14_en_0 & _T_7787; // @[MemPrimitives.scala 122:60:@51067.4]
  assign StickySelects_33_io_ins_7 = io_rPort_18_en_0 & _T_7793; // @[MemPrimitives.scala 122:60:@51068.4]
  assign StickySelects_33_io_ins_8 = io_rPort_20_en_0 & _T_7799; // @[MemPrimitives.scala 122:60:@51069.4]
  assign StickySelects_33_io_ins_9 = io_rPort_21_en_0 & _T_7805; // @[MemPrimitives.scala 122:60:@51070.4]
  assign StickySelects_33_io_ins_10 = io_rPort_23_en_0 & _T_7811; // @[MemPrimitives.scala 122:60:@51071.4]
  assign StickySelects_33_io_ins_11 = io_rPort_24_en_0 & _T_7817; // @[MemPrimitives.scala 122:60:@51072.4]
  assign StickySelects_33_io_ins_12 = io_rPort_25_en_0 & _T_7823; // @[MemPrimitives.scala 122:60:@51073.4]
  assign StickySelects_33_io_ins_13 = io_rPort_27_en_0 & _T_7829; // @[MemPrimitives.scala 122:60:@51074.4]
  assign StickySelects_33_io_ins_14 = io_rPort_28_en_0 & _T_7835; // @[MemPrimitives.scala 122:60:@51075.4]
  assign StickySelects_34_clock = clock; // @[:@51202.4]
  assign StickySelects_34_reset = reset; // @[:@51203.4]
  assign StickySelects_34_io_ins_0 = io_rPort_0_en_0 & _T_7903; // @[MemPrimitives.scala 122:60:@51204.4]
  assign StickySelects_34_io_ins_1 = io_rPort_1_en_0 & _T_7909; // @[MemPrimitives.scala 122:60:@51205.4]
  assign StickySelects_34_io_ins_2 = io_rPort_3_en_0 & _T_7915; // @[MemPrimitives.scala 122:60:@51206.4]
  assign StickySelects_34_io_ins_3 = io_rPort_4_en_0 & _T_7921; // @[MemPrimitives.scala 122:60:@51207.4]
  assign StickySelects_34_io_ins_4 = io_rPort_5_en_0 & _T_7927; // @[MemPrimitives.scala 122:60:@51208.4]
  assign StickySelects_34_io_ins_5 = io_rPort_9_en_0 & _T_7933; // @[MemPrimitives.scala 122:60:@51209.4]
  assign StickySelects_34_io_ins_6 = io_rPort_10_en_0 & _T_7939; // @[MemPrimitives.scala 122:60:@51210.4]
  assign StickySelects_34_io_ins_7 = io_rPort_13_en_0 & _T_7945; // @[MemPrimitives.scala 122:60:@51211.4]
  assign StickySelects_34_io_ins_8 = io_rPort_15_en_0 & _T_7951; // @[MemPrimitives.scala 122:60:@51212.4]
  assign StickySelects_34_io_ins_9 = io_rPort_16_en_0 & _T_7957; // @[MemPrimitives.scala 122:60:@51213.4]
  assign StickySelects_34_io_ins_10 = io_rPort_17_en_0 & _T_7963; // @[MemPrimitives.scala 122:60:@51214.4]
  assign StickySelects_34_io_ins_11 = io_rPort_19_en_0 & _T_7969; // @[MemPrimitives.scala 122:60:@51215.4]
  assign StickySelects_34_io_ins_12 = io_rPort_22_en_0 & _T_7975; // @[MemPrimitives.scala 122:60:@51216.4]
  assign StickySelects_34_io_ins_13 = io_rPort_26_en_0 & _T_7981; // @[MemPrimitives.scala 122:60:@51217.4]
  assign StickySelects_34_io_ins_14 = io_rPort_29_en_0 & _T_7987; // @[MemPrimitives.scala 122:60:@51218.4]
  assign StickySelects_35_clock = clock; // @[:@51345.4]
  assign StickySelects_35_reset = reset; // @[:@51346.4]
  assign StickySelects_35_io_ins_0 = io_rPort_2_en_0 & _T_8055; // @[MemPrimitives.scala 122:60:@51347.4]
  assign StickySelects_35_io_ins_1 = io_rPort_6_en_0 & _T_8061; // @[MemPrimitives.scala 122:60:@51348.4]
  assign StickySelects_35_io_ins_2 = io_rPort_7_en_0 & _T_8067; // @[MemPrimitives.scala 122:60:@51349.4]
  assign StickySelects_35_io_ins_3 = io_rPort_8_en_0 & _T_8073; // @[MemPrimitives.scala 122:60:@51350.4]
  assign StickySelects_35_io_ins_4 = io_rPort_11_en_0 & _T_8079; // @[MemPrimitives.scala 122:60:@51351.4]
  assign StickySelects_35_io_ins_5 = io_rPort_12_en_0 & _T_8085; // @[MemPrimitives.scala 122:60:@51352.4]
  assign StickySelects_35_io_ins_6 = io_rPort_14_en_0 & _T_8091; // @[MemPrimitives.scala 122:60:@51353.4]
  assign StickySelects_35_io_ins_7 = io_rPort_18_en_0 & _T_8097; // @[MemPrimitives.scala 122:60:@51354.4]
  assign StickySelects_35_io_ins_8 = io_rPort_20_en_0 & _T_8103; // @[MemPrimitives.scala 122:60:@51355.4]
  assign StickySelects_35_io_ins_9 = io_rPort_21_en_0 & _T_8109; // @[MemPrimitives.scala 122:60:@51356.4]
  assign StickySelects_35_io_ins_10 = io_rPort_23_en_0 & _T_8115; // @[MemPrimitives.scala 122:60:@51357.4]
  assign StickySelects_35_io_ins_11 = io_rPort_24_en_0 & _T_8121; // @[MemPrimitives.scala 122:60:@51358.4]
  assign StickySelects_35_io_ins_12 = io_rPort_25_en_0 & _T_8127; // @[MemPrimitives.scala 122:60:@51359.4]
  assign StickySelects_35_io_ins_13 = io_rPort_27_en_0 & _T_8133; // @[MemPrimitives.scala 122:60:@51360.4]
  assign StickySelects_35_io_ins_14 = io_rPort_28_en_0 & _T_8139; // @[MemPrimitives.scala 122:60:@51361.4]
  assign StickySelects_36_clock = clock; // @[:@51488.4]
  assign StickySelects_36_reset = reset; // @[:@51489.4]
  assign StickySelects_36_io_ins_0 = io_rPort_0_en_0 & _T_8207; // @[MemPrimitives.scala 122:60:@51490.4]
  assign StickySelects_36_io_ins_1 = io_rPort_1_en_0 & _T_8213; // @[MemPrimitives.scala 122:60:@51491.4]
  assign StickySelects_36_io_ins_2 = io_rPort_3_en_0 & _T_8219; // @[MemPrimitives.scala 122:60:@51492.4]
  assign StickySelects_36_io_ins_3 = io_rPort_4_en_0 & _T_8225; // @[MemPrimitives.scala 122:60:@51493.4]
  assign StickySelects_36_io_ins_4 = io_rPort_5_en_0 & _T_8231; // @[MemPrimitives.scala 122:60:@51494.4]
  assign StickySelects_36_io_ins_5 = io_rPort_9_en_0 & _T_8237; // @[MemPrimitives.scala 122:60:@51495.4]
  assign StickySelects_36_io_ins_6 = io_rPort_10_en_0 & _T_8243; // @[MemPrimitives.scala 122:60:@51496.4]
  assign StickySelects_36_io_ins_7 = io_rPort_13_en_0 & _T_8249; // @[MemPrimitives.scala 122:60:@51497.4]
  assign StickySelects_36_io_ins_8 = io_rPort_15_en_0 & _T_8255; // @[MemPrimitives.scala 122:60:@51498.4]
  assign StickySelects_36_io_ins_9 = io_rPort_16_en_0 & _T_8261; // @[MemPrimitives.scala 122:60:@51499.4]
  assign StickySelects_36_io_ins_10 = io_rPort_17_en_0 & _T_8267; // @[MemPrimitives.scala 122:60:@51500.4]
  assign StickySelects_36_io_ins_11 = io_rPort_19_en_0 & _T_8273; // @[MemPrimitives.scala 122:60:@51501.4]
  assign StickySelects_36_io_ins_12 = io_rPort_22_en_0 & _T_8279; // @[MemPrimitives.scala 122:60:@51502.4]
  assign StickySelects_36_io_ins_13 = io_rPort_26_en_0 & _T_8285; // @[MemPrimitives.scala 122:60:@51503.4]
  assign StickySelects_36_io_ins_14 = io_rPort_29_en_0 & _T_8291; // @[MemPrimitives.scala 122:60:@51504.4]
  assign StickySelects_37_clock = clock; // @[:@51631.4]
  assign StickySelects_37_reset = reset; // @[:@51632.4]
  assign StickySelects_37_io_ins_0 = io_rPort_2_en_0 & _T_8359; // @[MemPrimitives.scala 122:60:@51633.4]
  assign StickySelects_37_io_ins_1 = io_rPort_6_en_0 & _T_8365; // @[MemPrimitives.scala 122:60:@51634.4]
  assign StickySelects_37_io_ins_2 = io_rPort_7_en_0 & _T_8371; // @[MemPrimitives.scala 122:60:@51635.4]
  assign StickySelects_37_io_ins_3 = io_rPort_8_en_0 & _T_8377; // @[MemPrimitives.scala 122:60:@51636.4]
  assign StickySelects_37_io_ins_4 = io_rPort_11_en_0 & _T_8383; // @[MemPrimitives.scala 122:60:@51637.4]
  assign StickySelects_37_io_ins_5 = io_rPort_12_en_0 & _T_8389; // @[MemPrimitives.scala 122:60:@51638.4]
  assign StickySelects_37_io_ins_6 = io_rPort_14_en_0 & _T_8395; // @[MemPrimitives.scala 122:60:@51639.4]
  assign StickySelects_37_io_ins_7 = io_rPort_18_en_0 & _T_8401; // @[MemPrimitives.scala 122:60:@51640.4]
  assign StickySelects_37_io_ins_8 = io_rPort_20_en_0 & _T_8407; // @[MemPrimitives.scala 122:60:@51641.4]
  assign StickySelects_37_io_ins_9 = io_rPort_21_en_0 & _T_8413; // @[MemPrimitives.scala 122:60:@51642.4]
  assign StickySelects_37_io_ins_10 = io_rPort_23_en_0 & _T_8419; // @[MemPrimitives.scala 122:60:@51643.4]
  assign StickySelects_37_io_ins_11 = io_rPort_24_en_0 & _T_8425; // @[MemPrimitives.scala 122:60:@51644.4]
  assign StickySelects_37_io_ins_12 = io_rPort_25_en_0 & _T_8431; // @[MemPrimitives.scala 122:60:@51645.4]
  assign StickySelects_37_io_ins_13 = io_rPort_27_en_0 & _T_8437; // @[MemPrimitives.scala 122:60:@51646.4]
  assign StickySelects_37_io_ins_14 = io_rPort_28_en_0 & _T_8443; // @[MemPrimitives.scala 122:60:@51647.4]
  assign StickySelects_38_clock = clock; // @[:@51774.4]
  assign StickySelects_38_reset = reset; // @[:@51775.4]
  assign StickySelects_38_io_ins_0 = io_rPort_0_en_0 & _T_8511; // @[MemPrimitives.scala 122:60:@51776.4]
  assign StickySelects_38_io_ins_1 = io_rPort_1_en_0 & _T_8517; // @[MemPrimitives.scala 122:60:@51777.4]
  assign StickySelects_38_io_ins_2 = io_rPort_3_en_0 & _T_8523; // @[MemPrimitives.scala 122:60:@51778.4]
  assign StickySelects_38_io_ins_3 = io_rPort_4_en_0 & _T_8529; // @[MemPrimitives.scala 122:60:@51779.4]
  assign StickySelects_38_io_ins_4 = io_rPort_5_en_0 & _T_8535; // @[MemPrimitives.scala 122:60:@51780.4]
  assign StickySelects_38_io_ins_5 = io_rPort_9_en_0 & _T_8541; // @[MemPrimitives.scala 122:60:@51781.4]
  assign StickySelects_38_io_ins_6 = io_rPort_10_en_0 & _T_8547; // @[MemPrimitives.scala 122:60:@51782.4]
  assign StickySelects_38_io_ins_7 = io_rPort_13_en_0 & _T_8553; // @[MemPrimitives.scala 122:60:@51783.4]
  assign StickySelects_38_io_ins_8 = io_rPort_15_en_0 & _T_8559; // @[MemPrimitives.scala 122:60:@51784.4]
  assign StickySelects_38_io_ins_9 = io_rPort_16_en_0 & _T_8565; // @[MemPrimitives.scala 122:60:@51785.4]
  assign StickySelects_38_io_ins_10 = io_rPort_17_en_0 & _T_8571; // @[MemPrimitives.scala 122:60:@51786.4]
  assign StickySelects_38_io_ins_11 = io_rPort_19_en_0 & _T_8577; // @[MemPrimitives.scala 122:60:@51787.4]
  assign StickySelects_38_io_ins_12 = io_rPort_22_en_0 & _T_8583; // @[MemPrimitives.scala 122:60:@51788.4]
  assign StickySelects_38_io_ins_13 = io_rPort_26_en_0 & _T_8589; // @[MemPrimitives.scala 122:60:@51789.4]
  assign StickySelects_38_io_ins_14 = io_rPort_29_en_0 & _T_8595; // @[MemPrimitives.scala 122:60:@51790.4]
  assign StickySelects_39_clock = clock; // @[:@51917.4]
  assign StickySelects_39_reset = reset; // @[:@51918.4]
  assign StickySelects_39_io_ins_0 = io_rPort_2_en_0 & _T_8663; // @[MemPrimitives.scala 122:60:@51919.4]
  assign StickySelects_39_io_ins_1 = io_rPort_6_en_0 & _T_8669; // @[MemPrimitives.scala 122:60:@51920.4]
  assign StickySelects_39_io_ins_2 = io_rPort_7_en_0 & _T_8675; // @[MemPrimitives.scala 122:60:@51921.4]
  assign StickySelects_39_io_ins_3 = io_rPort_8_en_0 & _T_8681; // @[MemPrimitives.scala 122:60:@51922.4]
  assign StickySelects_39_io_ins_4 = io_rPort_11_en_0 & _T_8687; // @[MemPrimitives.scala 122:60:@51923.4]
  assign StickySelects_39_io_ins_5 = io_rPort_12_en_0 & _T_8693; // @[MemPrimitives.scala 122:60:@51924.4]
  assign StickySelects_39_io_ins_6 = io_rPort_14_en_0 & _T_8699; // @[MemPrimitives.scala 122:60:@51925.4]
  assign StickySelects_39_io_ins_7 = io_rPort_18_en_0 & _T_8705; // @[MemPrimitives.scala 122:60:@51926.4]
  assign StickySelects_39_io_ins_8 = io_rPort_20_en_0 & _T_8711; // @[MemPrimitives.scala 122:60:@51927.4]
  assign StickySelects_39_io_ins_9 = io_rPort_21_en_0 & _T_8717; // @[MemPrimitives.scala 122:60:@51928.4]
  assign StickySelects_39_io_ins_10 = io_rPort_23_en_0 & _T_8723; // @[MemPrimitives.scala 122:60:@51929.4]
  assign StickySelects_39_io_ins_11 = io_rPort_24_en_0 & _T_8729; // @[MemPrimitives.scala 122:60:@51930.4]
  assign StickySelects_39_io_ins_12 = io_rPort_25_en_0 & _T_8735; // @[MemPrimitives.scala 122:60:@51931.4]
  assign StickySelects_39_io_ins_13 = io_rPort_27_en_0 & _T_8741; // @[MemPrimitives.scala 122:60:@51932.4]
  assign StickySelects_39_io_ins_14 = io_rPort_28_en_0 & _T_8747; // @[MemPrimitives.scala 122:60:@51933.4]
  assign RetimeWrapper_clock = clock; // @[:@52061.4]
  assign RetimeWrapper_reset = reset; // @[:@52062.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52064.4]
  assign RetimeWrapper_io_in = _T_2735 & io_rPort_0_en_0; // @[package.scala 94:16:@52063.4]
  assign RetimeWrapper_1_clock = clock; // @[:@52069.4]
  assign RetimeWrapper_1_reset = reset; // @[:@52070.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52072.4]
  assign RetimeWrapper_1_io_in = _T_3039 & io_rPort_0_en_0; // @[package.scala 94:16:@52071.4]
  assign RetimeWrapper_2_clock = clock; // @[:@52077.4]
  assign RetimeWrapper_2_reset = reset; // @[:@52078.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52080.4]
  assign RetimeWrapper_2_io_in = _T_3343 & io_rPort_0_en_0; // @[package.scala 94:16:@52079.4]
  assign RetimeWrapper_3_clock = clock; // @[:@52085.4]
  assign RetimeWrapper_3_reset = reset; // @[:@52086.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52088.4]
  assign RetimeWrapper_3_io_in = _T_3647 & io_rPort_0_en_0; // @[package.scala 94:16:@52087.4]
  assign RetimeWrapper_4_clock = clock; // @[:@52093.4]
  assign RetimeWrapper_4_reset = reset; // @[:@52094.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52096.4]
  assign RetimeWrapper_4_io_in = _T_3951 & io_rPort_0_en_0; // @[package.scala 94:16:@52095.4]
  assign RetimeWrapper_5_clock = clock; // @[:@52101.4]
  assign RetimeWrapper_5_reset = reset; // @[:@52102.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52104.4]
  assign RetimeWrapper_5_io_in = _T_4255 & io_rPort_0_en_0; // @[package.scala 94:16:@52103.4]
  assign RetimeWrapper_6_clock = clock; // @[:@52109.4]
  assign RetimeWrapper_6_reset = reset; // @[:@52110.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52112.4]
  assign RetimeWrapper_6_io_in = _T_4559 & io_rPort_0_en_0; // @[package.scala 94:16:@52111.4]
  assign RetimeWrapper_7_clock = clock; // @[:@52117.4]
  assign RetimeWrapper_7_reset = reset; // @[:@52118.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52120.4]
  assign RetimeWrapper_7_io_in = _T_4863 & io_rPort_0_en_0; // @[package.scala 94:16:@52119.4]
  assign RetimeWrapper_8_clock = clock; // @[:@52125.4]
  assign RetimeWrapper_8_reset = reset; // @[:@52126.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52128.4]
  assign RetimeWrapper_8_io_in = _T_5167 & io_rPort_0_en_0; // @[package.scala 94:16:@52127.4]
  assign RetimeWrapper_9_clock = clock; // @[:@52133.4]
  assign RetimeWrapper_9_reset = reset; // @[:@52134.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52136.4]
  assign RetimeWrapper_9_io_in = _T_5471 & io_rPort_0_en_0; // @[package.scala 94:16:@52135.4]
  assign RetimeWrapper_10_clock = clock; // @[:@52141.4]
  assign RetimeWrapper_10_reset = reset; // @[:@52142.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52144.4]
  assign RetimeWrapper_10_io_in = _T_5775 & io_rPort_0_en_0; // @[package.scala 94:16:@52143.4]
  assign RetimeWrapper_11_clock = clock; // @[:@52149.4]
  assign RetimeWrapper_11_reset = reset; // @[:@52150.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52152.4]
  assign RetimeWrapper_11_io_in = _T_6079 & io_rPort_0_en_0; // @[package.scala 94:16:@52151.4]
  assign RetimeWrapper_12_clock = clock; // @[:@52157.4]
  assign RetimeWrapper_12_reset = reset; // @[:@52158.4]
  assign RetimeWrapper_12_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52160.4]
  assign RetimeWrapper_12_io_in = _T_6383 & io_rPort_0_en_0; // @[package.scala 94:16:@52159.4]
  assign RetimeWrapper_13_clock = clock; // @[:@52165.4]
  assign RetimeWrapper_13_reset = reset; // @[:@52166.4]
  assign RetimeWrapper_13_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52168.4]
  assign RetimeWrapper_13_io_in = _T_6687 & io_rPort_0_en_0; // @[package.scala 94:16:@52167.4]
  assign RetimeWrapper_14_clock = clock; // @[:@52173.4]
  assign RetimeWrapper_14_reset = reset; // @[:@52174.4]
  assign RetimeWrapper_14_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52176.4]
  assign RetimeWrapper_14_io_in = _T_6991 & io_rPort_0_en_0; // @[package.scala 94:16:@52175.4]
  assign RetimeWrapper_15_clock = clock; // @[:@52181.4]
  assign RetimeWrapper_15_reset = reset; // @[:@52182.4]
  assign RetimeWrapper_15_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52184.4]
  assign RetimeWrapper_15_io_in = _T_7295 & io_rPort_0_en_0; // @[package.scala 94:16:@52183.4]
  assign RetimeWrapper_16_clock = clock; // @[:@52189.4]
  assign RetimeWrapper_16_reset = reset; // @[:@52190.4]
  assign RetimeWrapper_16_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52192.4]
  assign RetimeWrapper_16_io_in = _T_7599 & io_rPort_0_en_0; // @[package.scala 94:16:@52191.4]
  assign RetimeWrapper_17_clock = clock; // @[:@52197.4]
  assign RetimeWrapper_17_reset = reset; // @[:@52198.4]
  assign RetimeWrapper_17_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52200.4]
  assign RetimeWrapper_17_io_in = _T_7903 & io_rPort_0_en_0; // @[package.scala 94:16:@52199.4]
  assign RetimeWrapper_18_clock = clock; // @[:@52205.4]
  assign RetimeWrapper_18_reset = reset; // @[:@52206.4]
  assign RetimeWrapper_18_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52208.4]
  assign RetimeWrapper_18_io_in = _T_8207 & io_rPort_0_en_0; // @[package.scala 94:16:@52207.4]
  assign RetimeWrapper_19_clock = clock; // @[:@52213.4]
  assign RetimeWrapper_19_reset = reset; // @[:@52214.4]
  assign RetimeWrapper_19_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@52216.4]
  assign RetimeWrapper_19_io_in = _T_8511 & io_rPort_0_en_0; // @[package.scala 94:16:@52215.4]
  assign RetimeWrapper_20_clock = clock; // @[:@52301.4]
  assign RetimeWrapper_20_reset = reset; // @[:@52302.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52304.4]
  assign RetimeWrapper_20_io_in = _T_2741 & io_rPort_1_en_0; // @[package.scala 94:16:@52303.4]
  assign RetimeWrapper_21_clock = clock; // @[:@52309.4]
  assign RetimeWrapper_21_reset = reset; // @[:@52310.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52312.4]
  assign RetimeWrapper_21_io_in = _T_3045 & io_rPort_1_en_0; // @[package.scala 94:16:@52311.4]
  assign RetimeWrapper_22_clock = clock; // @[:@52317.4]
  assign RetimeWrapper_22_reset = reset; // @[:@52318.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52320.4]
  assign RetimeWrapper_22_io_in = _T_3349 & io_rPort_1_en_0; // @[package.scala 94:16:@52319.4]
  assign RetimeWrapper_23_clock = clock; // @[:@52325.4]
  assign RetimeWrapper_23_reset = reset; // @[:@52326.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52328.4]
  assign RetimeWrapper_23_io_in = _T_3653 & io_rPort_1_en_0; // @[package.scala 94:16:@52327.4]
  assign RetimeWrapper_24_clock = clock; // @[:@52333.4]
  assign RetimeWrapper_24_reset = reset; // @[:@52334.4]
  assign RetimeWrapper_24_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52336.4]
  assign RetimeWrapper_24_io_in = _T_3957 & io_rPort_1_en_0; // @[package.scala 94:16:@52335.4]
  assign RetimeWrapper_25_clock = clock; // @[:@52341.4]
  assign RetimeWrapper_25_reset = reset; // @[:@52342.4]
  assign RetimeWrapper_25_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52344.4]
  assign RetimeWrapper_25_io_in = _T_4261 & io_rPort_1_en_0; // @[package.scala 94:16:@52343.4]
  assign RetimeWrapper_26_clock = clock; // @[:@52349.4]
  assign RetimeWrapper_26_reset = reset; // @[:@52350.4]
  assign RetimeWrapper_26_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52352.4]
  assign RetimeWrapper_26_io_in = _T_4565 & io_rPort_1_en_0; // @[package.scala 94:16:@52351.4]
  assign RetimeWrapper_27_clock = clock; // @[:@52357.4]
  assign RetimeWrapper_27_reset = reset; // @[:@52358.4]
  assign RetimeWrapper_27_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52360.4]
  assign RetimeWrapper_27_io_in = _T_4869 & io_rPort_1_en_0; // @[package.scala 94:16:@52359.4]
  assign RetimeWrapper_28_clock = clock; // @[:@52365.4]
  assign RetimeWrapper_28_reset = reset; // @[:@52366.4]
  assign RetimeWrapper_28_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52368.4]
  assign RetimeWrapper_28_io_in = _T_5173 & io_rPort_1_en_0; // @[package.scala 94:16:@52367.4]
  assign RetimeWrapper_29_clock = clock; // @[:@52373.4]
  assign RetimeWrapper_29_reset = reset; // @[:@52374.4]
  assign RetimeWrapper_29_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52376.4]
  assign RetimeWrapper_29_io_in = _T_5477 & io_rPort_1_en_0; // @[package.scala 94:16:@52375.4]
  assign RetimeWrapper_30_clock = clock; // @[:@52381.4]
  assign RetimeWrapper_30_reset = reset; // @[:@52382.4]
  assign RetimeWrapper_30_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52384.4]
  assign RetimeWrapper_30_io_in = _T_5781 & io_rPort_1_en_0; // @[package.scala 94:16:@52383.4]
  assign RetimeWrapper_31_clock = clock; // @[:@52389.4]
  assign RetimeWrapper_31_reset = reset; // @[:@52390.4]
  assign RetimeWrapper_31_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52392.4]
  assign RetimeWrapper_31_io_in = _T_6085 & io_rPort_1_en_0; // @[package.scala 94:16:@52391.4]
  assign RetimeWrapper_32_clock = clock; // @[:@52397.4]
  assign RetimeWrapper_32_reset = reset; // @[:@52398.4]
  assign RetimeWrapper_32_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52400.4]
  assign RetimeWrapper_32_io_in = _T_6389 & io_rPort_1_en_0; // @[package.scala 94:16:@52399.4]
  assign RetimeWrapper_33_clock = clock; // @[:@52405.4]
  assign RetimeWrapper_33_reset = reset; // @[:@52406.4]
  assign RetimeWrapper_33_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52408.4]
  assign RetimeWrapper_33_io_in = _T_6693 & io_rPort_1_en_0; // @[package.scala 94:16:@52407.4]
  assign RetimeWrapper_34_clock = clock; // @[:@52413.4]
  assign RetimeWrapper_34_reset = reset; // @[:@52414.4]
  assign RetimeWrapper_34_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52416.4]
  assign RetimeWrapper_34_io_in = _T_6997 & io_rPort_1_en_0; // @[package.scala 94:16:@52415.4]
  assign RetimeWrapper_35_clock = clock; // @[:@52421.4]
  assign RetimeWrapper_35_reset = reset; // @[:@52422.4]
  assign RetimeWrapper_35_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52424.4]
  assign RetimeWrapper_35_io_in = _T_7301 & io_rPort_1_en_0; // @[package.scala 94:16:@52423.4]
  assign RetimeWrapper_36_clock = clock; // @[:@52429.4]
  assign RetimeWrapper_36_reset = reset; // @[:@52430.4]
  assign RetimeWrapper_36_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52432.4]
  assign RetimeWrapper_36_io_in = _T_7605 & io_rPort_1_en_0; // @[package.scala 94:16:@52431.4]
  assign RetimeWrapper_37_clock = clock; // @[:@52437.4]
  assign RetimeWrapper_37_reset = reset; // @[:@52438.4]
  assign RetimeWrapper_37_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52440.4]
  assign RetimeWrapper_37_io_in = _T_7909 & io_rPort_1_en_0; // @[package.scala 94:16:@52439.4]
  assign RetimeWrapper_38_clock = clock; // @[:@52445.4]
  assign RetimeWrapper_38_reset = reset; // @[:@52446.4]
  assign RetimeWrapper_38_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52448.4]
  assign RetimeWrapper_38_io_in = _T_8213 & io_rPort_1_en_0; // @[package.scala 94:16:@52447.4]
  assign RetimeWrapper_39_clock = clock; // @[:@52453.4]
  assign RetimeWrapper_39_reset = reset; // @[:@52454.4]
  assign RetimeWrapper_39_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@52456.4]
  assign RetimeWrapper_39_io_in = _T_8517 & io_rPort_1_en_0; // @[package.scala 94:16:@52455.4]
  assign RetimeWrapper_40_clock = clock; // @[:@52541.4]
  assign RetimeWrapper_40_reset = reset; // @[:@52542.4]
  assign RetimeWrapper_40_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52544.4]
  assign RetimeWrapper_40_io_in = _T_2887 & io_rPort_2_en_0; // @[package.scala 94:16:@52543.4]
  assign RetimeWrapper_41_clock = clock; // @[:@52549.4]
  assign RetimeWrapper_41_reset = reset; // @[:@52550.4]
  assign RetimeWrapper_41_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52552.4]
  assign RetimeWrapper_41_io_in = _T_3191 & io_rPort_2_en_0; // @[package.scala 94:16:@52551.4]
  assign RetimeWrapper_42_clock = clock; // @[:@52557.4]
  assign RetimeWrapper_42_reset = reset; // @[:@52558.4]
  assign RetimeWrapper_42_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52560.4]
  assign RetimeWrapper_42_io_in = _T_3495 & io_rPort_2_en_0; // @[package.scala 94:16:@52559.4]
  assign RetimeWrapper_43_clock = clock; // @[:@52565.4]
  assign RetimeWrapper_43_reset = reset; // @[:@52566.4]
  assign RetimeWrapper_43_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52568.4]
  assign RetimeWrapper_43_io_in = _T_3799 & io_rPort_2_en_0; // @[package.scala 94:16:@52567.4]
  assign RetimeWrapper_44_clock = clock; // @[:@52573.4]
  assign RetimeWrapper_44_reset = reset; // @[:@52574.4]
  assign RetimeWrapper_44_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52576.4]
  assign RetimeWrapper_44_io_in = _T_4103 & io_rPort_2_en_0; // @[package.scala 94:16:@52575.4]
  assign RetimeWrapper_45_clock = clock; // @[:@52581.4]
  assign RetimeWrapper_45_reset = reset; // @[:@52582.4]
  assign RetimeWrapper_45_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52584.4]
  assign RetimeWrapper_45_io_in = _T_4407 & io_rPort_2_en_0; // @[package.scala 94:16:@52583.4]
  assign RetimeWrapper_46_clock = clock; // @[:@52589.4]
  assign RetimeWrapper_46_reset = reset; // @[:@52590.4]
  assign RetimeWrapper_46_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52592.4]
  assign RetimeWrapper_46_io_in = _T_4711 & io_rPort_2_en_0; // @[package.scala 94:16:@52591.4]
  assign RetimeWrapper_47_clock = clock; // @[:@52597.4]
  assign RetimeWrapper_47_reset = reset; // @[:@52598.4]
  assign RetimeWrapper_47_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52600.4]
  assign RetimeWrapper_47_io_in = _T_5015 & io_rPort_2_en_0; // @[package.scala 94:16:@52599.4]
  assign RetimeWrapper_48_clock = clock; // @[:@52605.4]
  assign RetimeWrapper_48_reset = reset; // @[:@52606.4]
  assign RetimeWrapper_48_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52608.4]
  assign RetimeWrapper_48_io_in = _T_5319 & io_rPort_2_en_0; // @[package.scala 94:16:@52607.4]
  assign RetimeWrapper_49_clock = clock; // @[:@52613.4]
  assign RetimeWrapper_49_reset = reset; // @[:@52614.4]
  assign RetimeWrapper_49_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52616.4]
  assign RetimeWrapper_49_io_in = _T_5623 & io_rPort_2_en_0; // @[package.scala 94:16:@52615.4]
  assign RetimeWrapper_50_clock = clock; // @[:@52621.4]
  assign RetimeWrapper_50_reset = reset; // @[:@52622.4]
  assign RetimeWrapper_50_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52624.4]
  assign RetimeWrapper_50_io_in = _T_5927 & io_rPort_2_en_0; // @[package.scala 94:16:@52623.4]
  assign RetimeWrapper_51_clock = clock; // @[:@52629.4]
  assign RetimeWrapper_51_reset = reset; // @[:@52630.4]
  assign RetimeWrapper_51_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52632.4]
  assign RetimeWrapper_51_io_in = _T_6231 & io_rPort_2_en_0; // @[package.scala 94:16:@52631.4]
  assign RetimeWrapper_52_clock = clock; // @[:@52637.4]
  assign RetimeWrapper_52_reset = reset; // @[:@52638.4]
  assign RetimeWrapper_52_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52640.4]
  assign RetimeWrapper_52_io_in = _T_6535 & io_rPort_2_en_0; // @[package.scala 94:16:@52639.4]
  assign RetimeWrapper_53_clock = clock; // @[:@52645.4]
  assign RetimeWrapper_53_reset = reset; // @[:@52646.4]
  assign RetimeWrapper_53_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52648.4]
  assign RetimeWrapper_53_io_in = _T_6839 & io_rPort_2_en_0; // @[package.scala 94:16:@52647.4]
  assign RetimeWrapper_54_clock = clock; // @[:@52653.4]
  assign RetimeWrapper_54_reset = reset; // @[:@52654.4]
  assign RetimeWrapper_54_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52656.4]
  assign RetimeWrapper_54_io_in = _T_7143 & io_rPort_2_en_0; // @[package.scala 94:16:@52655.4]
  assign RetimeWrapper_55_clock = clock; // @[:@52661.4]
  assign RetimeWrapper_55_reset = reset; // @[:@52662.4]
  assign RetimeWrapper_55_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52664.4]
  assign RetimeWrapper_55_io_in = _T_7447 & io_rPort_2_en_0; // @[package.scala 94:16:@52663.4]
  assign RetimeWrapper_56_clock = clock; // @[:@52669.4]
  assign RetimeWrapper_56_reset = reset; // @[:@52670.4]
  assign RetimeWrapper_56_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52672.4]
  assign RetimeWrapper_56_io_in = _T_7751 & io_rPort_2_en_0; // @[package.scala 94:16:@52671.4]
  assign RetimeWrapper_57_clock = clock; // @[:@52677.4]
  assign RetimeWrapper_57_reset = reset; // @[:@52678.4]
  assign RetimeWrapper_57_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52680.4]
  assign RetimeWrapper_57_io_in = _T_8055 & io_rPort_2_en_0; // @[package.scala 94:16:@52679.4]
  assign RetimeWrapper_58_clock = clock; // @[:@52685.4]
  assign RetimeWrapper_58_reset = reset; // @[:@52686.4]
  assign RetimeWrapper_58_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52688.4]
  assign RetimeWrapper_58_io_in = _T_8359 & io_rPort_2_en_0; // @[package.scala 94:16:@52687.4]
  assign RetimeWrapper_59_clock = clock; // @[:@52693.4]
  assign RetimeWrapper_59_reset = reset; // @[:@52694.4]
  assign RetimeWrapper_59_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@52696.4]
  assign RetimeWrapper_59_io_in = _T_8663 & io_rPort_2_en_0; // @[package.scala 94:16:@52695.4]
  assign RetimeWrapper_60_clock = clock; // @[:@52781.4]
  assign RetimeWrapper_60_reset = reset; // @[:@52782.4]
  assign RetimeWrapper_60_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52784.4]
  assign RetimeWrapper_60_io_in = _T_2747 & io_rPort_3_en_0; // @[package.scala 94:16:@52783.4]
  assign RetimeWrapper_61_clock = clock; // @[:@52789.4]
  assign RetimeWrapper_61_reset = reset; // @[:@52790.4]
  assign RetimeWrapper_61_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52792.4]
  assign RetimeWrapper_61_io_in = _T_3051 & io_rPort_3_en_0; // @[package.scala 94:16:@52791.4]
  assign RetimeWrapper_62_clock = clock; // @[:@52797.4]
  assign RetimeWrapper_62_reset = reset; // @[:@52798.4]
  assign RetimeWrapper_62_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52800.4]
  assign RetimeWrapper_62_io_in = _T_3355 & io_rPort_3_en_0; // @[package.scala 94:16:@52799.4]
  assign RetimeWrapper_63_clock = clock; // @[:@52805.4]
  assign RetimeWrapper_63_reset = reset; // @[:@52806.4]
  assign RetimeWrapper_63_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52808.4]
  assign RetimeWrapper_63_io_in = _T_3659 & io_rPort_3_en_0; // @[package.scala 94:16:@52807.4]
  assign RetimeWrapper_64_clock = clock; // @[:@52813.4]
  assign RetimeWrapper_64_reset = reset; // @[:@52814.4]
  assign RetimeWrapper_64_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52816.4]
  assign RetimeWrapper_64_io_in = _T_3963 & io_rPort_3_en_0; // @[package.scala 94:16:@52815.4]
  assign RetimeWrapper_65_clock = clock; // @[:@52821.4]
  assign RetimeWrapper_65_reset = reset; // @[:@52822.4]
  assign RetimeWrapper_65_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52824.4]
  assign RetimeWrapper_65_io_in = _T_4267 & io_rPort_3_en_0; // @[package.scala 94:16:@52823.4]
  assign RetimeWrapper_66_clock = clock; // @[:@52829.4]
  assign RetimeWrapper_66_reset = reset; // @[:@52830.4]
  assign RetimeWrapper_66_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52832.4]
  assign RetimeWrapper_66_io_in = _T_4571 & io_rPort_3_en_0; // @[package.scala 94:16:@52831.4]
  assign RetimeWrapper_67_clock = clock; // @[:@52837.4]
  assign RetimeWrapper_67_reset = reset; // @[:@52838.4]
  assign RetimeWrapper_67_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52840.4]
  assign RetimeWrapper_67_io_in = _T_4875 & io_rPort_3_en_0; // @[package.scala 94:16:@52839.4]
  assign RetimeWrapper_68_clock = clock; // @[:@52845.4]
  assign RetimeWrapper_68_reset = reset; // @[:@52846.4]
  assign RetimeWrapper_68_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52848.4]
  assign RetimeWrapper_68_io_in = _T_5179 & io_rPort_3_en_0; // @[package.scala 94:16:@52847.4]
  assign RetimeWrapper_69_clock = clock; // @[:@52853.4]
  assign RetimeWrapper_69_reset = reset; // @[:@52854.4]
  assign RetimeWrapper_69_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52856.4]
  assign RetimeWrapper_69_io_in = _T_5483 & io_rPort_3_en_0; // @[package.scala 94:16:@52855.4]
  assign RetimeWrapper_70_clock = clock; // @[:@52861.4]
  assign RetimeWrapper_70_reset = reset; // @[:@52862.4]
  assign RetimeWrapper_70_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52864.4]
  assign RetimeWrapper_70_io_in = _T_5787 & io_rPort_3_en_0; // @[package.scala 94:16:@52863.4]
  assign RetimeWrapper_71_clock = clock; // @[:@52869.4]
  assign RetimeWrapper_71_reset = reset; // @[:@52870.4]
  assign RetimeWrapper_71_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52872.4]
  assign RetimeWrapper_71_io_in = _T_6091 & io_rPort_3_en_0; // @[package.scala 94:16:@52871.4]
  assign RetimeWrapper_72_clock = clock; // @[:@52877.4]
  assign RetimeWrapper_72_reset = reset; // @[:@52878.4]
  assign RetimeWrapper_72_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52880.4]
  assign RetimeWrapper_72_io_in = _T_6395 & io_rPort_3_en_0; // @[package.scala 94:16:@52879.4]
  assign RetimeWrapper_73_clock = clock; // @[:@52885.4]
  assign RetimeWrapper_73_reset = reset; // @[:@52886.4]
  assign RetimeWrapper_73_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52888.4]
  assign RetimeWrapper_73_io_in = _T_6699 & io_rPort_3_en_0; // @[package.scala 94:16:@52887.4]
  assign RetimeWrapper_74_clock = clock; // @[:@52893.4]
  assign RetimeWrapper_74_reset = reset; // @[:@52894.4]
  assign RetimeWrapper_74_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52896.4]
  assign RetimeWrapper_74_io_in = _T_7003 & io_rPort_3_en_0; // @[package.scala 94:16:@52895.4]
  assign RetimeWrapper_75_clock = clock; // @[:@52901.4]
  assign RetimeWrapper_75_reset = reset; // @[:@52902.4]
  assign RetimeWrapper_75_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52904.4]
  assign RetimeWrapper_75_io_in = _T_7307 & io_rPort_3_en_0; // @[package.scala 94:16:@52903.4]
  assign RetimeWrapper_76_clock = clock; // @[:@52909.4]
  assign RetimeWrapper_76_reset = reset; // @[:@52910.4]
  assign RetimeWrapper_76_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52912.4]
  assign RetimeWrapper_76_io_in = _T_7611 & io_rPort_3_en_0; // @[package.scala 94:16:@52911.4]
  assign RetimeWrapper_77_clock = clock; // @[:@52917.4]
  assign RetimeWrapper_77_reset = reset; // @[:@52918.4]
  assign RetimeWrapper_77_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52920.4]
  assign RetimeWrapper_77_io_in = _T_7915 & io_rPort_3_en_0; // @[package.scala 94:16:@52919.4]
  assign RetimeWrapper_78_clock = clock; // @[:@52925.4]
  assign RetimeWrapper_78_reset = reset; // @[:@52926.4]
  assign RetimeWrapper_78_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52928.4]
  assign RetimeWrapper_78_io_in = _T_8219 & io_rPort_3_en_0; // @[package.scala 94:16:@52927.4]
  assign RetimeWrapper_79_clock = clock; // @[:@52933.4]
  assign RetimeWrapper_79_reset = reset; // @[:@52934.4]
  assign RetimeWrapper_79_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@52936.4]
  assign RetimeWrapper_79_io_in = _T_8523 & io_rPort_3_en_0; // @[package.scala 94:16:@52935.4]
  assign RetimeWrapper_80_clock = clock; // @[:@53021.4]
  assign RetimeWrapper_80_reset = reset; // @[:@53022.4]
  assign RetimeWrapper_80_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53024.4]
  assign RetimeWrapper_80_io_in = _T_2753 & io_rPort_4_en_0; // @[package.scala 94:16:@53023.4]
  assign RetimeWrapper_81_clock = clock; // @[:@53029.4]
  assign RetimeWrapper_81_reset = reset; // @[:@53030.4]
  assign RetimeWrapper_81_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53032.4]
  assign RetimeWrapper_81_io_in = _T_3057 & io_rPort_4_en_0; // @[package.scala 94:16:@53031.4]
  assign RetimeWrapper_82_clock = clock; // @[:@53037.4]
  assign RetimeWrapper_82_reset = reset; // @[:@53038.4]
  assign RetimeWrapper_82_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53040.4]
  assign RetimeWrapper_82_io_in = _T_3361 & io_rPort_4_en_0; // @[package.scala 94:16:@53039.4]
  assign RetimeWrapper_83_clock = clock; // @[:@53045.4]
  assign RetimeWrapper_83_reset = reset; // @[:@53046.4]
  assign RetimeWrapper_83_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53048.4]
  assign RetimeWrapper_83_io_in = _T_3665 & io_rPort_4_en_0; // @[package.scala 94:16:@53047.4]
  assign RetimeWrapper_84_clock = clock; // @[:@53053.4]
  assign RetimeWrapper_84_reset = reset; // @[:@53054.4]
  assign RetimeWrapper_84_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53056.4]
  assign RetimeWrapper_84_io_in = _T_3969 & io_rPort_4_en_0; // @[package.scala 94:16:@53055.4]
  assign RetimeWrapper_85_clock = clock; // @[:@53061.4]
  assign RetimeWrapper_85_reset = reset; // @[:@53062.4]
  assign RetimeWrapper_85_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53064.4]
  assign RetimeWrapper_85_io_in = _T_4273 & io_rPort_4_en_0; // @[package.scala 94:16:@53063.4]
  assign RetimeWrapper_86_clock = clock; // @[:@53069.4]
  assign RetimeWrapper_86_reset = reset; // @[:@53070.4]
  assign RetimeWrapper_86_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53072.4]
  assign RetimeWrapper_86_io_in = _T_4577 & io_rPort_4_en_0; // @[package.scala 94:16:@53071.4]
  assign RetimeWrapper_87_clock = clock; // @[:@53077.4]
  assign RetimeWrapper_87_reset = reset; // @[:@53078.4]
  assign RetimeWrapper_87_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53080.4]
  assign RetimeWrapper_87_io_in = _T_4881 & io_rPort_4_en_0; // @[package.scala 94:16:@53079.4]
  assign RetimeWrapper_88_clock = clock; // @[:@53085.4]
  assign RetimeWrapper_88_reset = reset; // @[:@53086.4]
  assign RetimeWrapper_88_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53088.4]
  assign RetimeWrapper_88_io_in = _T_5185 & io_rPort_4_en_0; // @[package.scala 94:16:@53087.4]
  assign RetimeWrapper_89_clock = clock; // @[:@53093.4]
  assign RetimeWrapper_89_reset = reset; // @[:@53094.4]
  assign RetimeWrapper_89_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53096.4]
  assign RetimeWrapper_89_io_in = _T_5489 & io_rPort_4_en_0; // @[package.scala 94:16:@53095.4]
  assign RetimeWrapper_90_clock = clock; // @[:@53101.4]
  assign RetimeWrapper_90_reset = reset; // @[:@53102.4]
  assign RetimeWrapper_90_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53104.4]
  assign RetimeWrapper_90_io_in = _T_5793 & io_rPort_4_en_0; // @[package.scala 94:16:@53103.4]
  assign RetimeWrapper_91_clock = clock; // @[:@53109.4]
  assign RetimeWrapper_91_reset = reset; // @[:@53110.4]
  assign RetimeWrapper_91_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53112.4]
  assign RetimeWrapper_91_io_in = _T_6097 & io_rPort_4_en_0; // @[package.scala 94:16:@53111.4]
  assign RetimeWrapper_92_clock = clock; // @[:@53117.4]
  assign RetimeWrapper_92_reset = reset; // @[:@53118.4]
  assign RetimeWrapper_92_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53120.4]
  assign RetimeWrapper_92_io_in = _T_6401 & io_rPort_4_en_0; // @[package.scala 94:16:@53119.4]
  assign RetimeWrapper_93_clock = clock; // @[:@53125.4]
  assign RetimeWrapper_93_reset = reset; // @[:@53126.4]
  assign RetimeWrapper_93_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53128.4]
  assign RetimeWrapper_93_io_in = _T_6705 & io_rPort_4_en_0; // @[package.scala 94:16:@53127.4]
  assign RetimeWrapper_94_clock = clock; // @[:@53133.4]
  assign RetimeWrapper_94_reset = reset; // @[:@53134.4]
  assign RetimeWrapper_94_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53136.4]
  assign RetimeWrapper_94_io_in = _T_7009 & io_rPort_4_en_0; // @[package.scala 94:16:@53135.4]
  assign RetimeWrapper_95_clock = clock; // @[:@53141.4]
  assign RetimeWrapper_95_reset = reset; // @[:@53142.4]
  assign RetimeWrapper_95_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53144.4]
  assign RetimeWrapper_95_io_in = _T_7313 & io_rPort_4_en_0; // @[package.scala 94:16:@53143.4]
  assign RetimeWrapper_96_clock = clock; // @[:@53149.4]
  assign RetimeWrapper_96_reset = reset; // @[:@53150.4]
  assign RetimeWrapper_96_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53152.4]
  assign RetimeWrapper_96_io_in = _T_7617 & io_rPort_4_en_0; // @[package.scala 94:16:@53151.4]
  assign RetimeWrapper_97_clock = clock; // @[:@53157.4]
  assign RetimeWrapper_97_reset = reset; // @[:@53158.4]
  assign RetimeWrapper_97_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53160.4]
  assign RetimeWrapper_97_io_in = _T_7921 & io_rPort_4_en_0; // @[package.scala 94:16:@53159.4]
  assign RetimeWrapper_98_clock = clock; // @[:@53165.4]
  assign RetimeWrapper_98_reset = reset; // @[:@53166.4]
  assign RetimeWrapper_98_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53168.4]
  assign RetimeWrapper_98_io_in = _T_8225 & io_rPort_4_en_0; // @[package.scala 94:16:@53167.4]
  assign RetimeWrapper_99_clock = clock; // @[:@53173.4]
  assign RetimeWrapper_99_reset = reset; // @[:@53174.4]
  assign RetimeWrapper_99_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@53176.4]
  assign RetimeWrapper_99_io_in = _T_8529 & io_rPort_4_en_0; // @[package.scala 94:16:@53175.4]
  assign RetimeWrapper_100_clock = clock; // @[:@53261.4]
  assign RetimeWrapper_100_reset = reset; // @[:@53262.4]
  assign RetimeWrapper_100_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53264.4]
  assign RetimeWrapper_100_io_in = _T_2759 & io_rPort_5_en_0; // @[package.scala 94:16:@53263.4]
  assign RetimeWrapper_101_clock = clock; // @[:@53269.4]
  assign RetimeWrapper_101_reset = reset; // @[:@53270.4]
  assign RetimeWrapper_101_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53272.4]
  assign RetimeWrapper_101_io_in = _T_3063 & io_rPort_5_en_0; // @[package.scala 94:16:@53271.4]
  assign RetimeWrapper_102_clock = clock; // @[:@53277.4]
  assign RetimeWrapper_102_reset = reset; // @[:@53278.4]
  assign RetimeWrapper_102_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53280.4]
  assign RetimeWrapper_102_io_in = _T_3367 & io_rPort_5_en_0; // @[package.scala 94:16:@53279.4]
  assign RetimeWrapper_103_clock = clock; // @[:@53285.4]
  assign RetimeWrapper_103_reset = reset; // @[:@53286.4]
  assign RetimeWrapper_103_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53288.4]
  assign RetimeWrapper_103_io_in = _T_3671 & io_rPort_5_en_0; // @[package.scala 94:16:@53287.4]
  assign RetimeWrapper_104_clock = clock; // @[:@53293.4]
  assign RetimeWrapper_104_reset = reset; // @[:@53294.4]
  assign RetimeWrapper_104_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53296.4]
  assign RetimeWrapper_104_io_in = _T_3975 & io_rPort_5_en_0; // @[package.scala 94:16:@53295.4]
  assign RetimeWrapper_105_clock = clock; // @[:@53301.4]
  assign RetimeWrapper_105_reset = reset; // @[:@53302.4]
  assign RetimeWrapper_105_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53304.4]
  assign RetimeWrapper_105_io_in = _T_4279 & io_rPort_5_en_0; // @[package.scala 94:16:@53303.4]
  assign RetimeWrapper_106_clock = clock; // @[:@53309.4]
  assign RetimeWrapper_106_reset = reset; // @[:@53310.4]
  assign RetimeWrapper_106_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53312.4]
  assign RetimeWrapper_106_io_in = _T_4583 & io_rPort_5_en_0; // @[package.scala 94:16:@53311.4]
  assign RetimeWrapper_107_clock = clock; // @[:@53317.4]
  assign RetimeWrapper_107_reset = reset; // @[:@53318.4]
  assign RetimeWrapper_107_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53320.4]
  assign RetimeWrapper_107_io_in = _T_4887 & io_rPort_5_en_0; // @[package.scala 94:16:@53319.4]
  assign RetimeWrapper_108_clock = clock; // @[:@53325.4]
  assign RetimeWrapper_108_reset = reset; // @[:@53326.4]
  assign RetimeWrapper_108_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53328.4]
  assign RetimeWrapper_108_io_in = _T_5191 & io_rPort_5_en_0; // @[package.scala 94:16:@53327.4]
  assign RetimeWrapper_109_clock = clock; // @[:@53333.4]
  assign RetimeWrapper_109_reset = reset; // @[:@53334.4]
  assign RetimeWrapper_109_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53336.4]
  assign RetimeWrapper_109_io_in = _T_5495 & io_rPort_5_en_0; // @[package.scala 94:16:@53335.4]
  assign RetimeWrapper_110_clock = clock; // @[:@53341.4]
  assign RetimeWrapper_110_reset = reset; // @[:@53342.4]
  assign RetimeWrapper_110_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53344.4]
  assign RetimeWrapper_110_io_in = _T_5799 & io_rPort_5_en_0; // @[package.scala 94:16:@53343.4]
  assign RetimeWrapper_111_clock = clock; // @[:@53349.4]
  assign RetimeWrapper_111_reset = reset; // @[:@53350.4]
  assign RetimeWrapper_111_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53352.4]
  assign RetimeWrapper_111_io_in = _T_6103 & io_rPort_5_en_0; // @[package.scala 94:16:@53351.4]
  assign RetimeWrapper_112_clock = clock; // @[:@53357.4]
  assign RetimeWrapper_112_reset = reset; // @[:@53358.4]
  assign RetimeWrapper_112_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53360.4]
  assign RetimeWrapper_112_io_in = _T_6407 & io_rPort_5_en_0; // @[package.scala 94:16:@53359.4]
  assign RetimeWrapper_113_clock = clock; // @[:@53365.4]
  assign RetimeWrapper_113_reset = reset; // @[:@53366.4]
  assign RetimeWrapper_113_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53368.4]
  assign RetimeWrapper_113_io_in = _T_6711 & io_rPort_5_en_0; // @[package.scala 94:16:@53367.4]
  assign RetimeWrapper_114_clock = clock; // @[:@53373.4]
  assign RetimeWrapper_114_reset = reset; // @[:@53374.4]
  assign RetimeWrapper_114_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53376.4]
  assign RetimeWrapper_114_io_in = _T_7015 & io_rPort_5_en_0; // @[package.scala 94:16:@53375.4]
  assign RetimeWrapper_115_clock = clock; // @[:@53381.4]
  assign RetimeWrapper_115_reset = reset; // @[:@53382.4]
  assign RetimeWrapper_115_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53384.4]
  assign RetimeWrapper_115_io_in = _T_7319 & io_rPort_5_en_0; // @[package.scala 94:16:@53383.4]
  assign RetimeWrapper_116_clock = clock; // @[:@53389.4]
  assign RetimeWrapper_116_reset = reset; // @[:@53390.4]
  assign RetimeWrapper_116_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53392.4]
  assign RetimeWrapper_116_io_in = _T_7623 & io_rPort_5_en_0; // @[package.scala 94:16:@53391.4]
  assign RetimeWrapper_117_clock = clock; // @[:@53397.4]
  assign RetimeWrapper_117_reset = reset; // @[:@53398.4]
  assign RetimeWrapper_117_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53400.4]
  assign RetimeWrapper_117_io_in = _T_7927 & io_rPort_5_en_0; // @[package.scala 94:16:@53399.4]
  assign RetimeWrapper_118_clock = clock; // @[:@53405.4]
  assign RetimeWrapper_118_reset = reset; // @[:@53406.4]
  assign RetimeWrapper_118_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53408.4]
  assign RetimeWrapper_118_io_in = _T_8231 & io_rPort_5_en_0; // @[package.scala 94:16:@53407.4]
  assign RetimeWrapper_119_clock = clock; // @[:@53413.4]
  assign RetimeWrapper_119_reset = reset; // @[:@53414.4]
  assign RetimeWrapper_119_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@53416.4]
  assign RetimeWrapper_119_io_in = _T_8535 & io_rPort_5_en_0; // @[package.scala 94:16:@53415.4]
  assign RetimeWrapper_120_clock = clock; // @[:@53501.4]
  assign RetimeWrapper_120_reset = reset; // @[:@53502.4]
  assign RetimeWrapper_120_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53504.4]
  assign RetimeWrapper_120_io_in = _T_2893 & io_rPort_6_en_0; // @[package.scala 94:16:@53503.4]
  assign RetimeWrapper_121_clock = clock; // @[:@53509.4]
  assign RetimeWrapper_121_reset = reset; // @[:@53510.4]
  assign RetimeWrapper_121_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53512.4]
  assign RetimeWrapper_121_io_in = _T_3197 & io_rPort_6_en_0; // @[package.scala 94:16:@53511.4]
  assign RetimeWrapper_122_clock = clock; // @[:@53517.4]
  assign RetimeWrapper_122_reset = reset; // @[:@53518.4]
  assign RetimeWrapper_122_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53520.4]
  assign RetimeWrapper_122_io_in = _T_3501 & io_rPort_6_en_0; // @[package.scala 94:16:@53519.4]
  assign RetimeWrapper_123_clock = clock; // @[:@53525.4]
  assign RetimeWrapper_123_reset = reset; // @[:@53526.4]
  assign RetimeWrapper_123_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53528.4]
  assign RetimeWrapper_123_io_in = _T_3805 & io_rPort_6_en_0; // @[package.scala 94:16:@53527.4]
  assign RetimeWrapper_124_clock = clock; // @[:@53533.4]
  assign RetimeWrapper_124_reset = reset; // @[:@53534.4]
  assign RetimeWrapper_124_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53536.4]
  assign RetimeWrapper_124_io_in = _T_4109 & io_rPort_6_en_0; // @[package.scala 94:16:@53535.4]
  assign RetimeWrapper_125_clock = clock; // @[:@53541.4]
  assign RetimeWrapper_125_reset = reset; // @[:@53542.4]
  assign RetimeWrapper_125_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53544.4]
  assign RetimeWrapper_125_io_in = _T_4413 & io_rPort_6_en_0; // @[package.scala 94:16:@53543.4]
  assign RetimeWrapper_126_clock = clock; // @[:@53549.4]
  assign RetimeWrapper_126_reset = reset; // @[:@53550.4]
  assign RetimeWrapper_126_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53552.4]
  assign RetimeWrapper_126_io_in = _T_4717 & io_rPort_6_en_0; // @[package.scala 94:16:@53551.4]
  assign RetimeWrapper_127_clock = clock; // @[:@53557.4]
  assign RetimeWrapper_127_reset = reset; // @[:@53558.4]
  assign RetimeWrapper_127_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53560.4]
  assign RetimeWrapper_127_io_in = _T_5021 & io_rPort_6_en_0; // @[package.scala 94:16:@53559.4]
  assign RetimeWrapper_128_clock = clock; // @[:@53565.4]
  assign RetimeWrapper_128_reset = reset; // @[:@53566.4]
  assign RetimeWrapper_128_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53568.4]
  assign RetimeWrapper_128_io_in = _T_5325 & io_rPort_6_en_0; // @[package.scala 94:16:@53567.4]
  assign RetimeWrapper_129_clock = clock; // @[:@53573.4]
  assign RetimeWrapper_129_reset = reset; // @[:@53574.4]
  assign RetimeWrapper_129_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53576.4]
  assign RetimeWrapper_129_io_in = _T_5629 & io_rPort_6_en_0; // @[package.scala 94:16:@53575.4]
  assign RetimeWrapper_130_clock = clock; // @[:@53581.4]
  assign RetimeWrapper_130_reset = reset; // @[:@53582.4]
  assign RetimeWrapper_130_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53584.4]
  assign RetimeWrapper_130_io_in = _T_5933 & io_rPort_6_en_0; // @[package.scala 94:16:@53583.4]
  assign RetimeWrapper_131_clock = clock; // @[:@53589.4]
  assign RetimeWrapper_131_reset = reset; // @[:@53590.4]
  assign RetimeWrapper_131_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53592.4]
  assign RetimeWrapper_131_io_in = _T_6237 & io_rPort_6_en_0; // @[package.scala 94:16:@53591.4]
  assign RetimeWrapper_132_clock = clock; // @[:@53597.4]
  assign RetimeWrapper_132_reset = reset; // @[:@53598.4]
  assign RetimeWrapper_132_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53600.4]
  assign RetimeWrapper_132_io_in = _T_6541 & io_rPort_6_en_0; // @[package.scala 94:16:@53599.4]
  assign RetimeWrapper_133_clock = clock; // @[:@53605.4]
  assign RetimeWrapper_133_reset = reset; // @[:@53606.4]
  assign RetimeWrapper_133_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53608.4]
  assign RetimeWrapper_133_io_in = _T_6845 & io_rPort_6_en_0; // @[package.scala 94:16:@53607.4]
  assign RetimeWrapper_134_clock = clock; // @[:@53613.4]
  assign RetimeWrapper_134_reset = reset; // @[:@53614.4]
  assign RetimeWrapper_134_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53616.4]
  assign RetimeWrapper_134_io_in = _T_7149 & io_rPort_6_en_0; // @[package.scala 94:16:@53615.4]
  assign RetimeWrapper_135_clock = clock; // @[:@53621.4]
  assign RetimeWrapper_135_reset = reset; // @[:@53622.4]
  assign RetimeWrapper_135_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53624.4]
  assign RetimeWrapper_135_io_in = _T_7453 & io_rPort_6_en_0; // @[package.scala 94:16:@53623.4]
  assign RetimeWrapper_136_clock = clock; // @[:@53629.4]
  assign RetimeWrapper_136_reset = reset; // @[:@53630.4]
  assign RetimeWrapper_136_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53632.4]
  assign RetimeWrapper_136_io_in = _T_7757 & io_rPort_6_en_0; // @[package.scala 94:16:@53631.4]
  assign RetimeWrapper_137_clock = clock; // @[:@53637.4]
  assign RetimeWrapper_137_reset = reset; // @[:@53638.4]
  assign RetimeWrapper_137_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53640.4]
  assign RetimeWrapper_137_io_in = _T_8061 & io_rPort_6_en_0; // @[package.scala 94:16:@53639.4]
  assign RetimeWrapper_138_clock = clock; // @[:@53645.4]
  assign RetimeWrapper_138_reset = reset; // @[:@53646.4]
  assign RetimeWrapper_138_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53648.4]
  assign RetimeWrapper_138_io_in = _T_8365 & io_rPort_6_en_0; // @[package.scala 94:16:@53647.4]
  assign RetimeWrapper_139_clock = clock; // @[:@53653.4]
  assign RetimeWrapper_139_reset = reset; // @[:@53654.4]
  assign RetimeWrapper_139_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@53656.4]
  assign RetimeWrapper_139_io_in = _T_8669 & io_rPort_6_en_0; // @[package.scala 94:16:@53655.4]
  assign RetimeWrapper_140_clock = clock; // @[:@53741.4]
  assign RetimeWrapper_140_reset = reset; // @[:@53742.4]
  assign RetimeWrapper_140_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53744.4]
  assign RetimeWrapper_140_io_in = _T_2899 & io_rPort_7_en_0; // @[package.scala 94:16:@53743.4]
  assign RetimeWrapper_141_clock = clock; // @[:@53749.4]
  assign RetimeWrapper_141_reset = reset; // @[:@53750.4]
  assign RetimeWrapper_141_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53752.4]
  assign RetimeWrapper_141_io_in = _T_3203 & io_rPort_7_en_0; // @[package.scala 94:16:@53751.4]
  assign RetimeWrapper_142_clock = clock; // @[:@53757.4]
  assign RetimeWrapper_142_reset = reset; // @[:@53758.4]
  assign RetimeWrapper_142_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53760.4]
  assign RetimeWrapper_142_io_in = _T_3507 & io_rPort_7_en_0; // @[package.scala 94:16:@53759.4]
  assign RetimeWrapper_143_clock = clock; // @[:@53765.4]
  assign RetimeWrapper_143_reset = reset; // @[:@53766.4]
  assign RetimeWrapper_143_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53768.4]
  assign RetimeWrapper_143_io_in = _T_3811 & io_rPort_7_en_0; // @[package.scala 94:16:@53767.4]
  assign RetimeWrapper_144_clock = clock; // @[:@53773.4]
  assign RetimeWrapper_144_reset = reset; // @[:@53774.4]
  assign RetimeWrapper_144_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53776.4]
  assign RetimeWrapper_144_io_in = _T_4115 & io_rPort_7_en_0; // @[package.scala 94:16:@53775.4]
  assign RetimeWrapper_145_clock = clock; // @[:@53781.4]
  assign RetimeWrapper_145_reset = reset; // @[:@53782.4]
  assign RetimeWrapper_145_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53784.4]
  assign RetimeWrapper_145_io_in = _T_4419 & io_rPort_7_en_0; // @[package.scala 94:16:@53783.4]
  assign RetimeWrapper_146_clock = clock; // @[:@53789.4]
  assign RetimeWrapper_146_reset = reset; // @[:@53790.4]
  assign RetimeWrapper_146_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53792.4]
  assign RetimeWrapper_146_io_in = _T_4723 & io_rPort_7_en_0; // @[package.scala 94:16:@53791.4]
  assign RetimeWrapper_147_clock = clock; // @[:@53797.4]
  assign RetimeWrapper_147_reset = reset; // @[:@53798.4]
  assign RetimeWrapper_147_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53800.4]
  assign RetimeWrapper_147_io_in = _T_5027 & io_rPort_7_en_0; // @[package.scala 94:16:@53799.4]
  assign RetimeWrapper_148_clock = clock; // @[:@53805.4]
  assign RetimeWrapper_148_reset = reset; // @[:@53806.4]
  assign RetimeWrapper_148_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53808.4]
  assign RetimeWrapper_148_io_in = _T_5331 & io_rPort_7_en_0; // @[package.scala 94:16:@53807.4]
  assign RetimeWrapper_149_clock = clock; // @[:@53813.4]
  assign RetimeWrapper_149_reset = reset; // @[:@53814.4]
  assign RetimeWrapper_149_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53816.4]
  assign RetimeWrapper_149_io_in = _T_5635 & io_rPort_7_en_0; // @[package.scala 94:16:@53815.4]
  assign RetimeWrapper_150_clock = clock; // @[:@53821.4]
  assign RetimeWrapper_150_reset = reset; // @[:@53822.4]
  assign RetimeWrapper_150_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53824.4]
  assign RetimeWrapper_150_io_in = _T_5939 & io_rPort_7_en_0; // @[package.scala 94:16:@53823.4]
  assign RetimeWrapper_151_clock = clock; // @[:@53829.4]
  assign RetimeWrapper_151_reset = reset; // @[:@53830.4]
  assign RetimeWrapper_151_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53832.4]
  assign RetimeWrapper_151_io_in = _T_6243 & io_rPort_7_en_0; // @[package.scala 94:16:@53831.4]
  assign RetimeWrapper_152_clock = clock; // @[:@53837.4]
  assign RetimeWrapper_152_reset = reset; // @[:@53838.4]
  assign RetimeWrapper_152_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53840.4]
  assign RetimeWrapper_152_io_in = _T_6547 & io_rPort_7_en_0; // @[package.scala 94:16:@53839.4]
  assign RetimeWrapper_153_clock = clock; // @[:@53845.4]
  assign RetimeWrapper_153_reset = reset; // @[:@53846.4]
  assign RetimeWrapper_153_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53848.4]
  assign RetimeWrapper_153_io_in = _T_6851 & io_rPort_7_en_0; // @[package.scala 94:16:@53847.4]
  assign RetimeWrapper_154_clock = clock; // @[:@53853.4]
  assign RetimeWrapper_154_reset = reset; // @[:@53854.4]
  assign RetimeWrapper_154_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53856.4]
  assign RetimeWrapper_154_io_in = _T_7155 & io_rPort_7_en_0; // @[package.scala 94:16:@53855.4]
  assign RetimeWrapper_155_clock = clock; // @[:@53861.4]
  assign RetimeWrapper_155_reset = reset; // @[:@53862.4]
  assign RetimeWrapper_155_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53864.4]
  assign RetimeWrapper_155_io_in = _T_7459 & io_rPort_7_en_0; // @[package.scala 94:16:@53863.4]
  assign RetimeWrapper_156_clock = clock; // @[:@53869.4]
  assign RetimeWrapper_156_reset = reset; // @[:@53870.4]
  assign RetimeWrapper_156_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53872.4]
  assign RetimeWrapper_156_io_in = _T_7763 & io_rPort_7_en_0; // @[package.scala 94:16:@53871.4]
  assign RetimeWrapper_157_clock = clock; // @[:@53877.4]
  assign RetimeWrapper_157_reset = reset; // @[:@53878.4]
  assign RetimeWrapper_157_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53880.4]
  assign RetimeWrapper_157_io_in = _T_8067 & io_rPort_7_en_0; // @[package.scala 94:16:@53879.4]
  assign RetimeWrapper_158_clock = clock; // @[:@53885.4]
  assign RetimeWrapper_158_reset = reset; // @[:@53886.4]
  assign RetimeWrapper_158_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53888.4]
  assign RetimeWrapper_158_io_in = _T_8371 & io_rPort_7_en_0; // @[package.scala 94:16:@53887.4]
  assign RetimeWrapper_159_clock = clock; // @[:@53893.4]
  assign RetimeWrapper_159_reset = reset; // @[:@53894.4]
  assign RetimeWrapper_159_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@53896.4]
  assign RetimeWrapper_159_io_in = _T_8675 & io_rPort_7_en_0; // @[package.scala 94:16:@53895.4]
  assign RetimeWrapper_160_clock = clock; // @[:@53981.4]
  assign RetimeWrapper_160_reset = reset; // @[:@53982.4]
  assign RetimeWrapper_160_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@53984.4]
  assign RetimeWrapper_160_io_in = _T_2905 & io_rPort_8_en_0; // @[package.scala 94:16:@53983.4]
  assign RetimeWrapper_161_clock = clock; // @[:@53989.4]
  assign RetimeWrapper_161_reset = reset; // @[:@53990.4]
  assign RetimeWrapper_161_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@53992.4]
  assign RetimeWrapper_161_io_in = _T_3209 & io_rPort_8_en_0; // @[package.scala 94:16:@53991.4]
  assign RetimeWrapper_162_clock = clock; // @[:@53997.4]
  assign RetimeWrapper_162_reset = reset; // @[:@53998.4]
  assign RetimeWrapper_162_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54000.4]
  assign RetimeWrapper_162_io_in = _T_3513 & io_rPort_8_en_0; // @[package.scala 94:16:@53999.4]
  assign RetimeWrapper_163_clock = clock; // @[:@54005.4]
  assign RetimeWrapper_163_reset = reset; // @[:@54006.4]
  assign RetimeWrapper_163_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54008.4]
  assign RetimeWrapper_163_io_in = _T_3817 & io_rPort_8_en_0; // @[package.scala 94:16:@54007.4]
  assign RetimeWrapper_164_clock = clock; // @[:@54013.4]
  assign RetimeWrapper_164_reset = reset; // @[:@54014.4]
  assign RetimeWrapper_164_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54016.4]
  assign RetimeWrapper_164_io_in = _T_4121 & io_rPort_8_en_0; // @[package.scala 94:16:@54015.4]
  assign RetimeWrapper_165_clock = clock; // @[:@54021.4]
  assign RetimeWrapper_165_reset = reset; // @[:@54022.4]
  assign RetimeWrapper_165_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54024.4]
  assign RetimeWrapper_165_io_in = _T_4425 & io_rPort_8_en_0; // @[package.scala 94:16:@54023.4]
  assign RetimeWrapper_166_clock = clock; // @[:@54029.4]
  assign RetimeWrapper_166_reset = reset; // @[:@54030.4]
  assign RetimeWrapper_166_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54032.4]
  assign RetimeWrapper_166_io_in = _T_4729 & io_rPort_8_en_0; // @[package.scala 94:16:@54031.4]
  assign RetimeWrapper_167_clock = clock; // @[:@54037.4]
  assign RetimeWrapper_167_reset = reset; // @[:@54038.4]
  assign RetimeWrapper_167_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54040.4]
  assign RetimeWrapper_167_io_in = _T_5033 & io_rPort_8_en_0; // @[package.scala 94:16:@54039.4]
  assign RetimeWrapper_168_clock = clock; // @[:@54045.4]
  assign RetimeWrapper_168_reset = reset; // @[:@54046.4]
  assign RetimeWrapper_168_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54048.4]
  assign RetimeWrapper_168_io_in = _T_5337 & io_rPort_8_en_0; // @[package.scala 94:16:@54047.4]
  assign RetimeWrapper_169_clock = clock; // @[:@54053.4]
  assign RetimeWrapper_169_reset = reset; // @[:@54054.4]
  assign RetimeWrapper_169_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54056.4]
  assign RetimeWrapper_169_io_in = _T_5641 & io_rPort_8_en_0; // @[package.scala 94:16:@54055.4]
  assign RetimeWrapper_170_clock = clock; // @[:@54061.4]
  assign RetimeWrapper_170_reset = reset; // @[:@54062.4]
  assign RetimeWrapper_170_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54064.4]
  assign RetimeWrapper_170_io_in = _T_5945 & io_rPort_8_en_0; // @[package.scala 94:16:@54063.4]
  assign RetimeWrapper_171_clock = clock; // @[:@54069.4]
  assign RetimeWrapper_171_reset = reset; // @[:@54070.4]
  assign RetimeWrapper_171_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54072.4]
  assign RetimeWrapper_171_io_in = _T_6249 & io_rPort_8_en_0; // @[package.scala 94:16:@54071.4]
  assign RetimeWrapper_172_clock = clock; // @[:@54077.4]
  assign RetimeWrapper_172_reset = reset; // @[:@54078.4]
  assign RetimeWrapper_172_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54080.4]
  assign RetimeWrapper_172_io_in = _T_6553 & io_rPort_8_en_0; // @[package.scala 94:16:@54079.4]
  assign RetimeWrapper_173_clock = clock; // @[:@54085.4]
  assign RetimeWrapper_173_reset = reset; // @[:@54086.4]
  assign RetimeWrapper_173_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54088.4]
  assign RetimeWrapper_173_io_in = _T_6857 & io_rPort_8_en_0; // @[package.scala 94:16:@54087.4]
  assign RetimeWrapper_174_clock = clock; // @[:@54093.4]
  assign RetimeWrapper_174_reset = reset; // @[:@54094.4]
  assign RetimeWrapper_174_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54096.4]
  assign RetimeWrapper_174_io_in = _T_7161 & io_rPort_8_en_0; // @[package.scala 94:16:@54095.4]
  assign RetimeWrapper_175_clock = clock; // @[:@54101.4]
  assign RetimeWrapper_175_reset = reset; // @[:@54102.4]
  assign RetimeWrapper_175_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54104.4]
  assign RetimeWrapper_175_io_in = _T_7465 & io_rPort_8_en_0; // @[package.scala 94:16:@54103.4]
  assign RetimeWrapper_176_clock = clock; // @[:@54109.4]
  assign RetimeWrapper_176_reset = reset; // @[:@54110.4]
  assign RetimeWrapper_176_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54112.4]
  assign RetimeWrapper_176_io_in = _T_7769 & io_rPort_8_en_0; // @[package.scala 94:16:@54111.4]
  assign RetimeWrapper_177_clock = clock; // @[:@54117.4]
  assign RetimeWrapper_177_reset = reset; // @[:@54118.4]
  assign RetimeWrapper_177_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54120.4]
  assign RetimeWrapper_177_io_in = _T_8073 & io_rPort_8_en_0; // @[package.scala 94:16:@54119.4]
  assign RetimeWrapper_178_clock = clock; // @[:@54125.4]
  assign RetimeWrapper_178_reset = reset; // @[:@54126.4]
  assign RetimeWrapper_178_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54128.4]
  assign RetimeWrapper_178_io_in = _T_8377 & io_rPort_8_en_0; // @[package.scala 94:16:@54127.4]
  assign RetimeWrapper_179_clock = clock; // @[:@54133.4]
  assign RetimeWrapper_179_reset = reset; // @[:@54134.4]
  assign RetimeWrapper_179_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@54136.4]
  assign RetimeWrapper_179_io_in = _T_8681 & io_rPort_8_en_0; // @[package.scala 94:16:@54135.4]
  assign RetimeWrapper_180_clock = clock; // @[:@54221.4]
  assign RetimeWrapper_180_reset = reset; // @[:@54222.4]
  assign RetimeWrapper_180_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54224.4]
  assign RetimeWrapper_180_io_in = _T_2765 & io_rPort_9_en_0; // @[package.scala 94:16:@54223.4]
  assign RetimeWrapper_181_clock = clock; // @[:@54229.4]
  assign RetimeWrapper_181_reset = reset; // @[:@54230.4]
  assign RetimeWrapper_181_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54232.4]
  assign RetimeWrapper_181_io_in = _T_3069 & io_rPort_9_en_0; // @[package.scala 94:16:@54231.4]
  assign RetimeWrapper_182_clock = clock; // @[:@54237.4]
  assign RetimeWrapper_182_reset = reset; // @[:@54238.4]
  assign RetimeWrapper_182_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54240.4]
  assign RetimeWrapper_182_io_in = _T_3373 & io_rPort_9_en_0; // @[package.scala 94:16:@54239.4]
  assign RetimeWrapper_183_clock = clock; // @[:@54245.4]
  assign RetimeWrapper_183_reset = reset; // @[:@54246.4]
  assign RetimeWrapper_183_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54248.4]
  assign RetimeWrapper_183_io_in = _T_3677 & io_rPort_9_en_0; // @[package.scala 94:16:@54247.4]
  assign RetimeWrapper_184_clock = clock; // @[:@54253.4]
  assign RetimeWrapper_184_reset = reset; // @[:@54254.4]
  assign RetimeWrapper_184_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54256.4]
  assign RetimeWrapper_184_io_in = _T_3981 & io_rPort_9_en_0; // @[package.scala 94:16:@54255.4]
  assign RetimeWrapper_185_clock = clock; // @[:@54261.4]
  assign RetimeWrapper_185_reset = reset; // @[:@54262.4]
  assign RetimeWrapper_185_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54264.4]
  assign RetimeWrapper_185_io_in = _T_4285 & io_rPort_9_en_0; // @[package.scala 94:16:@54263.4]
  assign RetimeWrapper_186_clock = clock; // @[:@54269.4]
  assign RetimeWrapper_186_reset = reset; // @[:@54270.4]
  assign RetimeWrapper_186_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54272.4]
  assign RetimeWrapper_186_io_in = _T_4589 & io_rPort_9_en_0; // @[package.scala 94:16:@54271.4]
  assign RetimeWrapper_187_clock = clock; // @[:@54277.4]
  assign RetimeWrapper_187_reset = reset; // @[:@54278.4]
  assign RetimeWrapper_187_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54280.4]
  assign RetimeWrapper_187_io_in = _T_4893 & io_rPort_9_en_0; // @[package.scala 94:16:@54279.4]
  assign RetimeWrapper_188_clock = clock; // @[:@54285.4]
  assign RetimeWrapper_188_reset = reset; // @[:@54286.4]
  assign RetimeWrapper_188_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54288.4]
  assign RetimeWrapper_188_io_in = _T_5197 & io_rPort_9_en_0; // @[package.scala 94:16:@54287.4]
  assign RetimeWrapper_189_clock = clock; // @[:@54293.4]
  assign RetimeWrapper_189_reset = reset; // @[:@54294.4]
  assign RetimeWrapper_189_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54296.4]
  assign RetimeWrapper_189_io_in = _T_5501 & io_rPort_9_en_0; // @[package.scala 94:16:@54295.4]
  assign RetimeWrapper_190_clock = clock; // @[:@54301.4]
  assign RetimeWrapper_190_reset = reset; // @[:@54302.4]
  assign RetimeWrapper_190_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54304.4]
  assign RetimeWrapper_190_io_in = _T_5805 & io_rPort_9_en_0; // @[package.scala 94:16:@54303.4]
  assign RetimeWrapper_191_clock = clock; // @[:@54309.4]
  assign RetimeWrapper_191_reset = reset; // @[:@54310.4]
  assign RetimeWrapper_191_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54312.4]
  assign RetimeWrapper_191_io_in = _T_6109 & io_rPort_9_en_0; // @[package.scala 94:16:@54311.4]
  assign RetimeWrapper_192_clock = clock; // @[:@54317.4]
  assign RetimeWrapper_192_reset = reset; // @[:@54318.4]
  assign RetimeWrapper_192_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54320.4]
  assign RetimeWrapper_192_io_in = _T_6413 & io_rPort_9_en_0; // @[package.scala 94:16:@54319.4]
  assign RetimeWrapper_193_clock = clock; // @[:@54325.4]
  assign RetimeWrapper_193_reset = reset; // @[:@54326.4]
  assign RetimeWrapper_193_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54328.4]
  assign RetimeWrapper_193_io_in = _T_6717 & io_rPort_9_en_0; // @[package.scala 94:16:@54327.4]
  assign RetimeWrapper_194_clock = clock; // @[:@54333.4]
  assign RetimeWrapper_194_reset = reset; // @[:@54334.4]
  assign RetimeWrapper_194_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54336.4]
  assign RetimeWrapper_194_io_in = _T_7021 & io_rPort_9_en_0; // @[package.scala 94:16:@54335.4]
  assign RetimeWrapper_195_clock = clock; // @[:@54341.4]
  assign RetimeWrapper_195_reset = reset; // @[:@54342.4]
  assign RetimeWrapper_195_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54344.4]
  assign RetimeWrapper_195_io_in = _T_7325 & io_rPort_9_en_0; // @[package.scala 94:16:@54343.4]
  assign RetimeWrapper_196_clock = clock; // @[:@54349.4]
  assign RetimeWrapper_196_reset = reset; // @[:@54350.4]
  assign RetimeWrapper_196_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54352.4]
  assign RetimeWrapper_196_io_in = _T_7629 & io_rPort_9_en_0; // @[package.scala 94:16:@54351.4]
  assign RetimeWrapper_197_clock = clock; // @[:@54357.4]
  assign RetimeWrapper_197_reset = reset; // @[:@54358.4]
  assign RetimeWrapper_197_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54360.4]
  assign RetimeWrapper_197_io_in = _T_7933 & io_rPort_9_en_0; // @[package.scala 94:16:@54359.4]
  assign RetimeWrapper_198_clock = clock; // @[:@54365.4]
  assign RetimeWrapper_198_reset = reset; // @[:@54366.4]
  assign RetimeWrapper_198_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54368.4]
  assign RetimeWrapper_198_io_in = _T_8237 & io_rPort_9_en_0; // @[package.scala 94:16:@54367.4]
  assign RetimeWrapper_199_clock = clock; // @[:@54373.4]
  assign RetimeWrapper_199_reset = reset; // @[:@54374.4]
  assign RetimeWrapper_199_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@54376.4]
  assign RetimeWrapper_199_io_in = _T_8541 & io_rPort_9_en_0; // @[package.scala 94:16:@54375.4]
  assign RetimeWrapper_200_clock = clock; // @[:@54461.4]
  assign RetimeWrapper_200_reset = reset; // @[:@54462.4]
  assign RetimeWrapper_200_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54464.4]
  assign RetimeWrapper_200_io_in = _T_2771 & io_rPort_10_en_0; // @[package.scala 94:16:@54463.4]
  assign RetimeWrapper_201_clock = clock; // @[:@54469.4]
  assign RetimeWrapper_201_reset = reset; // @[:@54470.4]
  assign RetimeWrapper_201_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54472.4]
  assign RetimeWrapper_201_io_in = _T_3075 & io_rPort_10_en_0; // @[package.scala 94:16:@54471.4]
  assign RetimeWrapper_202_clock = clock; // @[:@54477.4]
  assign RetimeWrapper_202_reset = reset; // @[:@54478.4]
  assign RetimeWrapper_202_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54480.4]
  assign RetimeWrapper_202_io_in = _T_3379 & io_rPort_10_en_0; // @[package.scala 94:16:@54479.4]
  assign RetimeWrapper_203_clock = clock; // @[:@54485.4]
  assign RetimeWrapper_203_reset = reset; // @[:@54486.4]
  assign RetimeWrapper_203_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54488.4]
  assign RetimeWrapper_203_io_in = _T_3683 & io_rPort_10_en_0; // @[package.scala 94:16:@54487.4]
  assign RetimeWrapper_204_clock = clock; // @[:@54493.4]
  assign RetimeWrapper_204_reset = reset; // @[:@54494.4]
  assign RetimeWrapper_204_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54496.4]
  assign RetimeWrapper_204_io_in = _T_3987 & io_rPort_10_en_0; // @[package.scala 94:16:@54495.4]
  assign RetimeWrapper_205_clock = clock; // @[:@54501.4]
  assign RetimeWrapper_205_reset = reset; // @[:@54502.4]
  assign RetimeWrapper_205_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54504.4]
  assign RetimeWrapper_205_io_in = _T_4291 & io_rPort_10_en_0; // @[package.scala 94:16:@54503.4]
  assign RetimeWrapper_206_clock = clock; // @[:@54509.4]
  assign RetimeWrapper_206_reset = reset; // @[:@54510.4]
  assign RetimeWrapper_206_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54512.4]
  assign RetimeWrapper_206_io_in = _T_4595 & io_rPort_10_en_0; // @[package.scala 94:16:@54511.4]
  assign RetimeWrapper_207_clock = clock; // @[:@54517.4]
  assign RetimeWrapper_207_reset = reset; // @[:@54518.4]
  assign RetimeWrapper_207_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54520.4]
  assign RetimeWrapper_207_io_in = _T_4899 & io_rPort_10_en_0; // @[package.scala 94:16:@54519.4]
  assign RetimeWrapper_208_clock = clock; // @[:@54525.4]
  assign RetimeWrapper_208_reset = reset; // @[:@54526.4]
  assign RetimeWrapper_208_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54528.4]
  assign RetimeWrapper_208_io_in = _T_5203 & io_rPort_10_en_0; // @[package.scala 94:16:@54527.4]
  assign RetimeWrapper_209_clock = clock; // @[:@54533.4]
  assign RetimeWrapper_209_reset = reset; // @[:@54534.4]
  assign RetimeWrapper_209_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54536.4]
  assign RetimeWrapper_209_io_in = _T_5507 & io_rPort_10_en_0; // @[package.scala 94:16:@54535.4]
  assign RetimeWrapper_210_clock = clock; // @[:@54541.4]
  assign RetimeWrapper_210_reset = reset; // @[:@54542.4]
  assign RetimeWrapper_210_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54544.4]
  assign RetimeWrapper_210_io_in = _T_5811 & io_rPort_10_en_0; // @[package.scala 94:16:@54543.4]
  assign RetimeWrapper_211_clock = clock; // @[:@54549.4]
  assign RetimeWrapper_211_reset = reset; // @[:@54550.4]
  assign RetimeWrapper_211_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54552.4]
  assign RetimeWrapper_211_io_in = _T_6115 & io_rPort_10_en_0; // @[package.scala 94:16:@54551.4]
  assign RetimeWrapper_212_clock = clock; // @[:@54557.4]
  assign RetimeWrapper_212_reset = reset; // @[:@54558.4]
  assign RetimeWrapper_212_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54560.4]
  assign RetimeWrapper_212_io_in = _T_6419 & io_rPort_10_en_0; // @[package.scala 94:16:@54559.4]
  assign RetimeWrapper_213_clock = clock; // @[:@54565.4]
  assign RetimeWrapper_213_reset = reset; // @[:@54566.4]
  assign RetimeWrapper_213_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54568.4]
  assign RetimeWrapper_213_io_in = _T_6723 & io_rPort_10_en_0; // @[package.scala 94:16:@54567.4]
  assign RetimeWrapper_214_clock = clock; // @[:@54573.4]
  assign RetimeWrapper_214_reset = reset; // @[:@54574.4]
  assign RetimeWrapper_214_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54576.4]
  assign RetimeWrapper_214_io_in = _T_7027 & io_rPort_10_en_0; // @[package.scala 94:16:@54575.4]
  assign RetimeWrapper_215_clock = clock; // @[:@54581.4]
  assign RetimeWrapper_215_reset = reset; // @[:@54582.4]
  assign RetimeWrapper_215_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54584.4]
  assign RetimeWrapper_215_io_in = _T_7331 & io_rPort_10_en_0; // @[package.scala 94:16:@54583.4]
  assign RetimeWrapper_216_clock = clock; // @[:@54589.4]
  assign RetimeWrapper_216_reset = reset; // @[:@54590.4]
  assign RetimeWrapper_216_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54592.4]
  assign RetimeWrapper_216_io_in = _T_7635 & io_rPort_10_en_0; // @[package.scala 94:16:@54591.4]
  assign RetimeWrapper_217_clock = clock; // @[:@54597.4]
  assign RetimeWrapper_217_reset = reset; // @[:@54598.4]
  assign RetimeWrapper_217_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54600.4]
  assign RetimeWrapper_217_io_in = _T_7939 & io_rPort_10_en_0; // @[package.scala 94:16:@54599.4]
  assign RetimeWrapper_218_clock = clock; // @[:@54605.4]
  assign RetimeWrapper_218_reset = reset; // @[:@54606.4]
  assign RetimeWrapper_218_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54608.4]
  assign RetimeWrapper_218_io_in = _T_8243 & io_rPort_10_en_0; // @[package.scala 94:16:@54607.4]
  assign RetimeWrapper_219_clock = clock; // @[:@54613.4]
  assign RetimeWrapper_219_reset = reset; // @[:@54614.4]
  assign RetimeWrapper_219_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@54616.4]
  assign RetimeWrapper_219_io_in = _T_8547 & io_rPort_10_en_0; // @[package.scala 94:16:@54615.4]
  assign RetimeWrapper_220_clock = clock; // @[:@54701.4]
  assign RetimeWrapper_220_reset = reset; // @[:@54702.4]
  assign RetimeWrapper_220_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54704.4]
  assign RetimeWrapper_220_io_in = _T_2911 & io_rPort_11_en_0; // @[package.scala 94:16:@54703.4]
  assign RetimeWrapper_221_clock = clock; // @[:@54709.4]
  assign RetimeWrapper_221_reset = reset; // @[:@54710.4]
  assign RetimeWrapper_221_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54712.4]
  assign RetimeWrapper_221_io_in = _T_3215 & io_rPort_11_en_0; // @[package.scala 94:16:@54711.4]
  assign RetimeWrapper_222_clock = clock; // @[:@54717.4]
  assign RetimeWrapper_222_reset = reset; // @[:@54718.4]
  assign RetimeWrapper_222_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54720.4]
  assign RetimeWrapper_222_io_in = _T_3519 & io_rPort_11_en_0; // @[package.scala 94:16:@54719.4]
  assign RetimeWrapper_223_clock = clock; // @[:@54725.4]
  assign RetimeWrapper_223_reset = reset; // @[:@54726.4]
  assign RetimeWrapper_223_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54728.4]
  assign RetimeWrapper_223_io_in = _T_3823 & io_rPort_11_en_0; // @[package.scala 94:16:@54727.4]
  assign RetimeWrapper_224_clock = clock; // @[:@54733.4]
  assign RetimeWrapper_224_reset = reset; // @[:@54734.4]
  assign RetimeWrapper_224_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54736.4]
  assign RetimeWrapper_224_io_in = _T_4127 & io_rPort_11_en_0; // @[package.scala 94:16:@54735.4]
  assign RetimeWrapper_225_clock = clock; // @[:@54741.4]
  assign RetimeWrapper_225_reset = reset; // @[:@54742.4]
  assign RetimeWrapper_225_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54744.4]
  assign RetimeWrapper_225_io_in = _T_4431 & io_rPort_11_en_0; // @[package.scala 94:16:@54743.4]
  assign RetimeWrapper_226_clock = clock; // @[:@54749.4]
  assign RetimeWrapper_226_reset = reset; // @[:@54750.4]
  assign RetimeWrapper_226_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54752.4]
  assign RetimeWrapper_226_io_in = _T_4735 & io_rPort_11_en_0; // @[package.scala 94:16:@54751.4]
  assign RetimeWrapper_227_clock = clock; // @[:@54757.4]
  assign RetimeWrapper_227_reset = reset; // @[:@54758.4]
  assign RetimeWrapper_227_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54760.4]
  assign RetimeWrapper_227_io_in = _T_5039 & io_rPort_11_en_0; // @[package.scala 94:16:@54759.4]
  assign RetimeWrapper_228_clock = clock; // @[:@54765.4]
  assign RetimeWrapper_228_reset = reset; // @[:@54766.4]
  assign RetimeWrapper_228_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54768.4]
  assign RetimeWrapper_228_io_in = _T_5343 & io_rPort_11_en_0; // @[package.scala 94:16:@54767.4]
  assign RetimeWrapper_229_clock = clock; // @[:@54773.4]
  assign RetimeWrapper_229_reset = reset; // @[:@54774.4]
  assign RetimeWrapper_229_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54776.4]
  assign RetimeWrapper_229_io_in = _T_5647 & io_rPort_11_en_0; // @[package.scala 94:16:@54775.4]
  assign RetimeWrapper_230_clock = clock; // @[:@54781.4]
  assign RetimeWrapper_230_reset = reset; // @[:@54782.4]
  assign RetimeWrapper_230_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54784.4]
  assign RetimeWrapper_230_io_in = _T_5951 & io_rPort_11_en_0; // @[package.scala 94:16:@54783.4]
  assign RetimeWrapper_231_clock = clock; // @[:@54789.4]
  assign RetimeWrapper_231_reset = reset; // @[:@54790.4]
  assign RetimeWrapper_231_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54792.4]
  assign RetimeWrapper_231_io_in = _T_6255 & io_rPort_11_en_0; // @[package.scala 94:16:@54791.4]
  assign RetimeWrapper_232_clock = clock; // @[:@54797.4]
  assign RetimeWrapper_232_reset = reset; // @[:@54798.4]
  assign RetimeWrapper_232_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54800.4]
  assign RetimeWrapper_232_io_in = _T_6559 & io_rPort_11_en_0; // @[package.scala 94:16:@54799.4]
  assign RetimeWrapper_233_clock = clock; // @[:@54805.4]
  assign RetimeWrapper_233_reset = reset; // @[:@54806.4]
  assign RetimeWrapper_233_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54808.4]
  assign RetimeWrapper_233_io_in = _T_6863 & io_rPort_11_en_0; // @[package.scala 94:16:@54807.4]
  assign RetimeWrapper_234_clock = clock; // @[:@54813.4]
  assign RetimeWrapper_234_reset = reset; // @[:@54814.4]
  assign RetimeWrapper_234_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54816.4]
  assign RetimeWrapper_234_io_in = _T_7167 & io_rPort_11_en_0; // @[package.scala 94:16:@54815.4]
  assign RetimeWrapper_235_clock = clock; // @[:@54821.4]
  assign RetimeWrapper_235_reset = reset; // @[:@54822.4]
  assign RetimeWrapper_235_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54824.4]
  assign RetimeWrapper_235_io_in = _T_7471 & io_rPort_11_en_0; // @[package.scala 94:16:@54823.4]
  assign RetimeWrapper_236_clock = clock; // @[:@54829.4]
  assign RetimeWrapper_236_reset = reset; // @[:@54830.4]
  assign RetimeWrapper_236_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54832.4]
  assign RetimeWrapper_236_io_in = _T_7775 & io_rPort_11_en_0; // @[package.scala 94:16:@54831.4]
  assign RetimeWrapper_237_clock = clock; // @[:@54837.4]
  assign RetimeWrapper_237_reset = reset; // @[:@54838.4]
  assign RetimeWrapper_237_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54840.4]
  assign RetimeWrapper_237_io_in = _T_8079 & io_rPort_11_en_0; // @[package.scala 94:16:@54839.4]
  assign RetimeWrapper_238_clock = clock; // @[:@54845.4]
  assign RetimeWrapper_238_reset = reset; // @[:@54846.4]
  assign RetimeWrapper_238_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54848.4]
  assign RetimeWrapper_238_io_in = _T_8383 & io_rPort_11_en_0; // @[package.scala 94:16:@54847.4]
  assign RetimeWrapper_239_clock = clock; // @[:@54853.4]
  assign RetimeWrapper_239_reset = reset; // @[:@54854.4]
  assign RetimeWrapper_239_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@54856.4]
  assign RetimeWrapper_239_io_in = _T_8687 & io_rPort_11_en_0; // @[package.scala 94:16:@54855.4]
  assign RetimeWrapper_240_clock = clock; // @[:@54941.4]
  assign RetimeWrapper_240_reset = reset; // @[:@54942.4]
  assign RetimeWrapper_240_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@54944.4]
  assign RetimeWrapper_240_io_in = _T_2917 & io_rPort_12_en_0; // @[package.scala 94:16:@54943.4]
  assign RetimeWrapper_241_clock = clock; // @[:@54949.4]
  assign RetimeWrapper_241_reset = reset; // @[:@54950.4]
  assign RetimeWrapper_241_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@54952.4]
  assign RetimeWrapper_241_io_in = _T_3221 & io_rPort_12_en_0; // @[package.scala 94:16:@54951.4]
  assign RetimeWrapper_242_clock = clock; // @[:@54957.4]
  assign RetimeWrapper_242_reset = reset; // @[:@54958.4]
  assign RetimeWrapper_242_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@54960.4]
  assign RetimeWrapper_242_io_in = _T_3525 & io_rPort_12_en_0; // @[package.scala 94:16:@54959.4]
  assign RetimeWrapper_243_clock = clock; // @[:@54965.4]
  assign RetimeWrapper_243_reset = reset; // @[:@54966.4]
  assign RetimeWrapper_243_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@54968.4]
  assign RetimeWrapper_243_io_in = _T_3829 & io_rPort_12_en_0; // @[package.scala 94:16:@54967.4]
  assign RetimeWrapper_244_clock = clock; // @[:@54973.4]
  assign RetimeWrapper_244_reset = reset; // @[:@54974.4]
  assign RetimeWrapper_244_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@54976.4]
  assign RetimeWrapper_244_io_in = _T_4133 & io_rPort_12_en_0; // @[package.scala 94:16:@54975.4]
  assign RetimeWrapper_245_clock = clock; // @[:@54981.4]
  assign RetimeWrapper_245_reset = reset; // @[:@54982.4]
  assign RetimeWrapper_245_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@54984.4]
  assign RetimeWrapper_245_io_in = _T_4437 & io_rPort_12_en_0; // @[package.scala 94:16:@54983.4]
  assign RetimeWrapper_246_clock = clock; // @[:@54989.4]
  assign RetimeWrapper_246_reset = reset; // @[:@54990.4]
  assign RetimeWrapper_246_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@54992.4]
  assign RetimeWrapper_246_io_in = _T_4741 & io_rPort_12_en_0; // @[package.scala 94:16:@54991.4]
  assign RetimeWrapper_247_clock = clock; // @[:@54997.4]
  assign RetimeWrapper_247_reset = reset; // @[:@54998.4]
  assign RetimeWrapper_247_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55000.4]
  assign RetimeWrapper_247_io_in = _T_5045 & io_rPort_12_en_0; // @[package.scala 94:16:@54999.4]
  assign RetimeWrapper_248_clock = clock; // @[:@55005.4]
  assign RetimeWrapper_248_reset = reset; // @[:@55006.4]
  assign RetimeWrapper_248_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55008.4]
  assign RetimeWrapper_248_io_in = _T_5349 & io_rPort_12_en_0; // @[package.scala 94:16:@55007.4]
  assign RetimeWrapper_249_clock = clock; // @[:@55013.4]
  assign RetimeWrapper_249_reset = reset; // @[:@55014.4]
  assign RetimeWrapper_249_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55016.4]
  assign RetimeWrapper_249_io_in = _T_5653 & io_rPort_12_en_0; // @[package.scala 94:16:@55015.4]
  assign RetimeWrapper_250_clock = clock; // @[:@55021.4]
  assign RetimeWrapper_250_reset = reset; // @[:@55022.4]
  assign RetimeWrapper_250_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55024.4]
  assign RetimeWrapper_250_io_in = _T_5957 & io_rPort_12_en_0; // @[package.scala 94:16:@55023.4]
  assign RetimeWrapper_251_clock = clock; // @[:@55029.4]
  assign RetimeWrapper_251_reset = reset; // @[:@55030.4]
  assign RetimeWrapper_251_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55032.4]
  assign RetimeWrapper_251_io_in = _T_6261 & io_rPort_12_en_0; // @[package.scala 94:16:@55031.4]
  assign RetimeWrapper_252_clock = clock; // @[:@55037.4]
  assign RetimeWrapper_252_reset = reset; // @[:@55038.4]
  assign RetimeWrapper_252_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55040.4]
  assign RetimeWrapper_252_io_in = _T_6565 & io_rPort_12_en_0; // @[package.scala 94:16:@55039.4]
  assign RetimeWrapper_253_clock = clock; // @[:@55045.4]
  assign RetimeWrapper_253_reset = reset; // @[:@55046.4]
  assign RetimeWrapper_253_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55048.4]
  assign RetimeWrapper_253_io_in = _T_6869 & io_rPort_12_en_0; // @[package.scala 94:16:@55047.4]
  assign RetimeWrapper_254_clock = clock; // @[:@55053.4]
  assign RetimeWrapper_254_reset = reset; // @[:@55054.4]
  assign RetimeWrapper_254_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55056.4]
  assign RetimeWrapper_254_io_in = _T_7173 & io_rPort_12_en_0; // @[package.scala 94:16:@55055.4]
  assign RetimeWrapper_255_clock = clock; // @[:@55061.4]
  assign RetimeWrapper_255_reset = reset; // @[:@55062.4]
  assign RetimeWrapper_255_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55064.4]
  assign RetimeWrapper_255_io_in = _T_7477 & io_rPort_12_en_0; // @[package.scala 94:16:@55063.4]
  assign RetimeWrapper_256_clock = clock; // @[:@55069.4]
  assign RetimeWrapper_256_reset = reset; // @[:@55070.4]
  assign RetimeWrapper_256_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55072.4]
  assign RetimeWrapper_256_io_in = _T_7781 & io_rPort_12_en_0; // @[package.scala 94:16:@55071.4]
  assign RetimeWrapper_257_clock = clock; // @[:@55077.4]
  assign RetimeWrapper_257_reset = reset; // @[:@55078.4]
  assign RetimeWrapper_257_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55080.4]
  assign RetimeWrapper_257_io_in = _T_8085 & io_rPort_12_en_0; // @[package.scala 94:16:@55079.4]
  assign RetimeWrapper_258_clock = clock; // @[:@55085.4]
  assign RetimeWrapper_258_reset = reset; // @[:@55086.4]
  assign RetimeWrapper_258_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55088.4]
  assign RetimeWrapper_258_io_in = _T_8389 & io_rPort_12_en_0; // @[package.scala 94:16:@55087.4]
  assign RetimeWrapper_259_clock = clock; // @[:@55093.4]
  assign RetimeWrapper_259_reset = reset; // @[:@55094.4]
  assign RetimeWrapper_259_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@55096.4]
  assign RetimeWrapper_259_io_in = _T_8693 & io_rPort_12_en_0; // @[package.scala 94:16:@55095.4]
  assign RetimeWrapper_260_clock = clock; // @[:@55181.4]
  assign RetimeWrapper_260_reset = reset; // @[:@55182.4]
  assign RetimeWrapper_260_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55184.4]
  assign RetimeWrapper_260_io_in = _T_2777 & io_rPort_13_en_0; // @[package.scala 94:16:@55183.4]
  assign RetimeWrapper_261_clock = clock; // @[:@55189.4]
  assign RetimeWrapper_261_reset = reset; // @[:@55190.4]
  assign RetimeWrapper_261_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55192.4]
  assign RetimeWrapper_261_io_in = _T_3081 & io_rPort_13_en_0; // @[package.scala 94:16:@55191.4]
  assign RetimeWrapper_262_clock = clock; // @[:@55197.4]
  assign RetimeWrapper_262_reset = reset; // @[:@55198.4]
  assign RetimeWrapper_262_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55200.4]
  assign RetimeWrapper_262_io_in = _T_3385 & io_rPort_13_en_0; // @[package.scala 94:16:@55199.4]
  assign RetimeWrapper_263_clock = clock; // @[:@55205.4]
  assign RetimeWrapper_263_reset = reset; // @[:@55206.4]
  assign RetimeWrapper_263_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55208.4]
  assign RetimeWrapper_263_io_in = _T_3689 & io_rPort_13_en_0; // @[package.scala 94:16:@55207.4]
  assign RetimeWrapper_264_clock = clock; // @[:@55213.4]
  assign RetimeWrapper_264_reset = reset; // @[:@55214.4]
  assign RetimeWrapper_264_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55216.4]
  assign RetimeWrapper_264_io_in = _T_3993 & io_rPort_13_en_0; // @[package.scala 94:16:@55215.4]
  assign RetimeWrapper_265_clock = clock; // @[:@55221.4]
  assign RetimeWrapper_265_reset = reset; // @[:@55222.4]
  assign RetimeWrapper_265_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55224.4]
  assign RetimeWrapper_265_io_in = _T_4297 & io_rPort_13_en_0; // @[package.scala 94:16:@55223.4]
  assign RetimeWrapper_266_clock = clock; // @[:@55229.4]
  assign RetimeWrapper_266_reset = reset; // @[:@55230.4]
  assign RetimeWrapper_266_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55232.4]
  assign RetimeWrapper_266_io_in = _T_4601 & io_rPort_13_en_0; // @[package.scala 94:16:@55231.4]
  assign RetimeWrapper_267_clock = clock; // @[:@55237.4]
  assign RetimeWrapper_267_reset = reset; // @[:@55238.4]
  assign RetimeWrapper_267_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55240.4]
  assign RetimeWrapper_267_io_in = _T_4905 & io_rPort_13_en_0; // @[package.scala 94:16:@55239.4]
  assign RetimeWrapper_268_clock = clock; // @[:@55245.4]
  assign RetimeWrapper_268_reset = reset; // @[:@55246.4]
  assign RetimeWrapper_268_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55248.4]
  assign RetimeWrapper_268_io_in = _T_5209 & io_rPort_13_en_0; // @[package.scala 94:16:@55247.4]
  assign RetimeWrapper_269_clock = clock; // @[:@55253.4]
  assign RetimeWrapper_269_reset = reset; // @[:@55254.4]
  assign RetimeWrapper_269_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55256.4]
  assign RetimeWrapper_269_io_in = _T_5513 & io_rPort_13_en_0; // @[package.scala 94:16:@55255.4]
  assign RetimeWrapper_270_clock = clock; // @[:@55261.4]
  assign RetimeWrapper_270_reset = reset; // @[:@55262.4]
  assign RetimeWrapper_270_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55264.4]
  assign RetimeWrapper_270_io_in = _T_5817 & io_rPort_13_en_0; // @[package.scala 94:16:@55263.4]
  assign RetimeWrapper_271_clock = clock; // @[:@55269.4]
  assign RetimeWrapper_271_reset = reset; // @[:@55270.4]
  assign RetimeWrapper_271_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55272.4]
  assign RetimeWrapper_271_io_in = _T_6121 & io_rPort_13_en_0; // @[package.scala 94:16:@55271.4]
  assign RetimeWrapper_272_clock = clock; // @[:@55277.4]
  assign RetimeWrapper_272_reset = reset; // @[:@55278.4]
  assign RetimeWrapper_272_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55280.4]
  assign RetimeWrapper_272_io_in = _T_6425 & io_rPort_13_en_0; // @[package.scala 94:16:@55279.4]
  assign RetimeWrapper_273_clock = clock; // @[:@55285.4]
  assign RetimeWrapper_273_reset = reset; // @[:@55286.4]
  assign RetimeWrapper_273_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55288.4]
  assign RetimeWrapper_273_io_in = _T_6729 & io_rPort_13_en_0; // @[package.scala 94:16:@55287.4]
  assign RetimeWrapper_274_clock = clock; // @[:@55293.4]
  assign RetimeWrapper_274_reset = reset; // @[:@55294.4]
  assign RetimeWrapper_274_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55296.4]
  assign RetimeWrapper_274_io_in = _T_7033 & io_rPort_13_en_0; // @[package.scala 94:16:@55295.4]
  assign RetimeWrapper_275_clock = clock; // @[:@55301.4]
  assign RetimeWrapper_275_reset = reset; // @[:@55302.4]
  assign RetimeWrapper_275_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55304.4]
  assign RetimeWrapper_275_io_in = _T_7337 & io_rPort_13_en_0; // @[package.scala 94:16:@55303.4]
  assign RetimeWrapper_276_clock = clock; // @[:@55309.4]
  assign RetimeWrapper_276_reset = reset; // @[:@55310.4]
  assign RetimeWrapper_276_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55312.4]
  assign RetimeWrapper_276_io_in = _T_7641 & io_rPort_13_en_0; // @[package.scala 94:16:@55311.4]
  assign RetimeWrapper_277_clock = clock; // @[:@55317.4]
  assign RetimeWrapper_277_reset = reset; // @[:@55318.4]
  assign RetimeWrapper_277_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55320.4]
  assign RetimeWrapper_277_io_in = _T_7945 & io_rPort_13_en_0; // @[package.scala 94:16:@55319.4]
  assign RetimeWrapper_278_clock = clock; // @[:@55325.4]
  assign RetimeWrapper_278_reset = reset; // @[:@55326.4]
  assign RetimeWrapper_278_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55328.4]
  assign RetimeWrapper_278_io_in = _T_8249 & io_rPort_13_en_0; // @[package.scala 94:16:@55327.4]
  assign RetimeWrapper_279_clock = clock; // @[:@55333.4]
  assign RetimeWrapper_279_reset = reset; // @[:@55334.4]
  assign RetimeWrapper_279_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@55336.4]
  assign RetimeWrapper_279_io_in = _T_8553 & io_rPort_13_en_0; // @[package.scala 94:16:@55335.4]
  assign RetimeWrapper_280_clock = clock; // @[:@55421.4]
  assign RetimeWrapper_280_reset = reset; // @[:@55422.4]
  assign RetimeWrapper_280_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55424.4]
  assign RetimeWrapper_280_io_in = _T_2923 & io_rPort_14_en_0; // @[package.scala 94:16:@55423.4]
  assign RetimeWrapper_281_clock = clock; // @[:@55429.4]
  assign RetimeWrapper_281_reset = reset; // @[:@55430.4]
  assign RetimeWrapper_281_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55432.4]
  assign RetimeWrapper_281_io_in = _T_3227 & io_rPort_14_en_0; // @[package.scala 94:16:@55431.4]
  assign RetimeWrapper_282_clock = clock; // @[:@55437.4]
  assign RetimeWrapper_282_reset = reset; // @[:@55438.4]
  assign RetimeWrapper_282_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55440.4]
  assign RetimeWrapper_282_io_in = _T_3531 & io_rPort_14_en_0; // @[package.scala 94:16:@55439.4]
  assign RetimeWrapper_283_clock = clock; // @[:@55445.4]
  assign RetimeWrapper_283_reset = reset; // @[:@55446.4]
  assign RetimeWrapper_283_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55448.4]
  assign RetimeWrapper_283_io_in = _T_3835 & io_rPort_14_en_0; // @[package.scala 94:16:@55447.4]
  assign RetimeWrapper_284_clock = clock; // @[:@55453.4]
  assign RetimeWrapper_284_reset = reset; // @[:@55454.4]
  assign RetimeWrapper_284_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55456.4]
  assign RetimeWrapper_284_io_in = _T_4139 & io_rPort_14_en_0; // @[package.scala 94:16:@55455.4]
  assign RetimeWrapper_285_clock = clock; // @[:@55461.4]
  assign RetimeWrapper_285_reset = reset; // @[:@55462.4]
  assign RetimeWrapper_285_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55464.4]
  assign RetimeWrapper_285_io_in = _T_4443 & io_rPort_14_en_0; // @[package.scala 94:16:@55463.4]
  assign RetimeWrapper_286_clock = clock; // @[:@55469.4]
  assign RetimeWrapper_286_reset = reset; // @[:@55470.4]
  assign RetimeWrapper_286_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55472.4]
  assign RetimeWrapper_286_io_in = _T_4747 & io_rPort_14_en_0; // @[package.scala 94:16:@55471.4]
  assign RetimeWrapper_287_clock = clock; // @[:@55477.4]
  assign RetimeWrapper_287_reset = reset; // @[:@55478.4]
  assign RetimeWrapper_287_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55480.4]
  assign RetimeWrapper_287_io_in = _T_5051 & io_rPort_14_en_0; // @[package.scala 94:16:@55479.4]
  assign RetimeWrapper_288_clock = clock; // @[:@55485.4]
  assign RetimeWrapper_288_reset = reset; // @[:@55486.4]
  assign RetimeWrapper_288_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55488.4]
  assign RetimeWrapper_288_io_in = _T_5355 & io_rPort_14_en_0; // @[package.scala 94:16:@55487.4]
  assign RetimeWrapper_289_clock = clock; // @[:@55493.4]
  assign RetimeWrapper_289_reset = reset; // @[:@55494.4]
  assign RetimeWrapper_289_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55496.4]
  assign RetimeWrapper_289_io_in = _T_5659 & io_rPort_14_en_0; // @[package.scala 94:16:@55495.4]
  assign RetimeWrapper_290_clock = clock; // @[:@55501.4]
  assign RetimeWrapper_290_reset = reset; // @[:@55502.4]
  assign RetimeWrapper_290_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55504.4]
  assign RetimeWrapper_290_io_in = _T_5963 & io_rPort_14_en_0; // @[package.scala 94:16:@55503.4]
  assign RetimeWrapper_291_clock = clock; // @[:@55509.4]
  assign RetimeWrapper_291_reset = reset; // @[:@55510.4]
  assign RetimeWrapper_291_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55512.4]
  assign RetimeWrapper_291_io_in = _T_6267 & io_rPort_14_en_0; // @[package.scala 94:16:@55511.4]
  assign RetimeWrapper_292_clock = clock; // @[:@55517.4]
  assign RetimeWrapper_292_reset = reset; // @[:@55518.4]
  assign RetimeWrapper_292_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55520.4]
  assign RetimeWrapper_292_io_in = _T_6571 & io_rPort_14_en_0; // @[package.scala 94:16:@55519.4]
  assign RetimeWrapper_293_clock = clock; // @[:@55525.4]
  assign RetimeWrapper_293_reset = reset; // @[:@55526.4]
  assign RetimeWrapper_293_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55528.4]
  assign RetimeWrapper_293_io_in = _T_6875 & io_rPort_14_en_0; // @[package.scala 94:16:@55527.4]
  assign RetimeWrapper_294_clock = clock; // @[:@55533.4]
  assign RetimeWrapper_294_reset = reset; // @[:@55534.4]
  assign RetimeWrapper_294_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55536.4]
  assign RetimeWrapper_294_io_in = _T_7179 & io_rPort_14_en_0; // @[package.scala 94:16:@55535.4]
  assign RetimeWrapper_295_clock = clock; // @[:@55541.4]
  assign RetimeWrapper_295_reset = reset; // @[:@55542.4]
  assign RetimeWrapper_295_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55544.4]
  assign RetimeWrapper_295_io_in = _T_7483 & io_rPort_14_en_0; // @[package.scala 94:16:@55543.4]
  assign RetimeWrapper_296_clock = clock; // @[:@55549.4]
  assign RetimeWrapper_296_reset = reset; // @[:@55550.4]
  assign RetimeWrapper_296_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55552.4]
  assign RetimeWrapper_296_io_in = _T_7787 & io_rPort_14_en_0; // @[package.scala 94:16:@55551.4]
  assign RetimeWrapper_297_clock = clock; // @[:@55557.4]
  assign RetimeWrapper_297_reset = reset; // @[:@55558.4]
  assign RetimeWrapper_297_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55560.4]
  assign RetimeWrapper_297_io_in = _T_8091 & io_rPort_14_en_0; // @[package.scala 94:16:@55559.4]
  assign RetimeWrapper_298_clock = clock; // @[:@55565.4]
  assign RetimeWrapper_298_reset = reset; // @[:@55566.4]
  assign RetimeWrapper_298_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55568.4]
  assign RetimeWrapper_298_io_in = _T_8395 & io_rPort_14_en_0; // @[package.scala 94:16:@55567.4]
  assign RetimeWrapper_299_clock = clock; // @[:@55573.4]
  assign RetimeWrapper_299_reset = reset; // @[:@55574.4]
  assign RetimeWrapper_299_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@55576.4]
  assign RetimeWrapper_299_io_in = _T_8699 & io_rPort_14_en_0; // @[package.scala 94:16:@55575.4]
  assign RetimeWrapper_300_clock = clock; // @[:@55661.4]
  assign RetimeWrapper_300_reset = reset; // @[:@55662.4]
  assign RetimeWrapper_300_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55664.4]
  assign RetimeWrapper_300_io_in = _T_2783 & io_rPort_15_en_0; // @[package.scala 94:16:@55663.4]
  assign RetimeWrapper_301_clock = clock; // @[:@55669.4]
  assign RetimeWrapper_301_reset = reset; // @[:@55670.4]
  assign RetimeWrapper_301_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55672.4]
  assign RetimeWrapper_301_io_in = _T_3087 & io_rPort_15_en_0; // @[package.scala 94:16:@55671.4]
  assign RetimeWrapper_302_clock = clock; // @[:@55677.4]
  assign RetimeWrapper_302_reset = reset; // @[:@55678.4]
  assign RetimeWrapper_302_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55680.4]
  assign RetimeWrapper_302_io_in = _T_3391 & io_rPort_15_en_0; // @[package.scala 94:16:@55679.4]
  assign RetimeWrapper_303_clock = clock; // @[:@55685.4]
  assign RetimeWrapper_303_reset = reset; // @[:@55686.4]
  assign RetimeWrapper_303_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55688.4]
  assign RetimeWrapper_303_io_in = _T_3695 & io_rPort_15_en_0; // @[package.scala 94:16:@55687.4]
  assign RetimeWrapper_304_clock = clock; // @[:@55693.4]
  assign RetimeWrapper_304_reset = reset; // @[:@55694.4]
  assign RetimeWrapper_304_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55696.4]
  assign RetimeWrapper_304_io_in = _T_3999 & io_rPort_15_en_0; // @[package.scala 94:16:@55695.4]
  assign RetimeWrapper_305_clock = clock; // @[:@55701.4]
  assign RetimeWrapper_305_reset = reset; // @[:@55702.4]
  assign RetimeWrapper_305_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55704.4]
  assign RetimeWrapper_305_io_in = _T_4303 & io_rPort_15_en_0; // @[package.scala 94:16:@55703.4]
  assign RetimeWrapper_306_clock = clock; // @[:@55709.4]
  assign RetimeWrapper_306_reset = reset; // @[:@55710.4]
  assign RetimeWrapper_306_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55712.4]
  assign RetimeWrapper_306_io_in = _T_4607 & io_rPort_15_en_0; // @[package.scala 94:16:@55711.4]
  assign RetimeWrapper_307_clock = clock; // @[:@55717.4]
  assign RetimeWrapper_307_reset = reset; // @[:@55718.4]
  assign RetimeWrapper_307_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55720.4]
  assign RetimeWrapper_307_io_in = _T_4911 & io_rPort_15_en_0; // @[package.scala 94:16:@55719.4]
  assign RetimeWrapper_308_clock = clock; // @[:@55725.4]
  assign RetimeWrapper_308_reset = reset; // @[:@55726.4]
  assign RetimeWrapper_308_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55728.4]
  assign RetimeWrapper_308_io_in = _T_5215 & io_rPort_15_en_0; // @[package.scala 94:16:@55727.4]
  assign RetimeWrapper_309_clock = clock; // @[:@55733.4]
  assign RetimeWrapper_309_reset = reset; // @[:@55734.4]
  assign RetimeWrapper_309_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55736.4]
  assign RetimeWrapper_309_io_in = _T_5519 & io_rPort_15_en_0; // @[package.scala 94:16:@55735.4]
  assign RetimeWrapper_310_clock = clock; // @[:@55741.4]
  assign RetimeWrapper_310_reset = reset; // @[:@55742.4]
  assign RetimeWrapper_310_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55744.4]
  assign RetimeWrapper_310_io_in = _T_5823 & io_rPort_15_en_0; // @[package.scala 94:16:@55743.4]
  assign RetimeWrapper_311_clock = clock; // @[:@55749.4]
  assign RetimeWrapper_311_reset = reset; // @[:@55750.4]
  assign RetimeWrapper_311_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55752.4]
  assign RetimeWrapper_311_io_in = _T_6127 & io_rPort_15_en_0; // @[package.scala 94:16:@55751.4]
  assign RetimeWrapper_312_clock = clock; // @[:@55757.4]
  assign RetimeWrapper_312_reset = reset; // @[:@55758.4]
  assign RetimeWrapper_312_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55760.4]
  assign RetimeWrapper_312_io_in = _T_6431 & io_rPort_15_en_0; // @[package.scala 94:16:@55759.4]
  assign RetimeWrapper_313_clock = clock; // @[:@55765.4]
  assign RetimeWrapper_313_reset = reset; // @[:@55766.4]
  assign RetimeWrapper_313_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55768.4]
  assign RetimeWrapper_313_io_in = _T_6735 & io_rPort_15_en_0; // @[package.scala 94:16:@55767.4]
  assign RetimeWrapper_314_clock = clock; // @[:@55773.4]
  assign RetimeWrapper_314_reset = reset; // @[:@55774.4]
  assign RetimeWrapper_314_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55776.4]
  assign RetimeWrapper_314_io_in = _T_7039 & io_rPort_15_en_0; // @[package.scala 94:16:@55775.4]
  assign RetimeWrapper_315_clock = clock; // @[:@55781.4]
  assign RetimeWrapper_315_reset = reset; // @[:@55782.4]
  assign RetimeWrapper_315_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55784.4]
  assign RetimeWrapper_315_io_in = _T_7343 & io_rPort_15_en_0; // @[package.scala 94:16:@55783.4]
  assign RetimeWrapper_316_clock = clock; // @[:@55789.4]
  assign RetimeWrapper_316_reset = reset; // @[:@55790.4]
  assign RetimeWrapper_316_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55792.4]
  assign RetimeWrapper_316_io_in = _T_7647 & io_rPort_15_en_0; // @[package.scala 94:16:@55791.4]
  assign RetimeWrapper_317_clock = clock; // @[:@55797.4]
  assign RetimeWrapper_317_reset = reset; // @[:@55798.4]
  assign RetimeWrapper_317_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55800.4]
  assign RetimeWrapper_317_io_in = _T_7951 & io_rPort_15_en_0; // @[package.scala 94:16:@55799.4]
  assign RetimeWrapper_318_clock = clock; // @[:@55805.4]
  assign RetimeWrapper_318_reset = reset; // @[:@55806.4]
  assign RetimeWrapper_318_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55808.4]
  assign RetimeWrapper_318_io_in = _T_8255 & io_rPort_15_en_0; // @[package.scala 94:16:@55807.4]
  assign RetimeWrapper_319_clock = clock; // @[:@55813.4]
  assign RetimeWrapper_319_reset = reset; // @[:@55814.4]
  assign RetimeWrapper_319_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@55816.4]
  assign RetimeWrapper_319_io_in = _T_8559 & io_rPort_15_en_0; // @[package.scala 94:16:@55815.4]
  assign RetimeWrapper_320_clock = clock; // @[:@55901.4]
  assign RetimeWrapper_320_reset = reset; // @[:@55902.4]
  assign RetimeWrapper_320_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55904.4]
  assign RetimeWrapper_320_io_in = _T_2789 & io_rPort_16_en_0; // @[package.scala 94:16:@55903.4]
  assign RetimeWrapper_321_clock = clock; // @[:@55909.4]
  assign RetimeWrapper_321_reset = reset; // @[:@55910.4]
  assign RetimeWrapper_321_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55912.4]
  assign RetimeWrapper_321_io_in = _T_3093 & io_rPort_16_en_0; // @[package.scala 94:16:@55911.4]
  assign RetimeWrapper_322_clock = clock; // @[:@55917.4]
  assign RetimeWrapper_322_reset = reset; // @[:@55918.4]
  assign RetimeWrapper_322_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55920.4]
  assign RetimeWrapper_322_io_in = _T_3397 & io_rPort_16_en_0; // @[package.scala 94:16:@55919.4]
  assign RetimeWrapper_323_clock = clock; // @[:@55925.4]
  assign RetimeWrapper_323_reset = reset; // @[:@55926.4]
  assign RetimeWrapper_323_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55928.4]
  assign RetimeWrapper_323_io_in = _T_3701 & io_rPort_16_en_0; // @[package.scala 94:16:@55927.4]
  assign RetimeWrapper_324_clock = clock; // @[:@55933.4]
  assign RetimeWrapper_324_reset = reset; // @[:@55934.4]
  assign RetimeWrapper_324_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55936.4]
  assign RetimeWrapper_324_io_in = _T_4005 & io_rPort_16_en_0; // @[package.scala 94:16:@55935.4]
  assign RetimeWrapper_325_clock = clock; // @[:@55941.4]
  assign RetimeWrapper_325_reset = reset; // @[:@55942.4]
  assign RetimeWrapper_325_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55944.4]
  assign RetimeWrapper_325_io_in = _T_4309 & io_rPort_16_en_0; // @[package.scala 94:16:@55943.4]
  assign RetimeWrapper_326_clock = clock; // @[:@55949.4]
  assign RetimeWrapper_326_reset = reset; // @[:@55950.4]
  assign RetimeWrapper_326_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55952.4]
  assign RetimeWrapper_326_io_in = _T_4613 & io_rPort_16_en_0; // @[package.scala 94:16:@55951.4]
  assign RetimeWrapper_327_clock = clock; // @[:@55957.4]
  assign RetimeWrapper_327_reset = reset; // @[:@55958.4]
  assign RetimeWrapper_327_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55960.4]
  assign RetimeWrapper_327_io_in = _T_4917 & io_rPort_16_en_0; // @[package.scala 94:16:@55959.4]
  assign RetimeWrapper_328_clock = clock; // @[:@55965.4]
  assign RetimeWrapper_328_reset = reset; // @[:@55966.4]
  assign RetimeWrapper_328_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55968.4]
  assign RetimeWrapper_328_io_in = _T_5221 & io_rPort_16_en_0; // @[package.scala 94:16:@55967.4]
  assign RetimeWrapper_329_clock = clock; // @[:@55973.4]
  assign RetimeWrapper_329_reset = reset; // @[:@55974.4]
  assign RetimeWrapper_329_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55976.4]
  assign RetimeWrapper_329_io_in = _T_5525 & io_rPort_16_en_0; // @[package.scala 94:16:@55975.4]
  assign RetimeWrapper_330_clock = clock; // @[:@55981.4]
  assign RetimeWrapper_330_reset = reset; // @[:@55982.4]
  assign RetimeWrapper_330_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55984.4]
  assign RetimeWrapper_330_io_in = _T_5829 & io_rPort_16_en_0; // @[package.scala 94:16:@55983.4]
  assign RetimeWrapper_331_clock = clock; // @[:@55989.4]
  assign RetimeWrapper_331_reset = reset; // @[:@55990.4]
  assign RetimeWrapper_331_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@55992.4]
  assign RetimeWrapper_331_io_in = _T_6133 & io_rPort_16_en_0; // @[package.scala 94:16:@55991.4]
  assign RetimeWrapper_332_clock = clock; // @[:@55997.4]
  assign RetimeWrapper_332_reset = reset; // @[:@55998.4]
  assign RetimeWrapper_332_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56000.4]
  assign RetimeWrapper_332_io_in = _T_6437 & io_rPort_16_en_0; // @[package.scala 94:16:@55999.4]
  assign RetimeWrapper_333_clock = clock; // @[:@56005.4]
  assign RetimeWrapper_333_reset = reset; // @[:@56006.4]
  assign RetimeWrapper_333_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56008.4]
  assign RetimeWrapper_333_io_in = _T_6741 & io_rPort_16_en_0; // @[package.scala 94:16:@56007.4]
  assign RetimeWrapper_334_clock = clock; // @[:@56013.4]
  assign RetimeWrapper_334_reset = reset; // @[:@56014.4]
  assign RetimeWrapper_334_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56016.4]
  assign RetimeWrapper_334_io_in = _T_7045 & io_rPort_16_en_0; // @[package.scala 94:16:@56015.4]
  assign RetimeWrapper_335_clock = clock; // @[:@56021.4]
  assign RetimeWrapper_335_reset = reset; // @[:@56022.4]
  assign RetimeWrapper_335_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56024.4]
  assign RetimeWrapper_335_io_in = _T_7349 & io_rPort_16_en_0; // @[package.scala 94:16:@56023.4]
  assign RetimeWrapper_336_clock = clock; // @[:@56029.4]
  assign RetimeWrapper_336_reset = reset; // @[:@56030.4]
  assign RetimeWrapper_336_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56032.4]
  assign RetimeWrapper_336_io_in = _T_7653 & io_rPort_16_en_0; // @[package.scala 94:16:@56031.4]
  assign RetimeWrapper_337_clock = clock; // @[:@56037.4]
  assign RetimeWrapper_337_reset = reset; // @[:@56038.4]
  assign RetimeWrapper_337_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56040.4]
  assign RetimeWrapper_337_io_in = _T_7957 & io_rPort_16_en_0; // @[package.scala 94:16:@56039.4]
  assign RetimeWrapper_338_clock = clock; // @[:@56045.4]
  assign RetimeWrapper_338_reset = reset; // @[:@56046.4]
  assign RetimeWrapper_338_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56048.4]
  assign RetimeWrapper_338_io_in = _T_8261 & io_rPort_16_en_0; // @[package.scala 94:16:@56047.4]
  assign RetimeWrapper_339_clock = clock; // @[:@56053.4]
  assign RetimeWrapper_339_reset = reset; // @[:@56054.4]
  assign RetimeWrapper_339_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@56056.4]
  assign RetimeWrapper_339_io_in = _T_8565 & io_rPort_16_en_0; // @[package.scala 94:16:@56055.4]
  assign RetimeWrapper_340_clock = clock; // @[:@56141.4]
  assign RetimeWrapper_340_reset = reset; // @[:@56142.4]
  assign RetimeWrapper_340_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56144.4]
  assign RetimeWrapper_340_io_in = _T_2795 & io_rPort_17_en_0; // @[package.scala 94:16:@56143.4]
  assign RetimeWrapper_341_clock = clock; // @[:@56149.4]
  assign RetimeWrapper_341_reset = reset; // @[:@56150.4]
  assign RetimeWrapper_341_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56152.4]
  assign RetimeWrapper_341_io_in = _T_3099 & io_rPort_17_en_0; // @[package.scala 94:16:@56151.4]
  assign RetimeWrapper_342_clock = clock; // @[:@56157.4]
  assign RetimeWrapper_342_reset = reset; // @[:@56158.4]
  assign RetimeWrapper_342_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56160.4]
  assign RetimeWrapper_342_io_in = _T_3403 & io_rPort_17_en_0; // @[package.scala 94:16:@56159.4]
  assign RetimeWrapper_343_clock = clock; // @[:@56165.4]
  assign RetimeWrapper_343_reset = reset; // @[:@56166.4]
  assign RetimeWrapper_343_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56168.4]
  assign RetimeWrapper_343_io_in = _T_3707 & io_rPort_17_en_0; // @[package.scala 94:16:@56167.4]
  assign RetimeWrapper_344_clock = clock; // @[:@56173.4]
  assign RetimeWrapper_344_reset = reset; // @[:@56174.4]
  assign RetimeWrapper_344_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56176.4]
  assign RetimeWrapper_344_io_in = _T_4011 & io_rPort_17_en_0; // @[package.scala 94:16:@56175.4]
  assign RetimeWrapper_345_clock = clock; // @[:@56181.4]
  assign RetimeWrapper_345_reset = reset; // @[:@56182.4]
  assign RetimeWrapper_345_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56184.4]
  assign RetimeWrapper_345_io_in = _T_4315 & io_rPort_17_en_0; // @[package.scala 94:16:@56183.4]
  assign RetimeWrapper_346_clock = clock; // @[:@56189.4]
  assign RetimeWrapper_346_reset = reset; // @[:@56190.4]
  assign RetimeWrapper_346_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56192.4]
  assign RetimeWrapper_346_io_in = _T_4619 & io_rPort_17_en_0; // @[package.scala 94:16:@56191.4]
  assign RetimeWrapper_347_clock = clock; // @[:@56197.4]
  assign RetimeWrapper_347_reset = reset; // @[:@56198.4]
  assign RetimeWrapper_347_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56200.4]
  assign RetimeWrapper_347_io_in = _T_4923 & io_rPort_17_en_0; // @[package.scala 94:16:@56199.4]
  assign RetimeWrapper_348_clock = clock; // @[:@56205.4]
  assign RetimeWrapper_348_reset = reset; // @[:@56206.4]
  assign RetimeWrapper_348_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56208.4]
  assign RetimeWrapper_348_io_in = _T_5227 & io_rPort_17_en_0; // @[package.scala 94:16:@56207.4]
  assign RetimeWrapper_349_clock = clock; // @[:@56213.4]
  assign RetimeWrapper_349_reset = reset; // @[:@56214.4]
  assign RetimeWrapper_349_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56216.4]
  assign RetimeWrapper_349_io_in = _T_5531 & io_rPort_17_en_0; // @[package.scala 94:16:@56215.4]
  assign RetimeWrapper_350_clock = clock; // @[:@56221.4]
  assign RetimeWrapper_350_reset = reset; // @[:@56222.4]
  assign RetimeWrapper_350_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56224.4]
  assign RetimeWrapper_350_io_in = _T_5835 & io_rPort_17_en_0; // @[package.scala 94:16:@56223.4]
  assign RetimeWrapper_351_clock = clock; // @[:@56229.4]
  assign RetimeWrapper_351_reset = reset; // @[:@56230.4]
  assign RetimeWrapper_351_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56232.4]
  assign RetimeWrapper_351_io_in = _T_6139 & io_rPort_17_en_0; // @[package.scala 94:16:@56231.4]
  assign RetimeWrapper_352_clock = clock; // @[:@56237.4]
  assign RetimeWrapper_352_reset = reset; // @[:@56238.4]
  assign RetimeWrapper_352_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56240.4]
  assign RetimeWrapper_352_io_in = _T_6443 & io_rPort_17_en_0; // @[package.scala 94:16:@56239.4]
  assign RetimeWrapper_353_clock = clock; // @[:@56245.4]
  assign RetimeWrapper_353_reset = reset; // @[:@56246.4]
  assign RetimeWrapper_353_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56248.4]
  assign RetimeWrapper_353_io_in = _T_6747 & io_rPort_17_en_0; // @[package.scala 94:16:@56247.4]
  assign RetimeWrapper_354_clock = clock; // @[:@56253.4]
  assign RetimeWrapper_354_reset = reset; // @[:@56254.4]
  assign RetimeWrapper_354_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56256.4]
  assign RetimeWrapper_354_io_in = _T_7051 & io_rPort_17_en_0; // @[package.scala 94:16:@56255.4]
  assign RetimeWrapper_355_clock = clock; // @[:@56261.4]
  assign RetimeWrapper_355_reset = reset; // @[:@56262.4]
  assign RetimeWrapper_355_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56264.4]
  assign RetimeWrapper_355_io_in = _T_7355 & io_rPort_17_en_0; // @[package.scala 94:16:@56263.4]
  assign RetimeWrapper_356_clock = clock; // @[:@56269.4]
  assign RetimeWrapper_356_reset = reset; // @[:@56270.4]
  assign RetimeWrapper_356_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56272.4]
  assign RetimeWrapper_356_io_in = _T_7659 & io_rPort_17_en_0; // @[package.scala 94:16:@56271.4]
  assign RetimeWrapper_357_clock = clock; // @[:@56277.4]
  assign RetimeWrapper_357_reset = reset; // @[:@56278.4]
  assign RetimeWrapper_357_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56280.4]
  assign RetimeWrapper_357_io_in = _T_7963 & io_rPort_17_en_0; // @[package.scala 94:16:@56279.4]
  assign RetimeWrapper_358_clock = clock; // @[:@56285.4]
  assign RetimeWrapper_358_reset = reset; // @[:@56286.4]
  assign RetimeWrapper_358_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56288.4]
  assign RetimeWrapper_358_io_in = _T_8267 & io_rPort_17_en_0; // @[package.scala 94:16:@56287.4]
  assign RetimeWrapper_359_clock = clock; // @[:@56293.4]
  assign RetimeWrapper_359_reset = reset; // @[:@56294.4]
  assign RetimeWrapper_359_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@56296.4]
  assign RetimeWrapper_359_io_in = _T_8571 & io_rPort_17_en_0; // @[package.scala 94:16:@56295.4]
  assign RetimeWrapper_360_clock = clock; // @[:@56381.4]
  assign RetimeWrapper_360_reset = reset; // @[:@56382.4]
  assign RetimeWrapper_360_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56384.4]
  assign RetimeWrapper_360_io_in = _T_2929 & io_rPort_18_en_0; // @[package.scala 94:16:@56383.4]
  assign RetimeWrapper_361_clock = clock; // @[:@56389.4]
  assign RetimeWrapper_361_reset = reset; // @[:@56390.4]
  assign RetimeWrapper_361_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56392.4]
  assign RetimeWrapper_361_io_in = _T_3233 & io_rPort_18_en_0; // @[package.scala 94:16:@56391.4]
  assign RetimeWrapper_362_clock = clock; // @[:@56397.4]
  assign RetimeWrapper_362_reset = reset; // @[:@56398.4]
  assign RetimeWrapper_362_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56400.4]
  assign RetimeWrapper_362_io_in = _T_3537 & io_rPort_18_en_0; // @[package.scala 94:16:@56399.4]
  assign RetimeWrapper_363_clock = clock; // @[:@56405.4]
  assign RetimeWrapper_363_reset = reset; // @[:@56406.4]
  assign RetimeWrapper_363_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56408.4]
  assign RetimeWrapper_363_io_in = _T_3841 & io_rPort_18_en_0; // @[package.scala 94:16:@56407.4]
  assign RetimeWrapper_364_clock = clock; // @[:@56413.4]
  assign RetimeWrapper_364_reset = reset; // @[:@56414.4]
  assign RetimeWrapper_364_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56416.4]
  assign RetimeWrapper_364_io_in = _T_4145 & io_rPort_18_en_0; // @[package.scala 94:16:@56415.4]
  assign RetimeWrapper_365_clock = clock; // @[:@56421.4]
  assign RetimeWrapper_365_reset = reset; // @[:@56422.4]
  assign RetimeWrapper_365_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56424.4]
  assign RetimeWrapper_365_io_in = _T_4449 & io_rPort_18_en_0; // @[package.scala 94:16:@56423.4]
  assign RetimeWrapper_366_clock = clock; // @[:@56429.4]
  assign RetimeWrapper_366_reset = reset; // @[:@56430.4]
  assign RetimeWrapper_366_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56432.4]
  assign RetimeWrapper_366_io_in = _T_4753 & io_rPort_18_en_0; // @[package.scala 94:16:@56431.4]
  assign RetimeWrapper_367_clock = clock; // @[:@56437.4]
  assign RetimeWrapper_367_reset = reset; // @[:@56438.4]
  assign RetimeWrapper_367_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56440.4]
  assign RetimeWrapper_367_io_in = _T_5057 & io_rPort_18_en_0; // @[package.scala 94:16:@56439.4]
  assign RetimeWrapper_368_clock = clock; // @[:@56445.4]
  assign RetimeWrapper_368_reset = reset; // @[:@56446.4]
  assign RetimeWrapper_368_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56448.4]
  assign RetimeWrapper_368_io_in = _T_5361 & io_rPort_18_en_0; // @[package.scala 94:16:@56447.4]
  assign RetimeWrapper_369_clock = clock; // @[:@56453.4]
  assign RetimeWrapper_369_reset = reset; // @[:@56454.4]
  assign RetimeWrapper_369_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56456.4]
  assign RetimeWrapper_369_io_in = _T_5665 & io_rPort_18_en_0; // @[package.scala 94:16:@56455.4]
  assign RetimeWrapper_370_clock = clock; // @[:@56461.4]
  assign RetimeWrapper_370_reset = reset; // @[:@56462.4]
  assign RetimeWrapper_370_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56464.4]
  assign RetimeWrapper_370_io_in = _T_5969 & io_rPort_18_en_0; // @[package.scala 94:16:@56463.4]
  assign RetimeWrapper_371_clock = clock; // @[:@56469.4]
  assign RetimeWrapper_371_reset = reset; // @[:@56470.4]
  assign RetimeWrapper_371_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56472.4]
  assign RetimeWrapper_371_io_in = _T_6273 & io_rPort_18_en_0; // @[package.scala 94:16:@56471.4]
  assign RetimeWrapper_372_clock = clock; // @[:@56477.4]
  assign RetimeWrapper_372_reset = reset; // @[:@56478.4]
  assign RetimeWrapper_372_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56480.4]
  assign RetimeWrapper_372_io_in = _T_6577 & io_rPort_18_en_0; // @[package.scala 94:16:@56479.4]
  assign RetimeWrapper_373_clock = clock; // @[:@56485.4]
  assign RetimeWrapper_373_reset = reset; // @[:@56486.4]
  assign RetimeWrapper_373_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56488.4]
  assign RetimeWrapper_373_io_in = _T_6881 & io_rPort_18_en_0; // @[package.scala 94:16:@56487.4]
  assign RetimeWrapper_374_clock = clock; // @[:@56493.4]
  assign RetimeWrapper_374_reset = reset; // @[:@56494.4]
  assign RetimeWrapper_374_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56496.4]
  assign RetimeWrapper_374_io_in = _T_7185 & io_rPort_18_en_0; // @[package.scala 94:16:@56495.4]
  assign RetimeWrapper_375_clock = clock; // @[:@56501.4]
  assign RetimeWrapper_375_reset = reset; // @[:@56502.4]
  assign RetimeWrapper_375_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56504.4]
  assign RetimeWrapper_375_io_in = _T_7489 & io_rPort_18_en_0; // @[package.scala 94:16:@56503.4]
  assign RetimeWrapper_376_clock = clock; // @[:@56509.4]
  assign RetimeWrapper_376_reset = reset; // @[:@56510.4]
  assign RetimeWrapper_376_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56512.4]
  assign RetimeWrapper_376_io_in = _T_7793 & io_rPort_18_en_0; // @[package.scala 94:16:@56511.4]
  assign RetimeWrapper_377_clock = clock; // @[:@56517.4]
  assign RetimeWrapper_377_reset = reset; // @[:@56518.4]
  assign RetimeWrapper_377_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56520.4]
  assign RetimeWrapper_377_io_in = _T_8097 & io_rPort_18_en_0; // @[package.scala 94:16:@56519.4]
  assign RetimeWrapper_378_clock = clock; // @[:@56525.4]
  assign RetimeWrapper_378_reset = reset; // @[:@56526.4]
  assign RetimeWrapper_378_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56528.4]
  assign RetimeWrapper_378_io_in = _T_8401 & io_rPort_18_en_0; // @[package.scala 94:16:@56527.4]
  assign RetimeWrapper_379_clock = clock; // @[:@56533.4]
  assign RetimeWrapper_379_reset = reset; // @[:@56534.4]
  assign RetimeWrapper_379_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@56536.4]
  assign RetimeWrapper_379_io_in = _T_8705 & io_rPort_18_en_0; // @[package.scala 94:16:@56535.4]
  assign RetimeWrapper_380_clock = clock; // @[:@56621.4]
  assign RetimeWrapper_380_reset = reset; // @[:@56622.4]
  assign RetimeWrapper_380_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56624.4]
  assign RetimeWrapper_380_io_in = _T_2801 & io_rPort_19_en_0; // @[package.scala 94:16:@56623.4]
  assign RetimeWrapper_381_clock = clock; // @[:@56629.4]
  assign RetimeWrapper_381_reset = reset; // @[:@56630.4]
  assign RetimeWrapper_381_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56632.4]
  assign RetimeWrapper_381_io_in = _T_3105 & io_rPort_19_en_0; // @[package.scala 94:16:@56631.4]
  assign RetimeWrapper_382_clock = clock; // @[:@56637.4]
  assign RetimeWrapper_382_reset = reset; // @[:@56638.4]
  assign RetimeWrapper_382_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56640.4]
  assign RetimeWrapper_382_io_in = _T_3409 & io_rPort_19_en_0; // @[package.scala 94:16:@56639.4]
  assign RetimeWrapper_383_clock = clock; // @[:@56645.4]
  assign RetimeWrapper_383_reset = reset; // @[:@56646.4]
  assign RetimeWrapper_383_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56648.4]
  assign RetimeWrapper_383_io_in = _T_3713 & io_rPort_19_en_0; // @[package.scala 94:16:@56647.4]
  assign RetimeWrapper_384_clock = clock; // @[:@56653.4]
  assign RetimeWrapper_384_reset = reset; // @[:@56654.4]
  assign RetimeWrapper_384_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56656.4]
  assign RetimeWrapper_384_io_in = _T_4017 & io_rPort_19_en_0; // @[package.scala 94:16:@56655.4]
  assign RetimeWrapper_385_clock = clock; // @[:@56661.4]
  assign RetimeWrapper_385_reset = reset; // @[:@56662.4]
  assign RetimeWrapper_385_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56664.4]
  assign RetimeWrapper_385_io_in = _T_4321 & io_rPort_19_en_0; // @[package.scala 94:16:@56663.4]
  assign RetimeWrapper_386_clock = clock; // @[:@56669.4]
  assign RetimeWrapper_386_reset = reset; // @[:@56670.4]
  assign RetimeWrapper_386_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56672.4]
  assign RetimeWrapper_386_io_in = _T_4625 & io_rPort_19_en_0; // @[package.scala 94:16:@56671.4]
  assign RetimeWrapper_387_clock = clock; // @[:@56677.4]
  assign RetimeWrapper_387_reset = reset; // @[:@56678.4]
  assign RetimeWrapper_387_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56680.4]
  assign RetimeWrapper_387_io_in = _T_4929 & io_rPort_19_en_0; // @[package.scala 94:16:@56679.4]
  assign RetimeWrapper_388_clock = clock; // @[:@56685.4]
  assign RetimeWrapper_388_reset = reset; // @[:@56686.4]
  assign RetimeWrapper_388_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56688.4]
  assign RetimeWrapper_388_io_in = _T_5233 & io_rPort_19_en_0; // @[package.scala 94:16:@56687.4]
  assign RetimeWrapper_389_clock = clock; // @[:@56693.4]
  assign RetimeWrapper_389_reset = reset; // @[:@56694.4]
  assign RetimeWrapper_389_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56696.4]
  assign RetimeWrapper_389_io_in = _T_5537 & io_rPort_19_en_0; // @[package.scala 94:16:@56695.4]
  assign RetimeWrapper_390_clock = clock; // @[:@56701.4]
  assign RetimeWrapper_390_reset = reset; // @[:@56702.4]
  assign RetimeWrapper_390_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56704.4]
  assign RetimeWrapper_390_io_in = _T_5841 & io_rPort_19_en_0; // @[package.scala 94:16:@56703.4]
  assign RetimeWrapper_391_clock = clock; // @[:@56709.4]
  assign RetimeWrapper_391_reset = reset; // @[:@56710.4]
  assign RetimeWrapper_391_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56712.4]
  assign RetimeWrapper_391_io_in = _T_6145 & io_rPort_19_en_0; // @[package.scala 94:16:@56711.4]
  assign RetimeWrapper_392_clock = clock; // @[:@56717.4]
  assign RetimeWrapper_392_reset = reset; // @[:@56718.4]
  assign RetimeWrapper_392_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56720.4]
  assign RetimeWrapper_392_io_in = _T_6449 & io_rPort_19_en_0; // @[package.scala 94:16:@56719.4]
  assign RetimeWrapper_393_clock = clock; // @[:@56725.4]
  assign RetimeWrapper_393_reset = reset; // @[:@56726.4]
  assign RetimeWrapper_393_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56728.4]
  assign RetimeWrapper_393_io_in = _T_6753 & io_rPort_19_en_0; // @[package.scala 94:16:@56727.4]
  assign RetimeWrapper_394_clock = clock; // @[:@56733.4]
  assign RetimeWrapper_394_reset = reset; // @[:@56734.4]
  assign RetimeWrapper_394_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56736.4]
  assign RetimeWrapper_394_io_in = _T_7057 & io_rPort_19_en_0; // @[package.scala 94:16:@56735.4]
  assign RetimeWrapper_395_clock = clock; // @[:@56741.4]
  assign RetimeWrapper_395_reset = reset; // @[:@56742.4]
  assign RetimeWrapper_395_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56744.4]
  assign RetimeWrapper_395_io_in = _T_7361 & io_rPort_19_en_0; // @[package.scala 94:16:@56743.4]
  assign RetimeWrapper_396_clock = clock; // @[:@56749.4]
  assign RetimeWrapper_396_reset = reset; // @[:@56750.4]
  assign RetimeWrapper_396_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56752.4]
  assign RetimeWrapper_396_io_in = _T_7665 & io_rPort_19_en_0; // @[package.scala 94:16:@56751.4]
  assign RetimeWrapper_397_clock = clock; // @[:@56757.4]
  assign RetimeWrapper_397_reset = reset; // @[:@56758.4]
  assign RetimeWrapper_397_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56760.4]
  assign RetimeWrapper_397_io_in = _T_7969 & io_rPort_19_en_0; // @[package.scala 94:16:@56759.4]
  assign RetimeWrapper_398_clock = clock; // @[:@56765.4]
  assign RetimeWrapper_398_reset = reset; // @[:@56766.4]
  assign RetimeWrapper_398_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56768.4]
  assign RetimeWrapper_398_io_in = _T_8273 & io_rPort_19_en_0; // @[package.scala 94:16:@56767.4]
  assign RetimeWrapper_399_clock = clock; // @[:@56773.4]
  assign RetimeWrapper_399_reset = reset; // @[:@56774.4]
  assign RetimeWrapper_399_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@56776.4]
  assign RetimeWrapper_399_io_in = _T_8577 & io_rPort_19_en_0; // @[package.scala 94:16:@56775.4]
  assign RetimeWrapper_400_clock = clock; // @[:@56861.4]
  assign RetimeWrapper_400_reset = reset; // @[:@56862.4]
  assign RetimeWrapper_400_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56864.4]
  assign RetimeWrapper_400_io_in = _T_2935 & io_rPort_20_en_0; // @[package.scala 94:16:@56863.4]
  assign RetimeWrapper_401_clock = clock; // @[:@56869.4]
  assign RetimeWrapper_401_reset = reset; // @[:@56870.4]
  assign RetimeWrapper_401_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56872.4]
  assign RetimeWrapper_401_io_in = _T_3239 & io_rPort_20_en_0; // @[package.scala 94:16:@56871.4]
  assign RetimeWrapper_402_clock = clock; // @[:@56877.4]
  assign RetimeWrapper_402_reset = reset; // @[:@56878.4]
  assign RetimeWrapper_402_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56880.4]
  assign RetimeWrapper_402_io_in = _T_3543 & io_rPort_20_en_0; // @[package.scala 94:16:@56879.4]
  assign RetimeWrapper_403_clock = clock; // @[:@56885.4]
  assign RetimeWrapper_403_reset = reset; // @[:@56886.4]
  assign RetimeWrapper_403_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56888.4]
  assign RetimeWrapper_403_io_in = _T_3847 & io_rPort_20_en_0; // @[package.scala 94:16:@56887.4]
  assign RetimeWrapper_404_clock = clock; // @[:@56893.4]
  assign RetimeWrapper_404_reset = reset; // @[:@56894.4]
  assign RetimeWrapper_404_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56896.4]
  assign RetimeWrapper_404_io_in = _T_4151 & io_rPort_20_en_0; // @[package.scala 94:16:@56895.4]
  assign RetimeWrapper_405_clock = clock; // @[:@56901.4]
  assign RetimeWrapper_405_reset = reset; // @[:@56902.4]
  assign RetimeWrapper_405_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56904.4]
  assign RetimeWrapper_405_io_in = _T_4455 & io_rPort_20_en_0; // @[package.scala 94:16:@56903.4]
  assign RetimeWrapper_406_clock = clock; // @[:@56909.4]
  assign RetimeWrapper_406_reset = reset; // @[:@56910.4]
  assign RetimeWrapper_406_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56912.4]
  assign RetimeWrapper_406_io_in = _T_4759 & io_rPort_20_en_0; // @[package.scala 94:16:@56911.4]
  assign RetimeWrapper_407_clock = clock; // @[:@56917.4]
  assign RetimeWrapper_407_reset = reset; // @[:@56918.4]
  assign RetimeWrapper_407_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56920.4]
  assign RetimeWrapper_407_io_in = _T_5063 & io_rPort_20_en_0; // @[package.scala 94:16:@56919.4]
  assign RetimeWrapper_408_clock = clock; // @[:@56925.4]
  assign RetimeWrapper_408_reset = reset; // @[:@56926.4]
  assign RetimeWrapper_408_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56928.4]
  assign RetimeWrapper_408_io_in = _T_5367 & io_rPort_20_en_0; // @[package.scala 94:16:@56927.4]
  assign RetimeWrapper_409_clock = clock; // @[:@56933.4]
  assign RetimeWrapper_409_reset = reset; // @[:@56934.4]
  assign RetimeWrapper_409_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56936.4]
  assign RetimeWrapper_409_io_in = _T_5671 & io_rPort_20_en_0; // @[package.scala 94:16:@56935.4]
  assign RetimeWrapper_410_clock = clock; // @[:@56941.4]
  assign RetimeWrapper_410_reset = reset; // @[:@56942.4]
  assign RetimeWrapper_410_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56944.4]
  assign RetimeWrapper_410_io_in = _T_5975 & io_rPort_20_en_0; // @[package.scala 94:16:@56943.4]
  assign RetimeWrapper_411_clock = clock; // @[:@56949.4]
  assign RetimeWrapper_411_reset = reset; // @[:@56950.4]
  assign RetimeWrapper_411_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56952.4]
  assign RetimeWrapper_411_io_in = _T_6279 & io_rPort_20_en_0; // @[package.scala 94:16:@56951.4]
  assign RetimeWrapper_412_clock = clock; // @[:@56957.4]
  assign RetimeWrapper_412_reset = reset; // @[:@56958.4]
  assign RetimeWrapper_412_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56960.4]
  assign RetimeWrapper_412_io_in = _T_6583 & io_rPort_20_en_0; // @[package.scala 94:16:@56959.4]
  assign RetimeWrapper_413_clock = clock; // @[:@56965.4]
  assign RetimeWrapper_413_reset = reset; // @[:@56966.4]
  assign RetimeWrapper_413_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56968.4]
  assign RetimeWrapper_413_io_in = _T_6887 & io_rPort_20_en_0; // @[package.scala 94:16:@56967.4]
  assign RetimeWrapper_414_clock = clock; // @[:@56973.4]
  assign RetimeWrapper_414_reset = reset; // @[:@56974.4]
  assign RetimeWrapper_414_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56976.4]
  assign RetimeWrapper_414_io_in = _T_7191 & io_rPort_20_en_0; // @[package.scala 94:16:@56975.4]
  assign RetimeWrapper_415_clock = clock; // @[:@56981.4]
  assign RetimeWrapper_415_reset = reset; // @[:@56982.4]
  assign RetimeWrapper_415_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56984.4]
  assign RetimeWrapper_415_io_in = _T_7495 & io_rPort_20_en_0; // @[package.scala 94:16:@56983.4]
  assign RetimeWrapper_416_clock = clock; // @[:@56989.4]
  assign RetimeWrapper_416_reset = reset; // @[:@56990.4]
  assign RetimeWrapper_416_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@56992.4]
  assign RetimeWrapper_416_io_in = _T_7799 & io_rPort_20_en_0; // @[package.scala 94:16:@56991.4]
  assign RetimeWrapper_417_clock = clock; // @[:@56997.4]
  assign RetimeWrapper_417_reset = reset; // @[:@56998.4]
  assign RetimeWrapper_417_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@57000.4]
  assign RetimeWrapper_417_io_in = _T_8103 & io_rPort_20_en_0; // @[package.scala 94:16:@56999.4]
  assign RetimeWrapper_418_clock = clock; // @[:@57005.4]
  assign RetimeWrapper_418_reset = reset; // @[:@57006.4]
  assign RetimeWrapper_418_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@57008.4]
  assign RetimeWrapper_418_io_in = _T_8407 & io_rPort_20_en_0; // @[package.scala 94:16:@57007.4]
  assign RetimeWrapper_419_clock = clock; // @[:@57013.4]
  assign RetimeWrapper_419_reset = reset; // @[:@57014.4]
  assign RetimeWrapper_419_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@57016.4]
  assign RetimeWrapper_419_io_in = _T_8711 & io_rPort_20_en_0; // @[package.scala 94:16:@57015.4]
  assign RetimeWrapper_420_clock = clock; // @[:@57101.4]
  assign RetimeWrapper_420_reset = reset; // @[:@57102.4]
  assign RetimeWrapper_420_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57104.4]
  assign RetimeWrapper_420_io_in = _T_2941 & io_rPort_21_en_0; // @[package.scala 94:16:@57103.4]
  assign RetimeWrapper_421_clock = clock; // @[:@57109.4]
  assign RetimeWrapper_421_reset = reset; // @[:@57110.4]
  assign RetimeWrapper_421_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57112.4]
  assign RetimeWrapper_421_io_in = _T_3245 & io_rPort_21_en_0; // @[package.scala 94:16:@57111.4]
  assign RetimeWrapper_422_clock = clock; // @[:@57117.4]
  assign RetimeWrapper_422_reset = reset; // @[:@57118.4]
  assign RetimeWrapper_422_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57120.4]
  assign RetimeWrapper_422_io_in = _T_3549 & io_rPort_21_en_0; // @[package.scala 94:16:@57119.4]
  assign RetimeWrapper_423_clock = clock; // @[:@57125.4]
  assign RetimeWrapper_423_reset = reset; // @[:@57126.4]
  assign RetimeWrapper_423_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57128.4]
  assign RetimeWrapper_423_io_in = _T_3853 & io_rPort_21_en_0; // @[package.scala 94:16:@57127.4]
  assign RetimeWrapper_424_clock = clock; // @[:@57133.4]
  assign RetimeWrapper_424_reset = reset; // @[:@57134.4]
  assign RetimeWrapper_424_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57136.4]
  assign RetimeWrapper_424_io_in = _T_4157 & io_rPort_21_en_0; // @[package.scala 94:16:@57135.4]
  assign RetimeWrapper_425_clock = clock; // @[:@57141.4]
  assign RetimeWrapper_425_reset = reset; // @[:@57142.4]
  assign RetimeWrapper_425_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57144.4]
  assign RetimeWrapper_425_io_in = _T_4461 & io_rPort_21_en_0; // @[package.scala 94:16:@57143.4]
  assign RetimeWrapper_426_clock = clock; // @[:@57149.4]
  assign RetimeWrapper_426_reset = reset; // @[:@57150.4]
  assign RetimeWrapper_426_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57152.4]
  assign RetimeWrapper_426_io_in = _T_4765 & io_rPort_21_en_0; // @[package.scala 94:16:@57151.4]
  assign RetimeWrapper_427_clock = clock; // @[:@57157.4]
  assign RetimeWrapper_427_reset = reset; // @[:@57158.4]
  assign RetimeWrapper_427_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57160.4]
  assign RetimeWrapper_427_io_in = _T_5069 & io_rPort_21_en_0; // @[package.scala 94:16:@57159.4]
  assign RetimeWrapper_428_clock = clock; // @[:@57165.4]
  assign RetimeWrapper_428_reset = reset; // @[:@57166.4]
  assign RetimeWrapper_428_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57168.4]
  assign RetimeWrapper_428_io_in = _T_5373 & io_rPort_21_en_0; // @[package.scala 94:16:@57167.4]
  assign RetimeWrapper_429_clock = clock; // @[:@57173.4]
  assign RetimeWrapper_429_reset = reset; // @[:@57174.4]
  assign RetimeWrapper_429_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57176.4]
  assign RetimeWrapper_429_io_in = _T_5677 & io_rPort_21_en_0; // @[package.scala 94:16:@57175.4]
  assign RetimeWrapper_430_clock = clock; // @[:@57181.4]
  assign RetimeWrapper_430_reset = reset; // @[:@57182.4]
  assign RetimeWrapper_430_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57184.4]
  assign RetimeWrapper_430_io_in = _T_5981 & io_rPort_21_en_0; // @[package.scala 94:16:@57183.4]
  assign RetimeWrapper_431_clock = clock; // @[:@57189.4]
  assign RetimeWrapper_431_reset = reset; // @[:@57190.4]
  assign RetimeWrapper_431_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57192.4]
  assign RetimeWrapper_431_io_in = _T_6285 & io_rPort_21_en_0; // @[package.scala 94:16:@57191.4]
  assign RetimeWrapper_432_clock = clock; // @[:@57197.4]
  assign RetimeWrapper_432_reset = reset; // @[:@57198.4]
  assign RetimeWrapper_432_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57200.4]
  assign RetimeWrapper_432_io_in = _T_6589 & io_rPort_21_en_0; // @[package.scala 94:16:@57199.4]
  assign RetimeWrapper_433_clock = clock; // @[:@57205.4]
  assign RetimeWrapper_433_reset = reset; // @[:@57206.4]
  assign RetimeWrapper_433_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57208.4]
  assign RetimeWrapper_433_io_in = _T_6893 & io_rPort_21_en_0; // @[package.scala 94:16:@57207.4]
  assign RetimeWrapper_434_clock = clock; // @[:@57213.4]
  assign RetimeWrapper_434_reset = reset; // @[:@57214.4]
  assign RetimeWrapper_434_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57216.4]
  assign RetimeWrapper_434_io_in = _T_7197 & io_rPort_21_en_0; // @[package.scala 94:16:@57215.4]
  assign RetimeWrapper_435_clock = clock; // @[:@57221.4]
  assign RetimeWrapper_435_reset = reset; // @[:@57222.4]
  assign RetimeWrapper_435_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57224.4]
  assign RetimeWrapper_435_io_in = _T_7501 & io_rPort_21_en_0; // @[package.scala 94:16:@57223.4]
  assign RetimeWrapper_436_clock = clock; // @[:@57229.4]
  assign RetimeWrapper_436_reset = reset; // @[:@57230.4]
  assign RetimeWrapper_436_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57232.4]
  assign RetimeWrapper_436_io_in = _T_7805 & io_rPort_21_en_0; // @[package.scala 94:16:@57231.4]
  assign RetimeWrapper_437_clock = clock; // @[:@57237.4]
  assign RetimeWrapper_437_reset = reset; // @[:@57238.4]
  assign RetimeWrapper_437_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57240.4]
  assign RetimeWrapper_437_io_in = _T_8109 & io_rPort_21_en_0; // @[package.scala 94:16:@57239.4]
  assign RetimeWrapper_438_clock = clock; // @[:@57245.4]
  assign RetimeWrapper_438_reset = reset; // @[:@57246.4]
  assign RetimeWrapper_438_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57248.4]
  assign RetimeWrapper_438_io_in = _T_8413 & io_rPort_21_en_0; // @[package.scala 94:16:@57247.4]
  assign RetimeWrapper_439_clock = clock; // @[:@57253.4]
  assign RetimeWrapper_439_reset = reset; // @[:@57254.4]
  assign RetimeWrapper_439_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@57256.4]
  assign RetimeWrapper_439_io_in = _T_8717 & io_rPort_21_en_0; // @[package.scala 94:16:@57255.4]
  assign RetimeWrapper_440_clock = clock; // @[:@57341.4]
  assign RetimeWrapper_440_reset = reset; // @[:@57342.4]
  assign RetimeWrapper_440_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57344.4]
  assign RetimeWrapper_440_io_in = _T_2807 & io_rPort_22_en_0; // @[package.scala 94:16:@57343.4]
  assign RetimeWrapper_441_clock = clock; // @[:@57349.4]
  assign RetimeWrapper_441_reset = reset; // @[:@57350.4]
  assign RetimeWrapper_441_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57352.4]
  assign RetimeWrapper_441_io_in = _T_3111 & io_rPort_22_en_0; // @[package.scala 94:16:@57351.4]
  assign RetimeWrapper_442_clock = clock; // @[:@57357.4]
  assign RetimeWrapper_442_reset = reset; // @[:@57358.4]
  assign RetimeWrapper_442_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57360.4]
  assign RetimeWrapper_442_io_in = _T_3415 & io_rPort_22_en_0; // @[package.scala 94:16:@57359.4]
  assign RetimeWrapper_443_clock = clock; // @[:@57365.4]
  assign RetimeWrapper_443_reset = reset; // @[:@57366.4]
  assign RetimeWrapper_443_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57368.4]
  assign RetimeWrapper_443_io_in = _T_3719 & io_rPort_22_en_0; // @[package.scala 94:16:@57367.4]
  assign RetimeWrapper_444_clock = clock; // @[:@57373.4]
  assign RetimeWrapper_444_reset = reset; // @[:@57374.4]
  assign RetimeWrapper_444_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57376.4]
  assign RetimeWrapper_444_io_in = _T_4023 & io_rPort_22_en_0; // @[package.scala 94:16:@57375.4]
  assign RetimeWrapper_445_clock = clock; // @[:@57381.4]
  assign RetimeWrapper_445_reset = reset; // @[:@57382.4]
  assign RetimeWrapper_445_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57384.4]
  assign RetimeWrapper_445_io_in = _T_4327 & io_rPort_22_en_0; // @[package.scala 94:16:@57383.4]
  assign RetimeWrapper_446_clock = clock; // @[:@57389.4]
  assign RetimeWrapper_446_reset = reset; // @[:@57390.4]
  assign RetimeWrapper_446_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57392.4]
  assign RetimeWrapper_446_io_in = _T_4631 & io_rPort_22_en_0; // @[package.scala 94:16:@57391.4]
  assign RetimeWrapper_447_clock = clock; // @[:@57397.4]
  assign RetimeWrapper_447_reset = reset; // @[:@57398.4]
  assign RetimeWrapper_447_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57400.4]
  assign RetimeWrapper_447_io_in = _T_4935 & io_rPort_22_en_0; // @[package.scala 94:16:@57399.4]
  assign RetimeWrapper_448_clock = clock; // @[:@57405.4]
  assign RetimeWrapper_448_reset = reset; // @[:@57406.4]
  assign RetimeWrapper_448_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57408.4]
  assign RetimeWrapper_448_io_in = _T_5239 & io_rPort_22_en_0; // @[package.scala 94:16:@57407.4]
  assign RetimeWrapper_449_clock = clock; // @[:@57413.4]
  assign RetimeWrapper_449_reset = reset; // @[:@57414.4]
  assign RetimeWrapper_449_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57416.4]
  assign RetimeWrapper_449_io_in = _T_5543 & io_rPort_22_en_0; // @[package.scala 94:16:@57415.4]
  assign RetimeWrapper_450_clock = clock; // @[:@57421.4]
  assign RetimeWrapper_450_reset = reset; // @[:@57422.4]
  assign RetimeWrapper_450_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57424.4]
  assign RetimeWrapper_450_io_in = _T_5847 & io_rPort_22_en_0; // @[package.scala 94:16:@57423.4]
  assign RetimeWrapper_451_clock = clock; // @[:@57429.4]
  assign RetimeWrapper_451_reset = reset; // @[:@57430.4]
  assign RetimeWrapper_451_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57432.4]
  assign RetimeWrapper_451_io_in = _T_6151 & io_rPort_22_en_0; // @[package.scala 94:16:@57431.4]
  assign RetimeWrapper_452_clock = clock; // @[:@57437.4]
  assign RetimeWrapper_452_reset = reset; // @[:@57438.4]
  assign RetimeWrapper_452_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57440.4]
  assign RetimeWrapper_452_io_in = _T_6455 & io_rPort_22_en_0; // @[package.scala 94:16:@57439.4]
  assign RetimeWrapper_453_clock = clock; // @[:@57445.4]
  assign RetimeWrapper_453_reset = reset; // @[:@57446.4]
  assign RetimeWrapper_453_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57448.4]
  assign RetimeWrapper_453_io_in = _T_6759 & io_rPort_22_en_0; // @[package.scala 94:16:@57447.4]
  assign RetimeWrapper_454_clock = clock; // @[:@57453.4]
  assign RetimeWrapper_454_reset = reset; // @[:@57454.4]
  assign RetimeWrapper_454_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57456.4]
  assign RetimeWrapper_454_io_in = _T_7063 & io_rPort_22_en_0; // @[package.scala 94:16:@57455.4]
  assign RetimeWrapper_455_clock = clock; // @[:@57461.4]
  assign RetimeWrapper_455_reset = reset; // @[:@57462.4]
  assign RetimeWrapper_455_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57464.4]
  assign RetimeWrapper_455_io_in = _T_7367 & io_rPort_22_en_0; // @[package.scala 94:16:@57463.4]
  assign RetimeWrapper_456_clock = clock; // @[:@57469.4]
  assign RetimeWrapper_456_reset = reset; // @[:@57470.4]
  assign RetimeWrapper_456_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57472.4]
  assign RetimeWrapper_456_io_in = _T_7671 & io_rPort_22_en_0; // @[package.scala 94:16:@57471.4]
  assign RetimeWrapper_457_clock = clock; // @[:@57477.4]
  assign RetimeWrapper_457_reset = reset; // @[:@57478.4]
  assign RetimeWrapper_457_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57480.4]
  assign RetimeWrapper_457_io_in = _T_7975 & io_rPort_22_en_0; // @[package.scala 94:16:@57479.4]
  assign RetimeWrapper_458_clock = clock; // @[:@57485.4]
  assign RetimeWrapper_458_reset = reset; // @[:@57486.4]
  assign RetimeWrapper_458_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57488.4]
  assign RetimeWrapper_458_io_in = _T_8279 & io_rPort_22_en_0; // @[package.scala 94:16:@57487.4]
  assign RetimeWrapper_459_clock = clock; // @[:@57493.4]
  assign RetimeWrapper_459_reset = reset; // @[:@57494.4]
  assign RetimeWrapper_459_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@57496.4]
  assign RetimeWrapper_459_io_in = _T_8583 & io_rPort_22_en_0; // @[package.scala 94:16:@57495.4]
  assign RetimeWrapper_460_clock = clock; // @[:@57581.4]
  assign RetimeWrapper_460_reset = reset; // @[:@57582.4]
  assign RetimeWrapper_460_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57584.4]
  assign RetimeWrapper_460_io_in = _T_2947 & io_rPort_23_en_0; // @[package.scala 94:16:@57583.4]
  assign RetimeWrapper_461_clock = clock; // @[:@57589.4]
  assign RetimeWrapper_461_reset = reset; // @[:@57590.4]
  assign RetimeWrapper_461_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57592.4]
  assign RetimeWrapper_461_io_in = _T_3251 & io_rPort_23_en_0; // @[package.scala 94:16:@57591.4]
  assign RetimeWrapper_462_clock = clock; // @[:@57597.4]
  assign RetimeWrapper_462_reset = reset; // @[:@57598.4]
  assign RetimeWrapper_462_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57600.4]
  assign RetimeWrapper_462_io_in = _T_3555 & io_rPort_23_en_0; // @[package.scala 94:16:@57599.4]
  assign RetimeWrapper_463_clock = clock; // @[:@57605.4]
  assign RetimeWrapper_463_reset = reset; // @[:@57606.4]
  assign RetimeWrapper_463_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57608.4]
  assign RetimeWrapper_463_io_in = _T_3859 & io_rPort_23_en_0; // @[package.scala 94:16:@57607.4]
  assign RetimeWrapper_464_clock = clock; // @[:@57613.4]
  assign RetimeWrapper_464_reset = reset; // @[:@57614.4]
  assign RetimeWrapper_464_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57616.4]
  assign RetimeWrapper_464_io_in = _T_4163 & io_rPort_23_en_0; // @[package.scala 94:16:@57615.4]
  assign RetimeWrapper_465_clock = clock; // @[:@57621.4]
  assign RetimeWrapper_465_reset = reset; // @[:@57622.4]
  assign RetimeWrapper_465_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57624.4]
  assign RetimeWrapper_465_io_in = _T_4467 & io_rPort_23_en_0; // @[package.scala 94:16:@57623.4]
  assign RetimeWrapper_466_clock = clock; // @[:@57629.4]
  assign RetimeWrapper_466_reset = reset; // @[:@57630.4]
  assign RetimeWrapper_466_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57632.4]
  assign RetimeWrapper_466_io_in = _T_4771 & io_rPort_23_en_0; // @[package.scala 94:16:@57631.4]
  assign RetimeWrapper_467_clock = clock; // @[:@57637.4]
  assign RetimeWrapper_467_reset = reset; // @[:@57638.4]
  assign RetimeWrapper_467_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57640.4]
  assign RetimeWrapper_467_io_in = _T_5075 & io_rPort_23_en_0; // @[package.scala 94:16:@57639.4]
  assign RetimeWrapper_468_clock = clock; // @[:@57645.4]
  assign RetimeWrapper_468_reset = reset; // @[:@57646.4]
  assign RetimeWrapper_468_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57648.4]
  assign RetimeWrapper_468_io_in = _T_5379 & io_rPort_23_en_0; // @[package.scala 94:16:@57647.4]
  assign RetimeWrapper_469_clock = clock; // @[:@57653.4]
  assign RetimeWrapper_469_reset = reset; // @[:@57654.4]
  assign RetimeWrapper_469_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57656.4]
  assign RetimeWrapper_469_io_in = _T_5683 & io_rPort_23_en_0; // @[package.scala 94:16:@57655.4]
  assign RetimeWrapper_470_clock = clock; // @[:@57661.4]
  assign RetimeWrapper_470_reset = reset; // @[:@57662.4]
  assign RetimeWrapper_470_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57664.4]
  assign RetimeWrapper_470_io_in = _T_5987 & io_rPort_23_en_0; // @[package.scala 94:16:@57663.4]
  assign RetimeWrapper_471_clock = clock; // @[:@57669.4]
  assign RetimeWrapper_471_reset = reset; // @[:@57670.4]
  assign RetimeWrapper_471_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57672.4]
  assign RetimeWrapper_471_io_in = _T_6291 & io_rPort_23_en_0; // @[package.scala 94:16:@57671.4]
  assign RetimeWrapper_472_clock = clock; // @[:@57677.4]
  assign RetimeWrapper_472_reset = reset; // @[:@57678.4]
  assign RetimeWrapper_472_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57680.4]
  assign RetimeWrapper_472_io_in = _T_6595 & io_rPort_23_en_0; // @[package.scala 94:16:@57679.4]
  assign RetimeWrapper_473_clock = clock; // @[:@57685.4]
  assign RetimeWrapper_473_reset = reset; // @[:@57686.4]
  assign RetimeWrapper_473_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57688.4]
  assign RetimeWrapper_473_io_in = _T_6899 & io_rPort_23_en_0; // @[package.scala 94:16:@57687.4]
  assign RetimeWrapper_474_clock = clock; // @[:@57693.4]
  assign RetimeWrapper_474_reset = reset; // @[:@57694.4]
  assign RetimeWrapper_474_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57696.4]
  assign RetimeWrapper_474_io_in = _T_7203 & io_rPort_23_en_0; // @[package.scala 94:16:@57695.4]
  assign RetimeWrapper_475_clock = clock; // @[:@57701.4]
  assign RetimeWrapper_475_reset = reset; // @[:@57702.4]
  assign RetimeWrapper_475_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57704.4]
  assign RetimeWrapper_475_io_in = _T_7507 & io_rPort_23_en_0; // @[package.scala 94:16:@57703.4]
  assign RetimeWrapper_476_clock = clock; // @[:@57709.4]
  assign RetimeWrapper_476_reset = reset; // @[:@57710.4]
  assign RetimeWrapper_476_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57712.4]
  assign RetimeWrapper_476_io_in = _T_7811 & io_rPort_23_en_0; // @[package.scala 94:16:@57711.4]
  assign RetimeWrapper_477_clock = clock; // @[:@57717.4]
  assign RetimeWrapper_477_reset = reset; // @[:@57718.4]
  assign RetimeWrapper_477_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57720.4]
  assign RetimeWrapper_477_io_in = _T_8115 & io_rPort_23_en_0; // @[package.scala 94:16:@57719.4]
  assign RetimeWrapper_478_clock = clock; // @[:@57725.4]
  assign RetimeWrapper_478_reset = reset; // @[:@57726.4]
  assign RetimeWrapper_478_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57728.4]
  assign RetimeWrapper_478_io_in = _T_8419 & io_rPort_23_en_0; // @[package.scala 94:16:@57727.4]
  assign RetimeWrapper_479_clock = clock; // @[:@57733.4]
  assign RetimeWrapper_479_reset = reset; // @[:@57734.4]
  assign RetimeWrapper_479_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@57736.4]
  assign RetimeWrapper_479_io_in = _T_8723 & io_rPort_23_en_0; // @[package.scala 94:16:@57735.4]
  assign RetimeWrapper_480_clock = clock; // @[:@57821.4]
  assign RetimeWrapper_480_reset = reset; // @[:@57822.4]
  assign RetimeWrapper_480_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57824.4]
  assign RetimeWrapper_480_io_in = _T_2953 & io_rPort_24_en_0; // @[package.scala 94:16:@57823.4]
  assign RetimeWrapper_481_clock = clock; // @[:@57829.4]
  assign RetimeWrapper_481_reset = reset; // @[:@57830.4]
  assign RetimeWrapper_481_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57832.4]
  assign RetimeWrapper_481_io_in = _T_3257 & io_rPort_24_en_0; // @[package.scala 94:16:@57831.4]
  assign RetimeWrapper_482_clock = clock; // @[:@57837.4]
  assign RetimeWrapper_482_reset = reset; // @[:@57838.4]
  assign RetimeWrapper_482_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57840.4]
  assign RetimeWrapper_482_io_in = _T_3561 & io_rPort_24_en_0; // @[package.scala 94:16:@57839.4]
  assign RetimeWrapper_483_clock = clock; // @[:@57845.4]
  assign RetimeWrapper_483_reset = reset; // @[:@57846.4]
  assign RetimeWrapper_483_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57848.4]
  assign RetimeWrapper_483_io_in = _T_3865 & io_rPort_24_en_0; // @[package.scala 94:16:@57847.4]
  assign RetimeWrapper_484_clock = clock; // @[:@57853.4]
  assign RetimeWrapper_484_reset = reset; // @[:@57854.4]
  assign RetimeWrapper_484_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57856.4]
  assign RetimeWrapper_484_io_in = _T_4169 & io_rPort_24_en_0; // @[package.scala 94:16:@57855.4]
  assign RetimeWrapper_485_clock = clock; // @[:@57861.4]
  assign RetimeWrapper_485_reset = reset; // @[:@57862.4]
  assign RetimeWrapper_485_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57864.4]
  assign RetimeWrapper_485_io_in = _T_4473 & io_rPort_24_en_0; // @[package.scala 94:16:@57863.4]
  assign RetimeWrapper_486_clock = clock; // @[:@57869.4]
  assign RetimeWrapper_486_reset = reset; // @[:@57870.4]
  assign RetimeWrapper_486_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57872.4]
  assign RetimeWrapper_486_io_in = _T_4777 & io_rPort_24_en_0; // @[package.scala 94:16:@57871.4]
  assign RetimeWrapper_487_clock = clock; // @[:@57877.4]
  assign RetimeWrapper_487_reset = reset; // @[:@57878.4]
  assign RetimeWrapper_487_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57880.4]
  assign RetimeWrapper_487_io_in = _T_5081 & io_rPort_24_en_0; // @[package.scala 94:16:@57879.4]
  assign RetimeWrapper_488_clock = clock; // @[:@57885.4]
  assign RetimeWrapper_488_reset = reset; // @[:@57886.4]
  assign RetimeWrapper_488_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57888.4]
  assign RetimeWrapper_488_io_in = _T_5385 & io_rPort_24_en_0; // @[package.scala 94:16:@57887.4]
  assign RetimeWrapper_489_clock = clock; // @[:@57893.4]
  assign RetimeWrapper_489_reset = reset; // @[:@57894.4]
  assign RetimeWrapper_489_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57896.4]
  assign RetimeWrapper_489_io_in = _T_5689 & io_rPort_24_en_0; // @[package.scala 94:16:@57895.4]
  assign RetimeWrapper_490_clock = clock; // @[:@57901.4]
  assign RetimeWrapper_490_reset = reset; // @[:@57902.4]
  assign RetimeWrapper_490_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57904.4]
  assign RetimeWrapper_490_io_in = _T_5993 & io_rPort_24_en_0; // @[package.scala 94:16:@57903.4]
  assign RetimeWrapper_491_clock = clock; // @[:@57909.4]
  assign RetimeWrapper_491_reset = reset; // @[:@57910.4]
  assign RetimeWrapper_491_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57912.4]
  assign RetimeWrapper_491_io_in = _T_6297 & io_rPort_24_en_0; // @[package.scala 94:16:@57911.4]
  assign RetimeWrapper_492_clock = clock; // @[:@57917.4]
  assign RetimeWrapper_492_reset = reset; // @[:@57918.4]
  assign RetimeWrapper_492_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57920.4]
  assign RetimeWrapper_492_io_in = _T_6601 & io_rPort_24_en_0; // @[package.scala 94:16:@57919.4]
  assign RetimeWrapper_493_clock = clock; // @[:@57925.4]
  assign RetimeWrapper_493_reset = reset; // @[:@57926.4]
  assign RetimeWrapper_493_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57928.4]
  assign RetimeWrapper_493_io_in = _T_6905 & io_rPort_24_en_0; // @[package.scala 94:16:@57927.4]
  assign RetimeWrapper_494_clock = clock; // @[:@57933.4]
  assign RetimeWrapper_494_reset = reset; // @[:@57934.4]
  assign RetimeWrapper_494_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57936.4]
  assign RetimeWrapper_494_io_in = _T_7209 & io_rPort_24_en_0; // @[package.scala 94:16:@57935.4]
  assign RetimeWrapper_495_clock = clock; // @[:@57941.4]
  assign RetimeWrapper_495_reset = reset; // @[:@57942.4]
  assign RetimeWrapper_495_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57944.4]
  assign RetimeWrapper_495_io_in = _T_7513 & io_rPort_24_en_0; // @[package.scala 94:16:@57943.4]
  assign RetimeWrapper_496_clock = clock; // @[:@57949.4]
  assign RetimeWrapper_496_reset = reset; // @[:@57950.4]
  assign RetimeWrapper_496_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57952.4]
  assign RetimeWrapper_496_io_in = _T_7817 & io_rPort_24_en_0; // @[package.scala 94:16:@57951.4]
  assign RetimeWrapper_497_clock = clock; // @[:@57957.4]
  assign RetimeWrapper_497_reset = reset; // @[:@57958.4]
  assign RetimeWrapper_497_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57960.4]
  assign RetimeWrapper_497_io_in = _T_8121 & io_rPort_24_en_0; // @[package.scala 94:16:@57959.4]
  assign RetimeWrapper_498_clock = clock; // @[:@57965.4]
  assign RetimeWrapper_498_reset = reset; // @[:@57966.4]
  assign RetimeWrapper_498_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57968.4]
  assign RetimeWrapper_498_io_in = _T_8425 & io_rPort_24_en_0; // @[package.scala 94:16:@57967.4]
  assign RetimeWrapper_499_clock = clock; // @[:@57973.4]
  assign RetimeWrapper_499_reset = reset; // @[:@57974.4]
  assign RetimeWrapper_499_io_flow = io_rPort_24_backpressure; // @[package.scala 95:18:@57976.4]
  assign RetimeWrapper_499_io_in = _T_8729 & io_rPort_24_en_0; // @[package.scala 94:16:@57975.4]
  assign RetimeWrapper_500_clock = clock; // @[:@58061.4]
  assign RetimeWrapper_500_reset = reset; // @[:@58062.4]
  assign RetimeWrapper_500_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58064.4]
  assign RetimeWrapper_500_io_in = _T_2959 & io_rPort_25_en_0; // @[package.scala 94:16:@58063.4]
  assign RetimeWrapper_501_clock = clock; // @[:@58069.4]
  assign RetimeWrapper_501_reset = reset; // @[:@58070.4]
  assign RetimeWrapper_501_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58072.4]
  assign RetimeWrapper_501_io_in = _T_3263 & io_rPort_25_en_0; // @[package.scala 94:16:@58071.4]
  assign RetimeWrapper_502_clock = clock; // @[:@58077.4]
  assign RetimeWrapper_502_reset = reset; // @[:@58078.4]
  assign RetimeWrapper_502_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58080.4]
  assign RetimeWrapper_502_io_in = _T_3567 & io_rPort_25_en_0; // @[package.scala 94:16:@58079.4]
  assign RetimeWrapper_503_clock = clock; // @[:@58085.4]
  assign RetimeWrapper_503_reset = reset; // @[:@58086.4]
  assign RetimeWrapper_503_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58088.4]
  assign RetimeWrapper_503_io_in = _T_3871 & io_rPort_25_en_0; // @[package.scala 94:16:@58087.4]
  assign RetimeWrapper_504_clock = clock; // @[:@58093.4]
  assign RetimeWrapper_504_reset = reset; // @[:@58094.4]
  assign RetimeWrapper_504_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58096.4]
  assign RetimeWrapper_504_io_in = _T_4175 & io_rPort_25_en_0; // @[package.scala 94:16:@58095.4]
  assign RetimeWrapper_505_clock = clock; // @[:@58101.4]
  assign RetimeWrapper_505_reset = reset; // @[:@58102.4]
  assign RetimeWrapper_505_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58104.4]
  assign RetimeWrapper_505_io_in = _T_4479 & io_rPort_25_en_0; // @[package.scala 94:16:@58103.4]
  assign RetimeWrapper_506_clock = clock; // @[:@58109.4]
  assign RetimeWrapper_506_reset = reset; // @[:@58110.4]
  assign RetimeWrapper_506_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58112.4]
  assign RetimeWrapper_506_io_in = _T_4783 & io_rPort_25_en_0; // @[package.scala 94:16:@58111.4]
  assign RetimeWrapper_507_clock = clock; // @[:@58117.4]
  assign RetimeWrapper_507_reset = reset; // @[:@58118.4]
  assign RetimeWrapper_507_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58120.4]
  assign RetimeWrapper_507_io_in = _T_5087 & io_rPort_25_en_0; // @[package.scala 94:16:@58119.4]
  assign RetimeWrapper_508_clock = clock; // @[:@58125.4]
  assign RetimeWrapper_508_reset = reset; // @[:@58126.4]
  assign RetimeWrapper_508_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58128.4]
  assign RetimeWrapper_508_io_in = _T_5391 & io_rPort_25_en_0; // @[package.scala 94:16:@58127.4]
  assign RetimeWrapper_509_clock = clock; // @[:@58133.4]
  assign RetimeWrapper_509_reset = reset; // @[:@58134.4]
  assign RetimeWrapper_509_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58136.4]
  assign RetimeWrapper_509_io_in = _T_5695 & io_rPort_25_en_0; // @[package.scala 94:16:@58135.4]
  assign RetimeWrapper_510_clock = clock; // @[:@58141.4]
  assign RetimeWrapper_510_reset = reset; // @[:@58142.4]
  assign RetimeWrapper_510_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58144.4]
  assign RetimeWrapper_510_io_in = _T_5999 & io_rPort_25_en_0; // @[package.scala 94:16:@58143.4]
  assign RetimeWrapper_511_clock = clock; // @[:@58149.4]
  assign RetimeWrapper_511_reset = reset; // @[:@58150.4]
  assign RetimeWrapper_511_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58152.4]
  assign RetimeWrapper_511_io_in = _T_6303 & io_rPort_25_en_0; // @[package.scala 94:16:@58151.4]
  assign RetimeWrapper_512_clock = clock; // @[:@58157.4]
  assign RetimeWrapper_512_reset = reset; // @[:@58158.4]
  assign RetimeWrapper_512_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58160.4]
  assign RetimeWrapper_512_io_in = _T_6607 & io_rPort_25_en_0; // @[package.scala 94:16:@58159.4]
  assign RetimeWrapper_513_clock = clock; // @[:@58165.4]
  assign RetimeWrapper_513_reset = reset; // @[:@58166.4]
  assign RetimeWrapper_513_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58168.4]
  assign RetimeWrapper_513_io_in = _T_6911 & io_rPort_25_en_0; // @[package.scala 94:16:@58167.4]
  assign RetimeWrapper_514_clock = clock; // @[:@58173.4]
  assign RetimeWrapper_514_reset = reset; // @[:@58174.4]
  assign RetimeWrapper_514_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58176.4]
  assign RetimeWrapper_514_io_in = _T_7215 & io_rPort_25_en_0; // @[package.scala 94:16:@58175.4]
  assign RetimeWrapper_515_clock = clock; // @[:@58181.4]
  assign RetimeWrapper_515_reset = reset; // @[:@58182.4]
  assign RetimeWrapper_515_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58184.4]
  assign RetimeWrapper_515_io_in = _T_7519 & io_rPort_25_en_0; // @[package.scala 94:16:@58183.4]
  assign RetimeWrapper_516_clock = clock; // @[:@58189.4]
  assign RetimeWrapper_516_reset = reset; // @[:@58190.4]
  assign RetimeWrapper_516_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58192.4]
  assign RetimeWrapper_516_io_in = _T_7823 & io_rPort_25_en_0; // @[package.scala 94:16:@58191.4]
  assign RetimeWrapper_517_clock = clock; // @[:@58197.4]
  assign RetimeWrapper_517_reset = reset; // @[:@58198.4]
  assign RetimeWrapper_517_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58200.4]
  assign RetimeWrapper_517_io_in = _T_8127 & io_rPort_25_en_0; // @[package.scala 94:16:@58199.4]
  assign RetimeWrapper_518_clock = clock; // @[:@58205.4]
  assign RetimeWrapper_518_reset = reset; // @[:@58206.4]
  assign RetimeWrapper_518_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58208.4]
  assign RetimeWrapper_518_io_in = _T_8431 & io_rPort_25_en_0; // @[package.scala 94:16:@58207.4]
  assign RetimeWrapper_519_clock = clock; // @[:@58213.4]
  assign RetimeWrapper_519_reset = reset; // @[:@58214.4]
  assign RetimeWrapper_519_io_flow = io_rPort_25_backpressure; // @[package.scala 95:18:@58216.4]
  assign RetimeWrapper_519_io_in = _T_8735 & io_rPort_25_en_0; // @[package.scala 94:16:@58215.4]
  assign RetimeWrapper_520_clock = clock; // @[:@58301.4]
  assign RetimeWrapper_520_reset = reset; // @[:@58302.4]
  assign RetimeWrapper_520_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58304.4]
  assign RetimeWrapper_520_io_in = _T_2813 & io_rPort_26_en_0; // @[package.scala 94:16:@58303.4]
  assign RetimeWrapper_521_clock = clock; // @[:@58309.4]
  assign RetimeWrapper_521_reset = reset; // @[:@58310.4]
  assign RetimeWrapper_521_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58312.4]
  assign RetimeWrapper_521_io_in = _T_3117 & io_rPort_26_en_0; // @[package.scala 94:16:@58311.4]
  assign RetimeWrapper_522_clock = clock; // @[:@58317.4]
  assign RetimeWrapper_522_reset = reset; // @[:@58318.4]
  assign RetimeWrapper_522_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58320.4]
  assign RetimeWrapper_522_io_in = _T_3421 & io_rPort_26_en_0; // @[package.scala 94:16:@58319.4]
  assign RetimeWrapper_523_clock = clock; // @[:@58325.4]
  assign RetimeWrapper_523_reset = reset; // @[:@58326.4]
  assign RetimeWrapper_523_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58328.4]
  assign RetimeWrapper_523_io_in = _T_3725 & io_rPort_26_en_0; // @[package.scala 94:16:@58327.4]
  assign RetimeWrapper_524_clock = clock; // @[:@58333.4]
  assign RetimeWrapper_524_reset = reset; // @[:@58334.4]
  assign RetimeWrapper_524_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58336.4]
  assign RetimeWrapper_524_io_in = _T_4029 & io_rPort_26_en_0; // @[package.scala 94:16:@58335.4]
  assign RetimeWrapper_525_clock = clock; // @[:@58341.4]
  assign RetimeWrapper_525_reset = reset; // @[:@58342.4]
  assign RetimeWrapper_525_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58344.4]
  assign RetimeWrapper_525_io_in = _T_4333 & io_rPort_26_en_0; // @[package.scala 94:16:@58343.4]
  assign RetimeWrapper_526_clock = clock; // @[:@58349.4]
  assign RetimeWrapper_526_reset = reset; // @[:@58350.4]
  assign RetimeWrapper_526_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58352.4]
  assign RetimeWrapper_526_io_in = _T_4637 & io_rPort_26_en_0; // @[package.scala 94:16:@58351.4]
  assign RetimeWrapper_527_clock = clock; // @[:@58357.4]
  assign RetimeWrapper_527_reset = reset; // @[:@58358.4]
  assign RetimeWrapper_527_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58360.4]
  assign RetimeWrapper_527_io_in = _T_4941 & io_rPort_26_en_0; // @[package.scala 94:16:@58359.4]
  assign RetimeWrapper_528_clock = clock; // @[:@58365.4]
  assign RetimeWrapper_528_reset = reset; // @[:@58366.4]
  assign RetimeWrapper_528_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58368.4]
  assign RetimeWrapper_528_io_in = _T_5245 & io_rPort_26_en_0; // @[package.scala 94:16:@58367.4]
  assign RetimeWrapper_529_clock = clock; // @[:@58373.4]
  assign RetimeWrapper_529_reset = reset; // @[:@58374.4]
  assign RetimeWrapper_529_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58376.4]
  assign RetimeWrapper_529_io_in = _T_5549 & io_rPort_26_en_0; // @[package.scala 94:16:@58375.4]
  assign RetimeWrapper_530_clock = clock; // @[:@58381.4]
  assign RetimeWrapper_530_reset = reset; // @[:@58382.4]
  assign RetimeWrapper_530_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58384.4]
  assign RetimeWrapper_530_io_in = _T_5853 & io_rPort_26_en_0; // @[package.scala 94:16:@58383.4]
  assign RetimeWrapper_531_clock = clock; // @[:@58389.4]
  assign RetimeWrapper_531_reset = reset; // @[:@58390.4]
  assign RetimeWrapper_531_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58392.4]
  assign RetimeWrapper_531_io_in = _T_6157 & io_rPort_26_en_0; // @[package.scala 94:16:@58391.4]
  assign RetimeWrapper_532_clock = clock; // @[:@58397.4]
  assign RetimeWrapper_532_reset = reset; // @[:@58398.4]
  assign RetimeWrapper_532_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58400.4]
  assign RetimeWrapper_532_io_in = _T_6461 & io_rPort_26_en_0; // @[package.scala 94:16:@58399.4]
  assign RetimeWrapper_533_clock = clock; // @[:@58405.4]
  assign RetimeWrapper_533_reset = reset; // @[:@58406.4]
  assign RetimeWrapper_533_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58408.4]
  assign RetimeWrapper_533_io_in = _T_6765 & io_rPort_26_en_0; // @[package.scala 94:16:@58407.4]
  assign RetimeWrapper_534_clock = clock; // @[:@58413.4]
  assign RetimeWrapper_534_reset = reset; // @[:@58414.4]
  assign RetimeWrapper_534_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58416.4]
  assign RetimeWrapper_534_io_in = _T_7069 & io_rPort_26_en_0; // @[package.scala 94:16:@58415.4]
  assign RetimeWrapper_535_clock = clock; // @[:@58421.4]
  assign RetimeWrapper_535_reset = reset; // @[:@58422.4]
  assign RetimeWrapper_535_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58424.4]
  assign RetimeWrapper_535_io_in = _T_7373 & io_rPort_26_en_0; // @[package.scala 94:16:@58423.4]
  assign RetimeWrapper_536_clock = clock; // @[:@58429.4]
  assign RetimeWrapper_536_reset = reset; // @[:@58430.4]
  assign RetimeWrapper_536_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58432.4]
  assign RetimeWrapper_536_io_in = _T_7677 & io_rPort_26_en_0; // @[package.scala 94:16:@58431.4]
  assign RetimeWrapper_537_clock = clock; // @[:@58437.4]
  assign RetimeWrapper_537_reset = reset; // @[:@58438.4]
  assign RetimeWrapper_537_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58440.4]
  assign RetimeWrapper_537_io_in = _T_7981 & io_rPort_26_en_0; // @[package.scala 94:16:@58439.4]
  assign RetimeWrapper_538_clock = clock; // @[:@58445.4]
  assign RetimeWrapper_538_reset = reset; // @[:@58446.4]
  assign RetimeWrapper_538_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58448.4]
  assign RetimeWrapper_538_io_in = _T_8285 & io_rPort_26_en_0; // @[package.scala 94:16:@58447.4]
  assign RetimeWrapper_539_clock = clock; // @[:@58453.4]
  assign RetimeWrapper_539_reset = reset; // @[:@58454.4]
  assign RetimeWrapper_539_io_flow = io_rPort_26_backpressure; // @[package.scala 95:18:@58456.4]
  assign RetimeWrapper_539_io_in = _T_8589 & io_rPort_26_en_0; // @[package.scala 94:16:@58455.4]
  assign RetimeWrapper_540_clock = clock; // @[:@58541.4]
  assign RetimeWrapper_540_reset = reset; // @[:@58542.4]
  assign RetimeWrapper_540_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58544.4]
  assign RetimeWrapper_540_io_in = _T_2965 & io_rPort_27_en_0; // @[package.scala 94:16:@58543.4]
  assign RetimeWrapper_541_clock = clock; // @[:@58549.4]
  assign RetimeWrapper_541_reset = reset; // @[:@58550.4]
  assign RetimeWrapper_541_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58552.4]
  assign RetimeWrapper_541_io_in = _T_3269 & io_rPort_27_en_0; // @[package.scala 94:16:@58551.4]
  assign RetimeWrapper_542_clock = clock; // @[:@58557.4]
  assign RetimeWrapper_542_reset = reset; // @[:@58558.4]
  assign RetimeWrapper_542_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58560.4]
  assign RetimeWrapper_542_io_in = _T_3573 & io_rPort_27_en_0; // @[package.scala 94:16:@58559.4]
  assign RetimeWrapper_543_clock = clock; // @[:@58565.4]
  assign RetimeWrapper_543_reset = reset; // @[:@58566.4]
  assign RetimeWrapper_543_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58568.4]
  assign RetimeWrapper_543_io_in = _T_3877 & io_rPort_27_en_0; // @[package.scala 94:16:@58567.4]
  assign RetimeWrapper_544_clock = clock; // @[:@58573.4]
  assign RetimeWrapper_544_reset = reset; // @[:@58574.4]
  assign RetimeWrapper_544_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58576.4]
  assign RetimeWrapper_544_io_in = _T_4181 & io_rPort_27_en_0; // @[package.scala 94:16:@58575.4]
  assign RetimeWrapper_545_clock = clock; // @[:@58581.4]
  assign RetimeWrapper_545_reset = reset; // @[:@58582.4]
  assign RetimeWrapper_545_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58584.4]
  assign RetimeWrapper_545_io_in = _T_4485 & io_rPort_27_en_0; // @[package.scala 94:16:@58583.4]
  assign RetimeWrapper_546_clock = clock; // @[:@58589.4]
  assign RetimeWrapper_546_reset = reset; // @[:@58590.4]
  assign RetimeWrapper_546_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58592.4]
  assign RetimeWrapper_546_io_in = _T_4789 & io_rPort_27_en_0; // @[package.scala 94:16:@58591.4]
  assign RetimeWrapper_547_clock = clock; // @[:@58597.4]
  assign RetimeWrapper_547_reset = reset; // @[:@58598.4]
  assign RetimeWrapper_547_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58600.4]
  assign RetimeWrapper_547_io_in = _T_5093 & io_rPort_27_en_0; // @[package.scala 94:16:@58599.4]
  assign RetimeWrapper_548_clock = clock; // @[:@58605.4]
  assign RetimeWrapper_548_reset = reset; // @[:@58606.4]
  assign RetimeWrapper_548_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58608.4]
  assign RetimeWrapper_548_io_in = _T_5397 & io_rPort_27_en_0; // @[package.scala 94:16:@58607.4]
  assign RetimeWrapper_549_clock = clock; // @[:@58613.4]
  assign RetimeWrapper_549_reset = reset; // @[:@58614.4]
  assign RetimeWrapper_549_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58616.4]
  assign RetimeWrapper_549_io_in = _T_5701 & io_rPort_27_en_0; // @[package.scala 94:16:@58615.4]
  assign RetimeWrapper_550_clock = clock; // @[:@58621.4]
  assign RetimeWrapper_550_reset = reset; // @[:@58622.4]
  assign RetimeWrapper_550_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58624.4]
  assign RetimeWrapper_550_io_in = _T_6005 & io_rPort_27_en_0; // @[package.scala 94:16:@58623.4]
  assign RetimeWrapper_551_clock = clock; // @[:@58629.4]
  assign RetimeWrapper_551_reset = reset; // @[:@58630.4]
  assign RetimeWrapper_551_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58632.4]
  assign RetimeWrapper_551_io_in = _T_6309 & io_rPort_27_en_0; // @[package.scala 94:16:@58631.4]
  assign RetimeWrapper_552_clock = clock; // @[:@58637.4]
  assign RetimeWrapper_552_reset = reset; // @[:@58638.4]
  assign RetimeWrapper_552_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58640.4]
  assign RetimeWrapper_552_io_in = _T_6613 & io_rPort_27_en_0; // @[package.scala 94:16:@58639.4]
  assign RetimeWrapper_553_clock = clock; // @[:@58645.4]
  assign RetimeWrapper_553_reset = reset; // @[:@58646.4]
  assign RetimeWrapper_553_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58648.4]
  assign RetimeWrapper_553_io_in = _T_6917 & io_rPort_27_en_0; // @[package.scala 94:16:@58647.4]
  assign RetimeWrapper_554_clock = clock; // @[:@58653.4]
  assign RetimeWrapper_554_reset = reset; // @[:@58654.4]
  assign RetimeWrapper_554_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58656.4]
  assign RetimeWrapper_554_io_in = _T_7221 & io_rPort_27_en_0; // @[package.scala 94:16:@58655.4]
  assign RetimeWrapper_555_clock = clock; // @[:@58661.4]
  assign RetimeWrapper_555_reset = reset; // @[:@58662.4]
  assign RetimeWrapper_555_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58664.4]
  assign RetimeWrapper_555_io_in = _T_7525 & io_rPort_27_en_0; // @[package.scala 94:16:@58663.4]
  assign RetimeWrapper_556_clock = clock; // @[:@58669.4]
  assign RetimeWrapper_556_reset = reset; // @[:@58670.4]
  assign RetimeWrapper_556_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58672.4]
  assign RetimeWrapper_556_io_in = _T_7829 & io_rPort_27_en_0; // @[package.scala 94:16:@58671.4]
  assign RetimeWrapper_557_clock = clock; // @[:@58677.4]
  assign RetimeWrapper_557_reset = reset; // @[:@58678.4]
  assign RetimeWrapper_557_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58680.4]
  assign RetimeWrapper_557_io_in = _T_8133 & io_rPort_27_en_0; // @[package.scala 94:16:@58679.4]
  assign RetimeWrapper_558_clock = clock; // @[:@58685.4]
  assign RetimeWrapper_558_reset = reset; // @[:@58686.4]
  assign RetimeWrapper_558_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58688.4]
  assign RetimeWrapper_558_io_in = _T_8437 & io_rPort_27_en_0; // @[package.scala 94:16:@58687.4]
  assign RetimeWrapper_559_clock = clock; // @[:@58693.4]
  assign RetimeWrapper_559_reset = reset; // @[:@58694.4]
  assign RetimeWrapper_559_io_flow = io_rPort_27_backpressure; // @[package.scala 95:18:@58696.4]
  assign RetimeWrapper_559_io_in = _T_8741 & io_rPort_27_en_0; // @[package.scala 94:16:@58695.4]
  assign RetimeWrapper_560_clock = clock; // @[:@58781.4]
  assign RetimeWrapper_560_reset = reset; // @[:@58782.4]
  assign RetimeWrapper_560_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58784.4]
  assign RetimeWrapper_560_io_in = _T_2971 & io_rPort_28_en_0; // @[package.scala 94:16:@58783.4]
  assign RetimeWrapper_561_clock = clock; // @[:@58789.4]
  assign RetimeWrapper_561_reset = reset; // @[:@58790.4]
  assign RetimeWrapper_561_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58792.4]
  assign RetimeWrapper_561_io_in = _T_3275 & io_rPort_28_en_0; // @[package.scala 94:16:@58791.4]
  assign RetimeWrapper_562_clock = clock; // @[:@58797.4]
  assign RetimeWrapper_562_reset = reset; // @[:@58798.4]
  assign RetimeWrapper_562_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58800.4]
  assign RetimeWrapper_562_io_in = _T_3579 & io_rPort_28_en_0; // @[package.scala 94:16:@58799.4]
  assign RetimeWrapper_563_clock = clock; // @[:@58805.4]
  assign RetimeWrapper_563_reset = reset; // @[:@58806.4]
  assign RetimeWrapper_563_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58808.4]
  assign RetimeWrapper_563_io_in = _T_3883 & io_rPort_28_en_0; // @[package.scala 94:16:@58807.4]
  assign RetimeWrapper_564_clock = clock; // @[:@58813.4]
  assign RetimeWrapper_564_reset = reset; // @[:@58814.4]
  assign RetimeWrapper_564_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58816.4]
  assign RetimeWrapper_564_io_in = _T_4187 & io_rPort_28_en_0; // @[package.scala 94:16:@58815.4]
  assign RetimeWrapper_565_clock = clock; // @[:@58821.4]
  assign RetimeWrapper_565_reset = reset; // @[:@58822.4]
  assign RetimeWrapper_565_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58824.4]
  assign RetimeWrapper_565_io_in = _T_4491 & io_rPort_28_en_0; // @[package.scala 94:16:@58823.4]
  assign RetimeWrapper_566_clock = clock; // @[:@58829.4]
  assign RetimeWrapper_566_reset = reset; // @[:@58830.4]
  assign RetimeWrapper_566_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58832.4]
  assign RetimeWrapper_566_io_in = _T_4795 & io_rPort_28_en_0; // @[package.scala 94:16:@58831.4]
  assign RetimeWrapper_567_clock = clock; // @[:@58837.4]
  assign RetimeWrapper_567_reset = reset; // @[:@58838.4]
  assign RetimeWrapper_567_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58840.4]
  assign RetimeWrapper_567_io_in = _T_5099 & io_rPort_28_en_0; // @[package.scala 94:16:@58839.4]
  assign RetimeWrapper_568_clock = clock; // @[:@58845.4]
  assign RetimeWrapper_568_reset = reset; // @[:@58846.4]
  assign RetimeWrapper_568_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58848.4]
  assign RetimeWrapper_568_io_in = _T_5403 & io_rPort_28_en_0; // @[package.scala 94:16:@58847.4]
  assign RetimeWrapper_569_clock = clock; // @[:@58853.4]
  assign RetimeWrapper_569_reset = reset; // @[:@58854.4]
  assign RetimeWrapper_569_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58856.4]
  assign RetimeWrapper_569_io_in = _T_5707 & io_rPort_28_en_0; // @[package.scala 94:16:@58855.4]
  assign RetimeWrapper_570_clock = clock; // @[:@58861.4]
  assign RetimeWrapper_570_reset = reset; // @[:@58862.4]
  assign RetimeWrapper_570_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58864.4]
  assign RetimeWrapper_570_io_in = _T_6011 & io_rPort_28_en_0; // @[package.scala 94:16:@58863.4]
  assign RetimeWrapper_571_clock = clock; // @[:@58869.4]
  assign RetimeWrapper_571_reset = reset; // @[:@58870.4]
  assign RetimeWrapper_571_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58872.4]
  assign RetimeWrapper_571_io_in = _T_6315 & io_rPort_28_en_0; // @[package.scala 94:16:@58871.4]
  assign RetimeWrapper_572_clock = clock; // @[:@58877.4]
  assign RetimeWrapper_572_reset = reset; // @[:@58878.4]
  assign RetimeWrapper_572_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58880.4]
  assign RetimeWrapper_572_io_in = _T_6619 & io_rPort_28_en_0; // @[package.scala 94:16:@58879.4]
  assign RetimeWrapper_573_clock = clock; // @[:@58885.4]
  assign RetimeWrapper_573_reset = reset; // @[:@58886.4]
  assign RetimeWrapper_573_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58888.4]
  assign RetimeWrapper_573_io_in = _T_6923 & io_rPort_28_en_0; // @[package.scala 94:16:@58887.4]
  assign RetimeWrapper_574_clock = clock; // @[:@58893.4]
  assign RetimeWrapper_574_reset = reset; // @[:@58894.4]
  assign RetimeWrapper_574_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58896.4]
  assign RetimeWrapper_574_io_in = _T_7227 & io_rPort_28_en_0; // @[package.scala 94:16:@58895.4]
  assign RetimeWrapper_575_clock = clock; // @[:@58901.4]
  assign RetimeWrapper_575_reset = reset; // @[:@58902.4]
  assign RetimeWrapper_575_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58904.4]
  assign RetimeWrapper_575_io_in = _T_7531 & io_rPort_28_en_0; // @[package.scala 94:16:@58903.4]
  assign RetimeWrapper_576_clock = clock; // @[:@58909.4]
  assign RetimeWrapper_576_reset = reset; // @[:@58910.4]
  assign RetimeWrapper_576_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58912.4]
  assign RetimeWrapper_576_io_in = _T_7835 & io_rPort_28_en_0; // @[package.scala 94:16:@58911.4]
  assign RetimeWrapper_577_clock = clock; // @[:@58917.4]
  assign RetimeWrapper_577_reset = reset; // @[:@58918.4]
  assign RetimeWrapper_577_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58920.4]
  assign RetimeWrapper_577_io_in = _T_8139 & io_rPort_28_en_0; // @[package.scala 94:16:@58919.4]
  assign RetimeWrapper_578_clock = clock; // @[:@58925.4]
  assign RetimeWrapper_578_reset = reset; // @[:@58926.4]
  assign RetimeWrapper_578_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58928.4]
  assign RetimeWrapper_578_io_in = _T_8443 & io_rPort_28_en_0; // @[package.scala 94:16:@58927.4]
  assign RetimeWrapper_579_clock = clock; // @[:@58933.4]
  assign RetimeWrapper_579_reset = reset; // @[:@58934.4]
  assign RetimeWrapper_579_io_flow = io_rPort_28_backpressure; // @[package.scala 95:18:@58936.4]
  assign RetimeWrapper_579_io_in = _T_8747 & io_rPort_28_en_0; // @[package.scala 94:16:@58935.4]
  assign RetimeWrapper_580_clock = clock; // @[:@59021.4]
  assign RetimeWrapper_580_reset = reset; // @[:@59022.4]
  assign RetimeWrapper_580_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59024.4]
  assign RetimeWrapper_580_io_in = _T_2819 & io_rPort_29_en_0; // @[package.scala 94:16:@59023.4]
  assign RetimeWrapper_581_clock = clock; // @[:@59029.4]
  assign RetimeWrapper_581_reset = reset; // @[:@59030.4]
  assign RetimeWrapper_581_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59032.4]
  assign RetimeWrapper_581_io_in = _T_3123 & io_rPort_29_en_0; // @[package.scala 94:16:@59031.4]
  assign RetimeWrapper_582_clock = clock; // @[:@59037.4]
  assign RetimeWrapper_582_reset = reset; // @[:@59038.4]
  assign RetimeWrapper_582_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59040.4]
  assign RetimeWrapper_582_io_in = _T_3427 & io_rPort_29_en_0; // @[package.scala 94:16:@59039.4]
  assign RetimeWrapper_583_clock = clock; // @[:@59045.4]
  assign RetimeWrapper_583_reset = reset; // @[:@59046.4]
  assign RetimeWrapper_583_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59048.4]
  assign RetimeWrapper_583_io_in = _T_3731 & io_rPort_29_en_0; // @[package.scala 94:16:@59047.4]
  assign RetimeWrapper_584_clock = clock; // @[:@59053.4]
  assign RetimeWrapper_584_reset = reset; // @[:@59054.4]
  assign RetimeWrapper_584_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59056.4]
  assign RetimeWrapper_584_io_in = _T_4035 & io_rPort_29_en_0; // @[package.scala 94:16:@59055.4]
  assign RetimeWrapper_585_clock = clock; // @[:@59061.4]
  assign RetimeWrapper_585_reset = reset; // @[:@59062.4]
  assign RetimeWrapper_585_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59064.4]
  assign RetimeWrapper_585_io_in = _T_4339 & io_rPort_29_en_0; // @[package.scala 94:16:@59063.4]
  assign RetimeWrapper_586_clock = clock; // @[:@59069.4]
  assign RetimeWrapper_586_reset = reset; // @[:@59070.4]
  assign RetimeWrapper_586_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59072.4]
  assign RetimeWrapper_586_io_in = _T_4643 & io_rPort_29_en_0; // @[package.scala 94:16:@59071.4]
  assign RetimeWrapper_587_clock = clock; // @[:@59077.4]
  assign RetimeWrapper_587_reset = reset; // @[:@59078.4]
  assign RetimeWrapper_587_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59080.4]
  assign RetimeWrapper_587_io_in = _T_4947 & io_rPort_29_en_0; // @[package.scala 94:16:@59079.4]
  assign RetimeWrapper_588_clock = clock; // @[:@59085.4]
  assign RetimeWrapper_588_reset = reset; // @[:@59086.4]
  assign RetimeWrapper_588_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59088.4]
  assign RetimeWrapper_588_io_in = _T_5251 & io_rPort_29_en_0; // @[package.scala 94:16:@59087.4]
  assign RetimeWrapper_589_clock = clock; // @[:@59093.4]
  assign RetimeWrapper_589_reset = reset; // @[:@59094.4]
  assign RetimeWrapper_589_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59096.4]
  assign RetimeWrapper_589_io_in = _T_5555 & io_rPort_29_en_0; // @[package.scala 94:16:@59095.4]
  assign RetimeWrapper_590_clock = clock; // @[:@59101.4]
  assign RetimeWrapper_590_reset = reset; // @[:@59102.4]
  assign RetimeWrapper_590_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59104.4]
  assign RetimeWrapper_590_io_in = _T_5859 & io_rPort_29_en_0; // @[package.scala 94:16:@59103.4]
  assign RetimeWrapper_591_clock = clock; // @[:@59109.4]
  assign RetimeWrapper_591_reset = reset; // @[:@59110.4]
  assign RetimeWrapper_591_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59112.4]
  assign RetimeWrapper_591_io_in = _T_6163 & io_rPort_29_en_0; // @[package.scala 94:16:@59111.4]
  assign RetimeWrapper_592_clock = clock; // @[:@59117.4]
  assign RetimeWrapper_592_reset = reset; // @[:@59118.4]
  assign RetimeWrapper_592_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59120.4]
  assign RetimeWrapper_592_io_in = _T_6467 & io_rPort_29_en_0; // @[package.scala 94:16:@59119.4]
  assign RetimeWrapper_593_clock = clock; // @[:@59125.4]
  assign RetimeWrapper_593_reset = reset; // @[:@59126.4]
  assign RetimeWrapper_593_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59128.4]
  assign RetimeWrapper_593_io_in = _T_6771 & io_rPort_29_en_0; // @[package.scala 94:16:@59127.4]
  assign RetimeWrapper_594_clock = clock; // @[:@59133.4]
  assign RetimeWrapper_594_reset = reset; // @[:@59134.4]
  assign RetimeWrapper_594_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59136.4]
  assign RetimeWrapper_594_io_in = _T_7075 & io_rPort_29_en_0; // @[package.scala 94:16:@59135.4]
  assign RetimeWrapper_595_clock = clock; // @[:@59141.4]
  assign RetimeWrapper_595_reset = reset; // @[:@59142.4]
  assign RetimeWrapper_595_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59144.4]
  assign RetimeWrapper_595_io_in = _T_7379 & io_rPort_29_en_0; // @[package.scala 94:16:@59143.4]
  assign RetimeWrapper_596_clock = clock; // @[:@59149.4]
  assign RetimeWrapper_596_reset = reset; // @[:@59150.4]
  assign RetimeWrapper_596_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59152.4]
  assign RetimeWrapper_596_io_in = _T_7683 & io_rPort_29_en_0; // @[package.scala 94:16:@59151.4]
  assign RetimeWrapper_597_clock = clock; // @[:@59157.4]
  assign RetimeWrapper_597_reset = reset; // @[:@59158.4]
  assign RetimeWrapper_597_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59160.4]
  assign RetimeWrapper_597_io_in = _T_7987 & io_rPort_29_en_0; // @[package.scala 94:16:@59159.4]
  assign RetimeWrapper_598_clock = clock; // @[:@59165.4]
  assign RetimeWrapper_598_reset = reset; // @[:@59166.4]
  assign RetimeWrapper_598_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59168.4]
  assign RetimeWrapper_598_io_in = _T_8291 & io_rPort_29_en_0; // @[package.scala 94:16:@59167.4]
  assign RetimeWrapper_599_clock = clock; // @[:@59173.4]
  assign RetimeWrapper_599_reset = reset; // @[:@59174.4]
  assign RetimeWrapper_599_io_flow = io_rPort_29_backpressure; // @[package.scala 95:18:@59176.4]
  assign RetimeWrapper_599_io_in = _T_8595 & io_rPort_29_en_0; // @[package.scala 94:16:@59175.4]
endmodule
module RetimeWrapper_705( // @[:@59212.2]
  input         clock, // @[:@59213.4]
  input         reset, // @[:@59214.4]
  input         io_flow, // @[:@59215.4]
  input  [31:0] io_in, // @[:@59215.4]
  output [31:0] io_out // @[:@59215.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59217.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59217.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59217.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59217.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59217.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59217.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@59217.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59230.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59229.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@59228.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59227.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59226.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59224.4]
endmodule
module RetimeWrapper_706( // @[:@59244.2]
  input         clock, // @[:@59245.4]
  input         reset, // @[:@59246.4]
  input         io_flow, // @[:@59247.4]
  input  [31:0] io_in, // @[:@59247.4]
  output [31:0] io_out // @[:@59247.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59249.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59249.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59249.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59249.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59249.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59249.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@59249.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59262.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59261.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@59260.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59259.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59258.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59256.4]
endmodule
module fix2fixBox_18( // @[:@59264.2]
  input  [63:0] io_a, // @[:@59267.4]
  output [31:0] io_b // @[:@59267.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@59280.4]
endmodule
module x814( // @[:@59282.2]
  input         clock, // @[:@59283.4]
  input         reset, // @[:@59284.4]
  input  [31:0] io_a, // @[:@59285.4]
  input         io_flow, // @[:@59285.4]
  output [31:0] io_result // @[:@59285.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@59294.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@59294.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@59294.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@59294.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@59294.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@59302.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@59302.4]
  wire [31:0] _T_19; // @[package.scala 96:25:@59299.4 package.scala 96:25:@59300.4]
  wire [31:0] _GEN_0; // @[package.scala 94:16:@59297.4]
  RetimeWrapper_706 RetimeWrapper ( // @[package.scala 93:22:@59294.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  fix2fixBox_18 fix2fixBox ( // @[Math.scala 357:30:@59302.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_19 = RetimeWrapper_io_out; // @[package.scala 96:25:@59299.4 package.scala 96:25:@59300.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@59310.4]
  assign RetimeWrapper_clock = clock; // @[:@59295.4]
  assign RetimeWrapper_reset = reset; // @[:@59296.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@59298.4]
  assign _GEN_0 = io_a % 32'ha; // @[package.scala 94:16:@59297.4]
  assign RetimeWrapper_io_in = _GEN_0[31:0]; // @[package.scala 94:16:@59297.4]
  assign fix2fixBox_io_a = {{32'd0}, _T_19}; // @[Math.scala 358:23:@59305.4]
endmodule
module RetimeWrapper_708( // @[:@59513.2]
  input         clock, // @[:@59514.4]
  input         reset, // @[:@59515.4]
  input         io_flow, // @[:@59516.4]
  input  [31:0] io_in, // @[:@59516.4]
  output [31:0] io_out // @[:@59516.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59518.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59518.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59518.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59518.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59518.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59518.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@59518.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59531.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59530.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@59529.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59528.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59527.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59525.4]
endmodule
module x817_div( // @[:@59574.2]
  input         clock, // @[:@59575.4]
  input         reset, // @[:@59576.4]
  input  [31:0] io_a, // @[:@59577.4]
  input         io_flow, // @[:@59577.4]
  output [31:0] io_result // @[:@59577.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@59586.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@59586.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@59586.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@59586.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@59586.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@59599.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@59599.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@59583.4]
  wire [32:0] _T_17; // @[BigIPSim.scala 23:39:@59585.4]
  wire [32:0] _T_18; // @[package.scala 94:23:@59589.4]
  wire [31:0] _T_21; // @[package.scala 96:25:@59593.4]
  RetimeWrapper_708 RetimeWrapper ( // @[package.scala 93:22:@59586.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ _ ( // @[Math.scala 709:24:@59599.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@59583.4]
  assign _T_17 = $signed(_T_15) / $signed(32'sha); // @[BigIPSim.scala 23:39:@59585.4]
  assign _T_18 = $unsigned(_T_17); // @[package.scala 94:23:@59589.4]
  assign _T_21 = $signed(RetimeWrapper_io_out); // @[package.scala 96:25:@59593.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@59607.4]
  assign RetimeWrapper_clock = clock; // @[:@59587.4]
  assign RetimeWrapper_reset = reset; // @[:@59588.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@59591.4]
  assign RetimeWrapper_io_in = _T_18[31:0]; // @[package.scala 94:16:@59590.4]
  assign __io_b = $unsigned(_T_21); // @[Math.scala 710:17:@59602.4]
endmodule
module RetimeWrapper_709( // @[:@59621.2]
  input         clock, // @[:@59622.4]
  input         reset, // @[:@59623.4]
  input         io_flow, // @[:@59624.4]
  input  [31:0] io_in, // @[:@59624.4]
  output [31:0] io_out // @[:@59624.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59626.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59626.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59626.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59626.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59626.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59626.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@59626.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59639.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59638.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@59637.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59636.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59635.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59633.4]
endmodule
module RetimeWrapper_711( // @[:@59842.2]
  input         clock, // @[:@59843.4]
  input         reset, // @[:@59844.4]
  input         io_flow, // @[:@59845.4]
  input  [31:0] io_in, // @[:@59845.4]
  output [31:0] io_out // @[:@59845.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59847.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59847.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59847.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59847.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59847.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59847.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@59847.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59860.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59859.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@59858.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59857.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59856.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59854.4]
endmodule
module RetimeWrapper_712( // @[:@59874.2]
  input   clock, // @[:@59875.4]
  input   reset, // @[:@59876.4]
  input   io_flow, // @[:@59877.4]
  input   io_in, // @[:@59877.4]
  output  io_out // @[:@59877.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@59879.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@59879.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@59879.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59879.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59879.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59879.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(28)) sr ( // @[RetimeShiftRegister.scala 15:20:@59879.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59892.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59891.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@59890.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59889.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59888.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59886.4]
endmodule
module RetimeWrapper_713( // @[:@59906.2]
  input         clock, // @[:@59907.4]
  input         reset, // @[:@59908.4]
  input         io_flow, // @[:@59909.4]
  input  [31:0] io_in, // @[:@59909.4]
  output [31:0] io_out // @[:@59909.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59911.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59911.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59911.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59911.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59911.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59911.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@59911.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59924.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59923.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@59922.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59921.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59920.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59918.4]
endmodule
module RetimeWrapper_714( // @[:@59938.2]
  input        clock, // @[:@59939.4]
  input        reset, // @[:@59940.4]
  input        io_flow, // @[:@59941.4]
  input  [7:0] io_in, // @[:@59941.4]
  output [7:0] io_out // @[:@59941.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59943.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59943.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59943.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59943.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59943.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59943.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@59943.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59956.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59955.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@59954.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59953.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59952.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59950.4]
endmodule
module RetimeWrapper_715( // @[:@59970.2]
  input         clock, // @[:@59971.4]
  input         reset, // @[:@59972.4]
  input         io_flow, // @[:@59973.4]
  input  [31:0] io_in, // @[:@59973.4]
  output [31:0] io_out // @[:@59973.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59975.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59975.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59975.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59975.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59975.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59975.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@59975.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59988.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59987.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@59986.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59985.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59984.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59982.4]
endmodule
module RetimeWrapper_721( // @[:@60443.2]
  input         clock, // @[:@60444.4]
  input         reset, // @[:@60445.4]
  input         io_flow, // @[:@60446.4]
  input  [31:0] io_in, // @[:@60446.4]
  output [31:0] io_out // @[:@60446.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@60448.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@60448.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@60448.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@60448.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@60448.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@60448.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@60448.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@60461.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@60460.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@60459.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@60458.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@60457.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@60455.4]
endmodule
module RetimeWrapper_724( // @[:@60696.2]
  input         clock, // @[:@60697.4]
  input         reset, // @[:@60698.4]
  input         io_flow, // @[:@60699.4]
  input  [31:0] io_in, // @[:@60699.4]
  output [31:0] io_out // @[:@60699.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@60701.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@60701.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@60701.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@60701.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@60701.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@60701.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@60701.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@60714.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@60713.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@60712.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@60711.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@60710.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@60708.4]
endmodule
module RetimeWrapper_725( // @[:@60728.2]
  input         clock, // @[:@60729.4]
  input         reset, // @[:@60730.4]
  input         io_flow, // @[:@60731.4]
  input  [31:0] io_in, // @[:@60731.4]
  output [31:0] io_out // @[:@60731.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@60733.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@60733.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@60733.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@60733.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@60733.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@60733.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@60733.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@60746.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@60745.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@60744.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@60743.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@60742.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@60740.4]
endmodule
module RetimeWrapper_775( // @[:@64956.2]
  input         clock, // @[:@64957.4]
  input         reset, // @[:@64958.4]
  input         io_flow, // @[:@64959.4]
  input  [31:0] io_in, // @[:@64959.4]
  output [31:0] io_out // @[:@64959.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@64961.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@64961.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@64961.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@64961.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@64961.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@64961.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(30)) sr ( // @[RetimeShiftRegister.scala 15:20:@64961.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@64974.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@64973.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@64972.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@64971.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@64970.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@64968.4]
endmodule
module RetimeWrapper_782( // @[:@65337.2]
  input         clock, // @[:@65338.4]
  input         reset, // @[:@65339.4]
  input         io_flow, // @[:@65340.4]
  input  [31:0] io_in, // @[:@65340.4]
  output [31:0] io_out // @[:@65340.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@65342.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@65342.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@65342.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@65342.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@65342.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@65342.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@65342.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@65355.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@65354.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@65353.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@65352.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@65351.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@65349.4]
endmodule
module RetimeWrapper_785( // @[:@65590.2]
  input         clock, // @[:@65591.4]
  input         reset, // @[:@65592.4]
  input         io_flow, // @[:@65593.4]
  input  [31:0] io_in, // @[:@65593.4]
  output [31:0] io_out // @[:@65593.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@65595.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@65595.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@65595.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@65595.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@65595.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@65595.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@65595.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@65608.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@65607.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@65606.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@65605.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@65604.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@65602.4]
endmodule
module RetimeWrapper_786( // @[:@65622.2]
  input   clock, // @[:@65623.4]
  input   reset, // @[:@65624.4]
  input   io_flow, // @[:@65625.4]
  input   io_in, // @[:@65625.4]
  output  io_out // @[:@65625.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@65627.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@65627.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@65627.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@65627.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@65627.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@65627.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(52)) sr ( // @[RetimeShiftRegister.scala 15:20:@65627.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@65640.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@65639.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@65638.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@65637.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@65636.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@65634.4]
endmodule
module RetimeWrapper_787( // @[:@65654.2]
  input         clock, // @[:@65655.4]
  input         reset, // @[:@65656.4]
  input         io_flow, // @[:@65657.4]
  input  [31:0] io_in, // @[:@65657.4]
  output [31:0] io_out // @[:@65657.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@65659.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@65659.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@65659.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@65659.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@65659.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@65659.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(35)) sr ( // @[RetimeShiftRegister.scala 15:20:@65659.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@65672.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@65671.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@65670.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@65669.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@65668.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@65666.4]
endmodule
module RetimeWrapper_788( // @[:@65686.2]
  input   clock, // @[:@65687.4]
  input   reset, // @[:@65688.4]
  input   io_flow, // @[:@65689.4]
  input   io_in, // @[:@65689.4]
  output  io_out // @[:@65689.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@65691.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@65691.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@65691.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@65691.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@65691.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@65691.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@65691.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@65704.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@65703.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@65702.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@65701.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@65700.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@65698.4]
endmodule
module RetimeWrapper_838( // @[:@68385.2]
  input         clock, // @[:@68386.4]
  input         reset, // @[:@68387.4]
  input         io_flow, // @[:@68388.4]
  input  [31:0] io_in, // @[:@68388.4]
  output [31:0] io_out // @[:@68388.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@68390.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@68390.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@68390.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@68390.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@68390.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@68390.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(36)) sr ( // @[RetimeShiftRegister.scala 15:20:@68390.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@68403.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@68402.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@68401.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@68400.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@68399.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@68397.4]
endmodule
module RetimeWrapper_840( // @[:@68449.2]
  input   clock, // @[:@68450.4]
  input   reset, // @[:@68451.4]
  input   io_flow, // @[:@68452.4]
  input   io_in, // @[:@68452.4]
  output  io_out // @[:@68452.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@68454.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@68454.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@68454.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@68454.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@68454.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@68454.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@68454.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@68467.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@68466.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@68465.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@68464.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@68463.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@68461.4]
endmodule
module RetimeWrapper_847( // @[:@69111.2]
  input         clock, // @[:@69112.4]
  input         reset, // @[:@69113.4]
  input         io_flow, // @[:@69114.4]
  input  [31:0] io_in, // @[:@69114.4]
  output [31:0] io_out // @[:@69114.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@69116.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@69116.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@69116.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@69116.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@69116.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@69116.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@69116.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@69129.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@69128.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@69127.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@69126.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@69125.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@69123.4]
endmodule
module RetimeWrapper_935( // @[:@76135.2]
  input        clock, // @[:@76136.4]
  input        reset, // @[:@76137.4]
  input        io_flow, // @[:@76138.4]
  input  [8:0] io_in, // @[:@76138.4]
  output [8:0] io_out // @[:@76138.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@76140.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@76140.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@76140.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@76140.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@76140.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@76140.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@76140.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@76153.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@76152.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@76151.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@76150.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@76149.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@76147.4]
endmodule
module RetimeWrapper_937( // @[:@76199.2]
  input        clock, // @[:@76200.4]
  input        reset, // @[:@76201.4]
  input        io_flow, // @[:@76202.4]
  input  [9:0] io_in, // @[:@76202.4]
  output [9:0] io_out // @[:@76202.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@76204.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@76204.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@76204.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@76204.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@76204.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@76204.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@76204.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@76217.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@76216.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@76215.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@76214.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@76213.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@76211.4]
endmodule
module SimBlackBoxesfix2fixBox_164( // @[:@76315.2]
  input  [7:0] io_a, // @[:@76318.4]
  output [8:0] io_b // @[:@76318.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@76332.4]
endmodule
module __156( // @[:@76334.2]
  input  [7:0] io_b, // @[:@76337.4]
  output [8:0] io_result // @[:@76337.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@76342.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@76342.4]
  SimBlackBoxesfix2fixBox_164 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@76342.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@76355.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@76350.4]
endmodule
module fix2fixBox_81( // @[:@76399.2]
  input  [8:0] io_a, // @[:@76402.4]
  output [7:0] io_b // @[:@76402.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@76415.4]
endmodule
module x1051_x15( // @[:@76417.2]
  input  [7:0] io_a, // @[:@76420.4]
  input  [7:0] io_b, // @[:@76420.4]
  output [7:0] io_result // @[:@76420.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@76428.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@76428.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@76435.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@76435.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@76445.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@76445.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@76433.4 Math.scala 713:14:@76434.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@76440.4 Math.scala 713:14:@76441.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@76442.4]
  __156 _ ( // @[Math.scala 709:24:@76428.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __156 __1 ( // @[Math.scala 709:24:@76435.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_81 fix2fixBox ( // @[Math.scala 141:30:@76445.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@76433.4 Math.scala 713:14:@76434.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@76440.4 Math.scala 713:14:@76441.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@76442.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@76453.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@76431.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@76438.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@76448.4]
endmodule
module fix2fixBox_88( // @[:@77507.2]
  input        clock, // @[:@77508.4]
  input        reset, // @[:@77509.4]
  input  [8:0] io_a, // @[:@77510.4]
  input        io_flow, // @[:@77510.4]
  output [7:0] io_b // @[:@77510.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@77523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@77523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@77523.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@77523.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@77523.4]
  RetimeWrapper_65 RetimeWrapper ( // @[package.scala 93:22:@77523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@77530.4]
  assign RetimeWrapper_clock = clock; // @[:@77524.4]
  assign RetimeWrapper_reset = reset; // @[:@77525.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@77527.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@77526.4]
endmodule
module x1058_sum( // @[:@77532.2]
  input        clock, // @[:@77533.4]
  input        reset, // @[:@77534.4]
  input  [7:0] io_a, // @[:@77535.4]
  input  [7:0] io_b, // @[:@77535.4]
  input        io_flow, // @[:@77535.4]
  output [7:0] io_result // @[:@77535.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@77543.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@77543.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@77550.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@77550.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@77560.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@77560.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@77560.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@77560.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@77560.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@77548.4 Math.scala 713:14:@77549.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@77555.4 Math.scala 713:14:@77556.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@77557.4]
  __156 _ ( // @[Math.scala 709:24:@77543.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __156 __1 ( // @[Math.scala 709:24:@77550.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_88 fix2fixBox ( // @[Math.scala 141:30:@77560.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@77548.4 Math.scala 713:14:@77549.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@77555.4 Math.scala 713:14:@77556.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@77557.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@77568.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@77546.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@77553.4]
  assign fix2fixBox_clock = clock; // @[:@77561.4]
  assign fix2fixBox_reset = reset; // @[:@77562.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@77563.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@77566.4]
endmodule
module RetimeWrapper_997( // @[:@87135.2]
  input         clock, // @[:@87136.4]
  input         reset, // @[:@87137.4]
  input         io_flow, // @[:@87138.4]
  input  [63:0] io_in, // @[:@87138.4]
  output [63:0] io_out // @[:@87138.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@87140.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@87140.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@87140.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@87140.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@87140.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@87140.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@87140.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@87153.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@87152.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@87151.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@87150.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@87149.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@87147.4]
endmodule
module x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@87251.2]
  input          clock, // @[:@87252.4]
  input          reset, // @[:@87253.4]
  output         io_in_x745_TVALID, // @[:@87254.4]
  input          io_in_x745_TREADY, // @[:@87254.4]
  output [255:0] io_in_x745_TDATA, // @[:@87254.4]
  output         io_in_x744_TREADY, // @[:@87254.4]
  input  [255:0] io_in_x744_TDATA, // @[:@87254.4]
  input  [7:0]   io_in_x744_TID, // @[:@87254.4]
  input  [7:0]   io_in_x744_TDEST, // @[:@87254.4]
  input          io_sigsIn_backpressure, // @[:@87254.4]
  input          io_sigsIn_datapathEn, // @[:@87254.4]
  input          io_sigsIn_break, // @[:@87254.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@87254.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@87254.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@87254.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@87254.4]
  input          io_rr // @[:@87254.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@87268.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@87268.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@87280.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@87280.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@87303.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@87303.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@87303.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@87303.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@87303.4]
  wire  x805_lb_0_clock; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_reset; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_29_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_29_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_29_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_29_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_29_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_29_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_28_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_28_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_28_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_28_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_28_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_28_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_27_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_27_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_27_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_27_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_27_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_27_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_26_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_26_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_26_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_26_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_26_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_26_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_25_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_25_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_25_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_25_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_25_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_25_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_24_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_24_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_24_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_24_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_24_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_24_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_23_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_23_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_23_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_23_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_23_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_23_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_22_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_22_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_22_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_22_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_22_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_22_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_21_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_21_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_21_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_21_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_21_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_21_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_20_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_20_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_20_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_20_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_20_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_20_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_19_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_19_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_19_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_19_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_19_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_19_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_18_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_18_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_18_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_18_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_18_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_18_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_17_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_17_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_17_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_17_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_17_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_17_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_16_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_16_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_16_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_16_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_16_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_16_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_15_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_15_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_15_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_15_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_15_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_15_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_14_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_14_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_14_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_14_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_14_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_14_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_13_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_13_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_13_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_13_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_13_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_13_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_12_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_12_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_12_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_12_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_12_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_12_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_11_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_11_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_11_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_11_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_11_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_11_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_10_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_10_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_10_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_10_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_10_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_10_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_9_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_9_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_9_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_9_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_9_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_9_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_8_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_8_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_8_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_8_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_8_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_8_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_7_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_7_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_7_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_7_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_7_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_7_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_6_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_6_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_6_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_6_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_6_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_6_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_5_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_5_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_5_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_5_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_5_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_5_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_4_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_4_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_4_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_4_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_4_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_4_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_3_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_3_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_3_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_3_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_3_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_3_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_2_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_2_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_2_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_2_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_2_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_2_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_1_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_1_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_1_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_1_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_1_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_1_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_rPort_0_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_rPort_0_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_0_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_0_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_rPort_0_backpressure; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_rPort_0_output_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_7_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_7_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_7_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_7_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_7_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_6_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_6_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_6_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_6_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_6_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_5_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_5_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_5_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_5_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_5_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_4_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_4_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_4_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_4_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_4_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_3_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_3_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_3_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_3_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_3_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_2_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_2_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_2_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_2_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_2_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_1_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_1_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_1_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_1_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_1_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [3:0] x805_lb_0_io_wPort_0_banks_1; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [2:0] x805_lb_0_io_wPort_0_banks_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_0_ofs_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire [7:0] x805_lb_0_io_wPort_0_data_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  x805_lb_0_io_wPort_0_en_0; // @[m_x805_lb_0.scala 63:17:@87313.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@87631.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@87631.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@87631.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@87631.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@87631.4]
  wire  x814_1_clock; // @[Math.scala 366:24:@87653.4]
  wire  x814_1_reset; // @[Math.scala 366:24:@87653.4]
  wire [31:0] x814_1_io_a; // @[Math.scala 366:24:@87653.4]
  wire  x814_1_io_flow; // @[Math.scala 366:24:@87653.4]
  wire [31:0] x814_1_io_result; // @[Math.scala 366:24:@87653.4]
  wire  x1235_sum_1_clock; // @[Math.scala 150:24:@87682.4]
  wire  x1235_sum_1_reset; // @[Math.scala 150:24:@87682.4]
  wire [31:0] x1235_sum_1_io_a; // @[Math.scala 150:24:@87682.4]
  wire [31:0] x1235_sum_1_io_b; // @[Math.scala 150:24:@87682.4]
  wire  x1235_sum_1_io_flow; // @[Math.scala 150:24:@87682.4]
  wire [31:0] x1235_sum_1_io_result; // @[Math.scala 150:24:@87682.4]
  wire  x817_div_1_clock; // @[Math.scala 327:24:@87694.4]
  wire  x817_div_1_reset; // @[Math.scala 327:24:@87694.4]
  wire [31:0] x817_div_1_io_a; // @[Math.scala 327:24:@87694.4]
  wire  x817_div_1_io_flow; // @[Math.scala 327:24:@87694.4]
  wire [31:0] x817_div_1_io_result; // @[Math.scala 327:24:@87694.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@87704.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@87704.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@87704.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@87704.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@87704.4]
  wire  x818_sum_1_clock; // @[Math.scala 150:24:@87713.4]
  wire  x818_sum_1_reset; // @[Math.scala 150:24:@87713.4]
  wire [31:0] x818_sum_1_io_a; // @[Math.scala 150:24:@87713.4]
  wire [31:0] x818_sum_1_io_b; // @[Math.scala 150:24:@87713.4]
  wire  x818_sum_1_io_flow; // @[Math.scala 150:24:@87713.4]
  wire [31:0] x818_sum_1_io_result; // @[Math.scala 150:24:@87713.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@87723.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@87723.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@87723.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@87723.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@87723.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@87732.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@87732.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@87732.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@87732.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@87732.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@87741.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@87741.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@87741.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@87741.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@87741.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@87750.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@87750.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@87750.4]
  wire [7:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@87750.4]
  wire [7:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@87750.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@87759.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@87759.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@87759.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@87759.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@87759.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@87768.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@87768.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@87768.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@87768.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@87768.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@87779.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@87779.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@87779.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@87779.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@87779.4]
  wire  x820_rdcol_1_clock; // @[Math.scala 150:24:@87802.4]
  wire  x820_rdcol_1_reset; // @[Math.scala 150:24:@87802.4]
  wire [31:0] x820_rdcol_1_io_a; // @[Math.scala 150:24:@87802.4]
  wire [31:0] x820_rdcol_1_io_b; // @[Math.scala 150:24:@87802.4]
  wire  x820_rdcol_1_io_flow; // @[Math.scala 150:24:@87802.4]
  wire [31:0] x820_rdcol_1_io_result; // @[Math.scala 150:24:@87802.4]
  wire  x822_1_clock; // @[Math.scala 366:24:@87816.4]
  wire  x822_1_reset; // @[Math.scala 366:24:@87816.4]
  wire [31:0] x822_1_io_a; // @[Math.scala 366:24:@87816.4]
  wire  x822_1_io_flow; // @[Math.scala 366:24:@87816.4]
  wire [31:0] x822_1_io_result; // @[Math.scala 366:24:@87816.4]
  wire  x823_div_1_clock; // @[Math.scala 327:24:@87828.4]
  wire  x823_div_1_reset; // @[Math.scala 327:24:@87828.4]
  wire [31:0] x823_div_1_io_a; // @[Math.scala 327:24:@87828.4]
  wire  x823_div_1_io_flow; // @[Math.scala 327:24:@87828.4]
  wire [31:0] x823_div_1_io_result; // @[Math.scala 327:24:@87828.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@87838.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@87838.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@87838.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@87838.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@87838.4]
  wire  x824_sum_1_clock; // @[Math.scala 150:24:@87847.4]
  wire  x824_sum_1_reset; // @[Math.scala 150:24:@87847.4]
  wire [31:0] x824_sum_1_io_a; // @[Math.scala 150:24:@87847.4]
  wire [31:0] x824_sum_1_io_b; // @[Math.scala 150:24:@87847.4]
  wire  x824_sum_1_io_flow; // @[Math.scala 150:24:@87847.4]
  wire [31:0] x824_sum_1_io_result; // @[Math.scala 150:24:@87847.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@87857.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@87857.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@87857.4]
  wire [7:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@87857.4]
  wire [7:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@87857.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@87866.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@87866.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@87866.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@87866.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@87866.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@87875.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@87875.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@87875.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@87875.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@87875.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@87886.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@87886.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@87886.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@87886.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@87886.4]
  wire  x826_rdcol_1_clock; // @[Math.scala 150:24:@87909.4]
  wire  x826_rdcol_1_reset; // @[Math.scala 150:24:@87909.4]
  wire [31:0] x826_rdcol_1_io_a; // @[Math.scala 150:24:@87909.4]
  wire [31:0] x826_rdcol_1_io_b; // @[Math.scala 150:24:@87909.4]
  wire  x826_rdcol_1_io_flow; // @[Math.scala 150:24:@87909.4]
  wire [31:0] x826_rdcol_1_io_result; // @[Math.scala 150:24:@87909.4]
  wire  x828_1_clock; // @[Math.scala 366:24:@87923.4]
  wire  x828_1_reset; // @[Math.scala 366:24:@87923.4]
  wire [31:0] x828_1_io_a; // @[Math.scala 366:24:@87923.4]
  wire  x828_1_io_flow; // @[Math.scala 366:24:@87923.4]
  wire [31:0] x828_1_io_result; // @[Math.scala 366:24:@87923.4]
  wire  x829_div_1_clock; // @[Math.scala 327:24:@87935.4]
  wire  x829_div_1_reset; // @[Math.scala 327:24:@87935.4]
  wire [31:0] x829_div_1_io_a; // @[Math.scala 327:24:@87935.4]
  wire  x829_div_1_io_flow; // @[Math.scala 327:24:@87935.4]
  wire [31:0] x829_div_1_io_result; // @[Math.scala 327:24:@87935.4]
  wire  x830_sum_1_clock; // @[Math.scala 150:24:@87945.4]
  wire  x830_sum_1_reset; // @[Math.scala 150:24:@87945.4]
  wire [31:0] x830_sum_1_io_a; // @[Math.scala 150:24:@87945.4]
  wire [31:0] x830_sum_1_io_b; // @[Math.scala 150:24:@87945.4]
  wire  x830_sum_1_io_flow; // @[Math.scala 150:24:@87945.4]
  wire [31:0] x830_sum_1_io_result; // @[Math.scala 150:24:@87945.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@87955.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@87955.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@87955.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@87955.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@87955.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@87964.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@87964.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@87964.4]
  wire [7:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@87964.4]
  wire [7:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@87964.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@87973.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@87973.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@87973.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@87973.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@87973.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@87984.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@87984.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@87984.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@87984.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@87984.4]
  wire  x832_rdcol_1_clock; // @[Math.scala 150:24:@88007.4]
  wire  x832_rdcol_1_reset; // @[Math.scala 150:24:@88007.4]
  wire [31:0] x832_rdcol_1_io_a; // @[Math.scala 150:24:@88007.4]
  wire [31:0] x832_rdcol_1_io_b; // @[Math.scala 150:24:@88007.4]
  wire  x832_rdcol_1_io_flow; // @[Math.scala 150:24:@88007.4]
  wire [31:0] x832_rdcol_1_io_result; // @[Math.scala 150:24:@88007.4]
  wire  x834_1_clock; // @[Math.scala 366:24:@88023.4]
  wire  x834_1_reset; // @[Math.scala 366:24:@88023.4]
  wire [31:0] x834_1_io_a; // @[Math.scala 366:24:@88023.4]
  wire  x834_1_io_flow; // @[Math.scala 366:24:@88023.4]
  wire [31:0] x834_1_io_result; // @[Math.scala 366:24:@88023.4]
  wire  x835_div_1_clock; // @[Math.scala 327:24:@88035.4]
  wire  x835_div_1_reset; // @[Math.scala 327:24:@88035.4]
  wire [31:0] x835_div_1_io_a; // @[Math.scala 327:24:@88035.4]
  wire  x835_div_1_io_flow; // @[Math.scala 327:24:@88035.4]
  wire [31:0] x835_div_1_io_result; // @[Math.scala 327:24:@88035.4]
  wire  x836_sum_1_clock; // @[Math.scala 150:24:@88045.4]
  wire  x836_sum_1_reset; // @[Math.scala 150:24:@88045.4]
  wire [31:0] x836_sum_1_io_a; // @[Math.scala 150:24:@88045.4]
  wire [31:0] x836_sum_1_io_b; // @[Math.scala 150:24:@88045.4]
  wire  x836_sum_1_io_flow; // @[Math.scala 150:24:@88045.4]
  wire [31:0] x836_sum_1_io_result; // @[Math.scala 150:24:@88045.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@88055.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@88055.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@88055.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@88055.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@88055.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@88064.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@88064.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@88064.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@88064.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@88064.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@88073.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@88073.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@88073.4]
  wire [7:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@88073.4]
  wire [7:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@88073.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@88084.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@88084.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@88084.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@88084.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@88084.4]
  wire  x838_rdcol_1_clock; // @[Math.scala 150:24:@88107.4]
  wire  x838_rdcol_1_reset; // @[Math.scala 150:24:@88107.4]
  wire [31:0] x838_rdcol_1_io_a; // @[Math.scala 150:24:@88107.4]
  wire [31:0] x838_rdcol_1_io_b; // @[Math.scala 150:24:@88107.4]
  wire  x838_rdcol_1_io_flow; // @[Math.scala 150:24:@88107.4]
  wire [31:0] x838_rdcol_1_io_result; // @[Math.scala 150:24:@88107.4]
  wire  x840_1_clock; // @[Math.scala 366:24:@88121.4]
  wire  x840_1_reset; // @[Math.scala 366:24:@88121.4]
  wire [31:0] x840_1_io_a; // @[Math.scala 366:24:@88121.4]
  wire  x840_1_io_flow; // @[Math.scala 366:24:@88121.4]
  wire [31:0] x840_1_io_result; // @[Math.scala 366:24:@88121.4]
  wire  x841_div_1_clock; // @[Math.scala 327:24:@88133.4]
  wire  x841_div_1_reset; // @[Math.scala 327:24:@88133.4]
  wire [31:0] x841_div_1_io_a; // @[Math.scala 327:24:@88133.4]
  wire  x841_div_1_io_flow; // @[Math.scala 327:24:@88133.4]
  wire [31:0] x841_div_1_io_result; // @[Math.scala 327:24:@88133.4]
  wire  x842_sum_1_clock; // @[Math.scala 150:24:@88143.4]
  wire  x842_sum_1_reset; // @[Math.scala 150:24:@88143.4]
  wire [31:0] x842_sum_1_io_a; // @[Math.scala 150:24:@88143.4]
  wire [31:0] x842_sum_1_io_b; // @[Math.scala 150:24:@88143.4]
  wire  x842_sum_1_io_flow; // @[Math.scala 150:24:@88143.4]
  wire [31:0] x842_sum_1_io_result; // @[Math.scala 150:24:@88143.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@88153.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@88153.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@88153.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@88153.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@88153.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@88162.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@88162.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@88162.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@88162.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@88162.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@88171.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@88171.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@88171.4]
  wire [7:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@88171.4]
  wire [7:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@88171.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@88182.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@88182.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@88182.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@88182.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@88182.4]
  wire  x844_rdcol_1_clock; // @[Math.scala 150:24:@88205.4]
  wire  x844_rdcol_1_reset; // @[Math.scala 150:24:@88205.4]
  wire [31:0] x844_rdcol_1_io_a; // @[Math.scala 150:24:@88205.4]
  wire [31:0] x844_rdcol_1_io_b; // @[Math.scala 150:24:@88205.4]
  wire  x844_rdcol_1_io_flow; // @[Math.scala 150:24:@88205.4]
  wire [31:0] x844_rdcol_1_io_result; // @[Math.scala 150:24:@88205.4]
  wire  x846_1_clock; // @[Math.scala 366:24:@88219.4]
  wire  x846_1_reset; // @[Math.scala 366:24:@88219.4]
  wire [31:0] x846_1_io_a; // @[Math.scala 366:24:@88219.4]
  wire  x846_1_io_flow; // @[Math.scala 366:24:@88219.4]
  wire [31:0] x846_1_io_result; // @[Math.scala 366:24:@88219.4]
  wire  x847_div_1_clock; // @[Math.scala 327:24:@88231.4]
  wire  x847_div_1_reset; // @[Math.scala 327:24:@88231.4]
  wire [31:0] x847_div_1_io_a; // @[Math.scala 327:24:@88231.4]
  wire  x847_div_1_io_flow; // @[Math.scala 327:24:@88231.4]
  wire [31:0] x847_div_1_io_result; // @[Math.scala 327:24:@88231.4]
  wire  x848_sum_1_clock; // @[Math.scala 150:24:@88241.4]
  wire  x848_sum_1_reset; // @[Math.scala 150:24:@88241.4]
  wire [31:0] x848_sum_1_io_a; // @[Math.scala 150:24:@88241.4]
  wire [31:0] x848_sum_1_io_b; // @[Math.scala 150:24:@88241.4]
  wire  x848_sum_1_io_flow; // @[Math.scala 150:24:@88241.4]
  wire [31:0] x848_sum_1_io_result; // @[Math.scala 150:24:@88241.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@88251.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@88251.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@88251.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@88251.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@88251.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@88260.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@88260.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@88260.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@88260.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@88260.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@88269.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@88269.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@88269.4]
  wire [7:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@88269.4]
  wire [7:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@88269.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@88280.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@88280.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@88280.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@88280.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@88280.4]
  wire  x850_rdcol_1_clock; // @[Math.scala 150:24:@88303.4]
  wire  x850_rdcol_1_reset; // @[Math.scala 150:24:@88303.4]
  wire [31:0] x850_rdcol_1_io_a; // @[Math.scala 150:24:@88303.4]
  wire [31:0] x850_rdcol_1_io_b; // @[Math.scala 150:24:@88303.4]
  wire  x850_rdcol_1_io_flow; // @[Math.scala 150:24:@88303.4]
  wire [31:0] x850_rdcol_1_io_result; // @[Math.scala 150:24:@88303.4]
  wire  x852_1_clock; // @[Math.scala 366:24:@88317.4]
  wire  x852_1_reset; // @[Math.scala 366:24:@88317.4]
  wire [31:0] x852_1_io_a; // @[Math.scala 366:24:@88317.4]
  wire  x852_1_io_flow; // @[Math.scala 366:24:@88317.4]
  wire [31:0] x852_1_io_result; // @[Math.scala 366:24:@88317.4]
  wire  x853_div_1_clock; // @[Math.scala 327:24:@88329.4]
  wire  x853_div_1_reset; // @[Math.scala 327:24:@88329.4]
  wire [31:0] x853_div_1_io_a; // @[Math.scala 327:24:@88329.4]
  wire  x853_div_1_io_flow; // @[Math.scala 327:24:@88329.4]
  wire [31:0] x853_div_1_io_result; // @[Math.scala 327:24:@88329.4]
  wire  x854_sum_1_clock; // @[Math.scala 150:24:@88339.4]
  wire  x854_sum_1_reset; // @[Math.scala 150:24:@88339.4]
  wire [31:0] x854_sum_1_io_a; // @[Math.scala 150:24:@88339.4]
  wire [31:0] x854_sum_1_io_b; // @[Math.scala 150:24:@88339.4]
  wire  x854_sum_1_io_flow; // @[Math.scala 150:24:@88339.4]
  wire [31:0] x854_sum_1_io_result; // @[Math.scala 150:24:@88339.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@88349.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@88349.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@88349.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@88349.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@88349.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@88358.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@88358.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@88358.4]
  wire [7:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@88358.4]
  wire [7:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@88358.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@88367.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@88367.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@88367.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@88367.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@88367.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@88378.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@88378.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@88378.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@88378.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@88378.4]
  wire  x856_rdcol_1_clock; // @[Math.scala 150:24:@88401.4]
  wire  x856_rdcol_1_reset; // @[Math.scala 150:24:@88401.4]
  wire [31:0] x856_rdcol_1_io_a; // @[Math.scala 150:24:@88401.4]
  wire [31:0] x856_rdcol_1_io_b; // @[Math.scala 150:24:@88401.4]
  wire  x856_rdcol_1_io_flow; // @[Math.scala 150:24:@88401.4]
  wire [31:0] x856_rdcol_1_io_result; // @[Math.scala 150:24:@88401.4]
  wire  x858_1_clock; // @[Math.scala 366:24:@88415.4]
  wire  x858_1_reset; // @[Math.scala 366:24:@88415.4]
  wire [31:0] x858_1_io_a; // @[Math.scala 366:24:@88415.4]
  wire  x858_1_io_flow; // @[Math.scala 366:24:@88415.4]
  wire [31:0] x858_1_io_result; // @[Math.scala 366:24:@88415.4]
  wire  x859_div_1_clock; // @[Math.scala 327:24:@88427.4]
  wire  x859_div_1_reset; // @[Math.scala 327:24:@88427.4]
  wire [31:0] x859_div_1_io_a; // @[Math.scala 327:24:@88427.4]
  wire  x859_div_1_io_flow; // @[Math.scala 327:24:@88427.4]
  wire [31:0] x859_div_1_io_result; // @[Math.scala 327:24:@88427.4]
  wire  x860_sum_1_clock; // @[Math.scala 150:24:@88437.4]
  wire  x860_sum_1_reset; // @[Math.scala 150:24:@88437.4]
  wire [31:0] x860_sum_1_io_a; // @[Math.scala 150:24:@88437.4]
  wire [31:0] x860_sum_1_io_b; // @[Math.scala 150:24:@88437.4]
  wire  x860_sum_1_io_flow; // @[Math.scala 150:24:@88437.4]
  wire [31:0] x860_sum_1_io_result; // @[Math.scala 150:24:@88437.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@88447.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@88447.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@88447.4]
  wire [7:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@88447.4]
  wire [7:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@88447.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@88456.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@88456.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@88456.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@88456.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@88456.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@88465.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@88465.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@88465.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@88465.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@88465.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@88476.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@88476.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@88476.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@88476.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@88476.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@88497.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@88497.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@88497.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@88497.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@88497.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@88513.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@88513.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@88513.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@88513.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@88513.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@88531.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@88531.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@88531.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@88531.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@88531.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@88540.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@88540.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@88540.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@88540.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@88540.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@88554.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@88554.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@88554.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@88554.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@88554.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@88563.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@88563.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@88563.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@88563.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@88563.4]
  wire  x1240_sum_1_clock; // @[Math.scala 150:24:@88610.4]
  wire  x1240_sum_1_reset; // @[Math.scala 150:24:@88610.4]
  wire [31:0] x1240_sum_1_io_a; // @[Math.scala 150:24:@88610.4]
  wire [31:0] x1240_sum_1_io_b; // @[Math.scala 150:24:@88610.4]
  wire  x1240_sum_1_io_flow; // @[Math.scala 150:24:@88610.4]
  wire [31:0] x1240_sum_1_io_result; // @[Math.scala 150:24:@88610.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@88620.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@88620.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@88620.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@88620.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@88620.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@88629.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@88629.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@88629.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@88629.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@88629.4]
  wire  x871_sum_1_clock; // @[Math.scala 150:24:@88638.4]
  wire  x871_sum_1_reset; // @[Math.scala 150:24:@88638.4]
  wire [31:0] x871_sum_1_io_a; // @[Math.scala 150:24:@88638.4]
  wire [31:0] x871_sum_1_io_b; // @[Math.scala 150:24:@88638.4]
  wire  x871_sum_1_io_flow; // @[Math.scala 150:24:@88638.4]
  wire [31:0] x871_sum_1_io_result; // @[Math.scala 150:24:@88638.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@88648.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@88648.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@88648.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@88648.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@88648.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@88657.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@88657.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@88657.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@88657.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@88657.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@88666.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@88666.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@88666.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@88666.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@88666.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@88675.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@88675.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@88675.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@88675.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@88675.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@88684.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@88684.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@88684.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@88684.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@88684.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@88696.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@88696.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@88696.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@88696.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@88696.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@88717.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@88717.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@88717.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@88717.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@88717.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@88731.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@88731.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@88731.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@88731.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@88731.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@88746.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@88746.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@88746.4]
  wire [31:0] RetimeWrapper_55_io_in; // @[package.scala 93:22:@88746.4]
  wire [31:0] RetimeWrapper_55_io_out; // @[package.scala 93:22:@88746.4]
  wire  x877_sum_1_clock; // @[Math.scala 150:24:@88755.4]
  wire  x877_sum_1_reset; // @[Math.scala 150:24:@88755.4]
  wire [31:0] x877_sum_1_io_a; // @[Math.scala 150:24:@88755.4]
  wire [31:0] x877_sum_1_io_b; // @[Math.scala 150:24:@88755.4]
  wire  x877_sum_1_io_flow; // @[Math.scala 150:24:@88755.4]
  wire [31:0] x877_sum_1_io_result; // @[Math.scala 150:24:@88755.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@88765.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@88765.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@88765.4]
  wire [31:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@88765.4]
  wire [31:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@88765.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@88774.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@88774.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@88774.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@88774.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@88774.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@88786.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@88786.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@88786.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@88786.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@88786.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@88807.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@88807.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@88807.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@88807.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@88807.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@88821.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@88821.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@88821.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@88821.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@88821.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@88836.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@88836.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@88836.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@88836.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@88836.4]
  wire  x883_sum_1_clock; // @[Math.scala 150:24:@88845.4]
  wire  x883_sum_1_reset; // @[Math.scala 150:24:@88845.4]
  wire [31:0] x883_sum_1_io_a; // @[Math.scala 150:24:@88845.4]
  wire [31:0] x883_sum_1_io_b; // @[Math.scala 150:24:@88845.4]
  wire  x883_sum_1_io_flow; // @[Math.scala 150:24:@88845.4]
  wire [31:0] x883_sum_1_io_result; // @[Math.scala 150:24:@88845.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@88855.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@88855.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@88855.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@88855.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@88855.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@88864.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@88864.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@88864.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@88864.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@88864.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@88876.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@88876.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@88876.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@88876.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@88876.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@88897.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@88897.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@88897.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@88897.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@88897.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@88911.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@88911.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@88911.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@88911.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@88911.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@88926.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@88926.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@88926.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@88926.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@88926.4]
  wire  x889_sum_1_clock; // @[Math.scala 150:24:@88935.4]
  wire  x889_sum_1_reset; // @[Math.scala 150:24:@88935.4]
  wire [31:0] x889_sum_1_io_a; // @[Math.scala 150:24:@88935.4]
  wire [31:0] x889_sum_1_io_b; // @[Math.scala 150:24:@88935.4]
  wire  x889_sum_1_io_flow; // @[Math.scala 150:24:@88935.4]
  wire [31:0] x889_sum_1_io_result; // @[Math.scala 150:24:@88935.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@88945.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@88945.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@88945.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@88945.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@88945.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@88954.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@88954.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@88954.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@88954.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@88954.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@88966.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@88966.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@88966.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@88966.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@88966.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@88987.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@88987.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@88987.4]
  wire [31:0] RetimeWrapper_71_io_in; // @[package.scala 93:22:@88987.4]
  wire [31:0] RetimeWrapper_71_io_out; // @[package.scala 93:22:@88987.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@89003.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@89003.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@89003.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@89003.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@89003.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@89018.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@89018.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@89018.4]
  wire [31:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@89018.4]
  wire [31:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@89018.4]
  wire  x895_sum_1_clock; // @[Math.scala 150:24:@89027.4]
  wire  x895_sum_1_reset; // @[Math.scala 150:24:@89027.4]
  wire [31:0] x895_sum_1_io_a; // @[Math.scala 150:24:@89027.4]
  wire [31:0] x895_sum_1_io_b; // @[Math.scala 150:24:@89027.4]
  wire  x895_sum_1_io_flow; // @[Math.scala 150:24:@89027.4]
  wire [31:0] x895_sum_1_io_result; // @[Math.scala 150:24:@89027.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@89037.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@89037.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@89037.4]
  wire [31:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@89037.4]
  wire [31:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@89037.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@89046.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@89046.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@89046.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@89046.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@89046.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@89058.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@89058.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@89058.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@89058.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@89058.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@89079.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@89079.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@89079.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@89079.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@89079.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@89093.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@89093.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@89093.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@89093.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@89093.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@89108.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@89108.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@89108.4]
  wire [31:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@89108.4]
  wire [31:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@89108.4]
  wire  x901_sum_1_clock; // @[Math.scala 150:24:@89117.4]
  wire  x901_sum_1_reset; // @[Math.scala 150:24:@89117.4]
  wire [31:0] x901_sum_1_io_a; // @[Math.scala 150:24:@89117.4]
  wire [31:0] x901_sum_1_io_b; // @[Math.scala 150:24:@89117.4]
  wire  x901_sum_1_io_flow; // @[Math.scala 150:24:@89117.4]
  wire [31:0] x901_sum_1_io_result; // @[Math.scala 150:24:@89117.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@89127.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@89127.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@89127.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@89127.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@89127.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@89136.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@89136.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@89136.4]
  wire [31:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@89136.4]
  wire [31:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@89136.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@89148.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@89148.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@89148.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@89148.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@89148.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@89169.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@89169.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@89169.4]
  wire [31:0] RetimeWrapper_83_io_in; // @[package.scala 93:22:@89169.4]
  wire [31:0] RetimeWrapper_83_io_out; // @[package.scala 93:22:@89169.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@89183.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@89183.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@89183.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@89183.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@89183.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@89198.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@89198.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@89198.4]
  wire [31:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@89198.4]
  wire [31:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@89198.4]
  wire  x907_sum_1_clock; // @[Math.scala 150:24:@89207.4]
  wire  x907_sum_1_reset; // @[Math.scala 150:24:@89207.4]
  wire [31:0] x907_sum_1_io_a; // @[Math.scala 150:24:@89207.4]
  wire [31:0] x907_sum_1_io_b; // @[Math.scala 150:24:@89207.4]
  wire  x907_sum_1_io_flow; // @[Math.scala 150:24:@89207.4]
  wire [31:0] x907_sum_1_io_result; // @[Math.scala 150:24:@89207.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@89217.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@89217.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@89217.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@89217.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@89217.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@89226.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@89226.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@89226.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@89226.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@89226.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@89238.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@89238.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@89238.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@89238.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@89238.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@89259.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@89259.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@89259.4]
  wire [31:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@89259.4]
  wire [31:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@89259.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@89273.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@89273.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@89273.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@89273.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@89273.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@89288.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@89288.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@89288.4]
  wire [31:0] RetimeWrapper_91_io_in; // @[package.scala 93:22:@89288.4]
  wire [31:0] RetimeWrapper_91_io_out; // @[package.scala 93:22:@89288.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@89297.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@89297.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@89297.4]
  wire [31:0] RetimeWrapper_92_io_in; // @[package.scala 93:22:@89297.4]
  wire [31:0] RetimeWrapper_92_io_out; // @[package.scala 93:22:@89297.4]
  wire  x913_sum_1_clock; // @[Math.scala 150:24:@89306.4]
  wire  x913_sum_1_reset; // @[Math.scala 150:24:@89306.4]
  wire [31:0] x913_sum_1_io_a; // @[Math.scala 150:24:@89306.4]
  wire [31:0] x913_sum_1_io_b; // @[Math.scala 150:24:@89306.4]
  wire  x913_sum_1_io_flow; // @[Math.scala 150:24:@89306.4]
  wire [31:0] x913_sum_1_io_result; // @[Math.scala 150:24:@89306.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@89316.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@89316.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@89316.4]
  wire [31:0] RetimeWrapper_93_io_in; // @[package.scala 93:22:@89316.4]
  wire [31:0] RetimeWrapper_93_io_out; // @[package.scala 93:22:@89316.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@89325.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@89325.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@89325.4]
  wire [31:0] RetimeWrapper_94_io_in; // @[package.scala 93:22:@89325.4]
  wire [31:0] RetimeWrapper_94_io_out; // @[package.scala 93:22:@89325.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@89334.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@89334.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@89334.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@89334.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@89334.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@89346.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@89346.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@89346.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@89346.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@89346.4]
  wire  x916_rdcol_1_clock; // @[Math.scala 150:24:@89369.4]
  wire  x916_rdcol_1_reset; // @[Math.scala 150:24:@89369.4]
  wire [31:0] x916_rdcol_1_io_a; // @[Math.scala 150:24:@89369.4]
  wire [31:0] x916_rdcol_1_io_b; // @[Math.scala 150:24:@89369.4]
  wire  x916_rdcol_1_io_flow; // @[Math.scala 150:24:@89369.4]
  wire [31:0] x916_rdcol_1_io_result; // @[Math.scala 150:24:@89369.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@89384.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@89384.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@89384.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@89384.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@89384.4]
  wire  x920_1_clock; // @[Math.scala 366:24:@89401.4]
  wire  x920_1_reset; // @[Math.scala 366:24:@89401.4]
  wire [31:0] x920_1_io_a; // @[Math.scala 366:24:@89401.4]
  wire  x920_1_io_flow; // @[Math.scala 366:24:@89401.4]
  wire [31:0] x920_1_io_result; // @[Math.scala 366:24:@89401.4]
  wire  x921_div_1_clock; // @[Math.scala 327:24:@89413.4]
  wire  x921_div_1_reset; // @[Math.scala 327:24:@89413.4]
  wire [31:0] x921_div_1_io_a; // @[Math.scala 327:24:@89413.4]
  wire  x921_div_1_io_flow; // @[Math.scala 327:24:@89413.4]
  wire [31:0] x921_div_1_io_result; // @[Math.scala 327:24:@89413.4]
  wire  x922_sum_1_clock; // @[Math.scala 150:24:@89423.4]
  wire  x922_sum_1_reset; // @[Math.scala 150:24:@89423.4]
  wire [31:0] x922_sum_1_io_a; // @[Math.scala 150:24:@89423.4]
  wire [31:0] x922_sum_1_io_b; // @[Math.scala 150:24:@89423.4]
  wire  x922_sum_1_io_flow; // @[Math.scala 150:24:@89423.4]
  wire [31:0] x922_sum_1_io_result; // @[Math.scala 150:24:@89423.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@89433.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@89433.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@89433.4]
  wire [31:0] RetimeWrapper_98_io_in; // @[package.scala 93:22:@89433.4]
  wire [31:0] RetimeWrapper_98_io_out; // @[package.scala 93:22:@89433.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@89442.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@89442.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@89442.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@89442.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@89442.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@89454.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@89454.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@89454.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@89454.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@89454.4]
  wire  x925_rdcol_1_clock; // @[Math.scala 150:24:@89479.4]
  wire  x925_rdcol_1_reset; // @[Math.scala 150:24:@89479.4]
  wire [31:0] x925_rdcol_1_io_a; // @[Math.scala 150:24:@89479.4]
  wire [31:0] x925_rdcol_1_io_b; // @[Math.scala 150:24:@89479.4]
  wire  x925_rdcol_1_io_flow; // @[Math.scala 150:24:@89479.4]
  wire [31:0] x925_rdcol_1_io_result; // @[Math.scala 150:24:@89479.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@89494.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@89494.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@89494.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@89494.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@89494.4]
  wire  x929_1_clock; // @[Math.scala 366:24:@89511.4]
  wire  x929_1_reset; // @[Math.scala 366:24:@89511.4]
  wire [31:0] x929_1_io_a; // @[Math.scala 366:24:@89511.4]
  wire  x929_1_io_flow; // @[Math.scala 366:24:@89511.4]
  wire [31:0] x929_1_io_result; // @[Math.scala 366:24:@89511.4]
  wire  x930_div_1_clock; // @[Math.scala 327:24:@89523.4]
  wire  x930_div_1_reset; // @[Math.scala 327:24:@89523.4]
  wire [31:0] x930_div_1_io_a; // @[Math.scala 327:24:@89523.4]
  wire  x930_div_1_io_flow; // @[Math.scala 327:24:@89523.4]
  wire [31:0] x930_div_1_io_result; // @[Math.scala 327:24:@89523.4]
  wire  x931_sum_1_clock; // @[Math.scala 150:24:@89533.4]
  wire  x931_sum_1_reset; // @[Math.scala 150:24:@89533.4]
  wire [31:0] x931_sum_1_io_a; // @[Math.scala 150:24:@89533.4]
  wire [31:0] x931_sum_1_io_b; // @[Math.scala 150:24:@89533.4]
  wire  x931_sum_1_io_flow; // @[Math.scala 150:24:@89533.4]
  wire [31:0] x931_sum_1_io_result; // @[Math.scala 150:24:@89533.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@89543.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@89543.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@89543.4]
  wire [31:0] RetimeWrapper_102_io_in; // @[package.scala 93:22:@89543.4]
  wire [31:0] RetimeWrapper_102_io_out; // @[package.scala 93:22:@89543.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@89552.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@89552.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@89552.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@89552.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@89552.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@89564.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@89564.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@89564.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@89564.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@89564.4]
  wire  x934_rdrow_1_clock; // @[Math.scala 191:24:@89587.4]
  wire  x934_rdrow_1_reset; // @[Math.scala 191:24:@89587.4]
  wire [31:0] x934_rdrow_1_io_a; // @[Math.scala 191:24:@89587.4]
  wire [31:0] x934_rdrow_1_io_b; // @[Math.scala 191:24:@89587.4]
  wire  x934_rdrow_1_io_flow; // @[Math.scala 191:24:@89587.4]
  wire [31:0] x934_rdrow_1_io_result; // @[Math.scala 191:24:@89587.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@89604.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@89604.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@89604.4]
  wire [31:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@89604.4]
  wire [31:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@89604.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@89622.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@89622.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@89622.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@89622.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@89622.4]
  wire  x1245_sum_1_clock; // @[Math.scala 150:24:@89667.4]
  wire  x1245_sum_1_reset; // @[Math.scala 150:24:@89667.4]
  wire [31:0] x1245_sum_1_io_a; // @[Math.scala 150:24:@89667.4]
  wire [31:0] x1245_sum_1_io_b; // @[Math.scala 150:24:@89667.4]
  wire  x1245_sum_1_io_flow; // @[Math.scala 150:24:@89667.4]
  wire [31:0] x1245_sum_1_io_result; // @[Math.scala 150:24:@89667.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@89677.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@89677.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@89677.4]
  wire [31:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@89677.4]
  wire [31:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@89677.4]
  wire  x942_sum_1_clock; // @[Math.scala 150:24:@89686.4]
  wire  x942_sum_1_reset; // @[Math.scala 150:24:@89686.4]
  wire [31:0] x942_sum_1_io_a; // @[Math.scala 150:24:@89686.4]
  wire [31:0] x942_sum_1_io_b; // @[Math.scala 150:24:@89686.4]
  wire  x942_sum_1_io_flow; // @[Math.scala 150:24:@89686.4]
  wire [31:0] x942_sum_1_io_result; // @[Math.scala 150:24:@89686.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@89696.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@89696.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@89696.4]
  wire [31:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@89696.4]
  wire [31:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@89696.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@89705.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@89705.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@89705.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@89705.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@89705.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@89717.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@89717.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@89717.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@89717.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@89717.4]
  wire  x947_sum_1_clock; // @[Math.scala 150:24:@89744.4]
  wire  x947_sum_1_reset; // @[Math.scala 150:24:@89744.4]
  wire [31:0] x947_sum_1_io_a; // @[Math.scala 150:24:@89744.4]
  wire [31:0] x947_sum_1_io_b; // @[Math.scala 150:24:@89744.4]
  wire  x947_sum_1_io_flow; // @[Math.scala 150:24:@89744.4]
  wire [31:0] x947_sum_1_io_result; // @[Math.scala 150:24:@89744.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@89754.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@89754.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@89754.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@89754.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@89754.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@89766.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@89766.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@89766.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@89766.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@89766.4]
  wire  x952_sum_1_clock; // @[Math.scala 150:24:@89793.4]
  wire  x952_sum_1_reset; // @[Math.scala 150:24:@89793.4]
  wire [31:0] x952_sum_1_io_a; // @[Math.scala 150:24:@89793.4]
  wire [31:0] x952_sum_1_io_b; // @[Math.scala 150:24:@89793.4]
  wire  x952_sum_1_io_flow; // @[Math.scala 150:24:@89793.4]
  wire [31:0] x952_sum_1_io_result; // @[Math.scala 150:24:@89793.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@89803.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@89803.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@89803.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@89803.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@89803.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@89815.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@89815.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@89815.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@89815.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@89815.4]
  wire  x957_sum_1_clock; // @[Math.scala 150:24:@89842.4]
  wire  x957_sum_1_reset; // @[Math.scala 150:24:@89842.4]
  wire [31:0] x957_sum_1_io_a; // @[Math.scala 150:24:@89842.4]
  wire [31:0] x957_sum_1_io_b; // @[Math.scala 150:24:@89842.4]
  wire  x957_sum_1_io_flow; // @[Math.scala 150:24:@89842.4]
  wire [31:0] x957_sum_1_io_result; // @[Math.scala 150:24:@89842.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@89852.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@89852.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@89852.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@89852.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@89852.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@89864.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@89864.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@89864.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@89864.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@89864.4]
  wire  x962_sum_1_clock; // @[Math.scala 150:24:@89893.4]
  wire  x962_sum_1_reset; // @[Math.scala 150:24:@89893.4]
  wire [31:0] x962_sum_1_io_a; // @[Math.scala 150:24:@89893.4]
  wire [31:0] x962_sum_1_io_b; // @[Math.scala 150:24:@89893.4]
  wire  x962_sum_1_io_flow; // @[Math.scala 150:24:@89893.4]
  wire [31:0] x962_sum_1_io_result; // @[Math.scala 150:24:@89893.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@89903.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@89903.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@89903.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@89903.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@89903.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@89915.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@89915.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@89915.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@89915.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@89915.4]
  wire  x967_sum_1_clock; // @[Math.scala 150:24:@89942.4]
  wire  x967_sum_1_reset; // @[Math.scala 150:24:@89942.4]
  wire [31:0] x967_sum_1_io_a; // @[Math.scala 150:24:@89942.4]
  wire [31:0] x967_sum_1_io_b; // @[Math.scala 150:24:@89942.4]
  wire  x967_sum_1_io_flow; // @[Math.scala 150:24:@89942.4]
  wire [31:0] x967_sum_1_io_result; // @[Math.scala 150:24:@89942.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@89952.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@89952.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@89952.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@89952.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@89952.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@89964.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@89964.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@89964.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@89964.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@89964.4]
  wire  x972_sum_1_clock; // @[Math.scala 150:24:@89991.4]
  wire  x972_sum_1_reset; // @[Math.scala 150:24:@89991.4]
  wire [31:0] x972_sum_1_io_a; // @[Math.scala 150:24:@89991.4]
  wire [31:0] x972_sum_1_io_b; // @[Math.scala 150:24:@89991.4]
  wire  x972_sum_1_io_flow; // @[Math.scala 150:24:@89991.4]
  wire [31:0] x972_sum_1_io_result; // @[Math.scala 150:24:@89991.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@90001.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@90001.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@90001.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@90001.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@90001.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@90013.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@90013.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@90013.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@90013.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@90013.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@90034.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@90034.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@90034.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@90034.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@90034.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@90049.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@90049.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@90049.4]
  wire [31:0] RetimeWrapper_124_io_in; // @[package.scala 93:22:@90049.4]
  wire [31:0] RetimeWrapper_124_io_out; // @[package.scala 93:22:@90049.4]
  wire  x977_sum_1_clock; // @[Math.scala 150:24:@90058.4]
  wire  x977_sum_1_reset; // @[Math.scala 150:24:@90058.4]
  wire [31:0] x977_sum_1_io_a; // @[Math.scala 150:24:@90058.4]
  wire [31:0] x977_sum_1_io_b; // @[Math.scala 150:24:@90058.4]
  wire  x977_sum_1_io_flow; // @[Math.scala 150:24:@90058.4]
  wire [31:0] x977_sum_1_io_result; // @[Math.scala 150:24:@90058.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@90068.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@90068.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@90068.4]
  wire [31:0] RetimeWrapper_125_io_in; // @[package.scala 93:22:@90068.4]
  wire [31:0] RetimeWrapper_125_io_out; // @[package.scala 93:22:@90068.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@90077.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@90077.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@90077.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@90077.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@90077.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@90089.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@90089.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@90089.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@90089.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@90089.4]
  wire  x982_sum_1_clock; // @[Math.scala 150:24:@90116.4]
  wire  x982_sum_1_reset; // @[Math.scala 150:24:@90116.4]
  wire [31:0] x982_sum_1_io_a; // @[Math.scala 150:24:@90116.4]
  wire [31:0] x982_sum_1_io_b; // @[Math.scala 150:24:@90116.4]
  wire  x982_sum_1_io_flow; // @[Math.scala 150:24:@90116.4]
  wire [31:0] x982_sum_1_io_result; // @[Math.scala 150:24:@90116.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@90126.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@90126.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@90126.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@90126.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@90126.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@90138.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@90138.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@90138.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@90138.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@90138.4]
  wire  x987_sum_1_clock; // @[Math.scala 150:24:@90165.4]
  wire  x987_sum_1_reset; // @[Math.scala 150:24:@90165.4]
  wire [31:0] x987_sum_1_io_a; // @[Math.scala 150:24:@90165.4]
  wire [31:0] x987_sum_1_io_b; // @[Math.scala 150:24:@90165.4]
  wire  x987_sum_1_io_flow; // @[Math.scala 150:24:@90165.4]
  wire [31:0] x987_sum_1_io_result; // @[Math.scala 150:24:@90165.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@90175.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@90175.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@90175.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@90175.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@90175.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@90187.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@90187.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@90187.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@90187.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@90187.4]
  wire  x990_rdrow_1_clock; // @[Math.scala 191:24:@90210.4]
  wire  x990_rdrow_1_reset; // @[Math.scala 191:24:@90210.4]
  wire [31:0] x990_rdrow_1_io_a; // @[Math.scala 191:24:@90210.4]
  wire [31:0] x990_rdrow_1_io_b; // @[Math.scala 191:24:@90210.4]
  wire  x990_rdrow_1_io_flow; // @[Math.scala 191:24:@90210.4]
  wire [31:0] x990_rdrow_1_io_result; // @[Math.scala 191:24:@90210.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@90227.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@90227.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@90227.4]
  wire [31:0] RetimeWrapper_132_io_in; // @[package.scala 93:22:@90227.4]
  wire [31:0] RetimeWrapper_132_io_out; // @[package.scala 93:22:@90227.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@90245.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@90245.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@90245.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@90245.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@90245.4]
  wire  x1250_sum_1_clock; // @[Math.scala 150:24:@90290.4]
  wire  x1250_sum_1_reset; // @[Math.scala 150:24:@90290.4]
  wire [31:0] x1250_sum_1_io_a; // @[Math.scala 150:24:@90290.4]
  wire [31:0] x1250_sum_1_io_b; // @[Math.scala 150:24:@90290.4]
  wire  x1250_sum_1_io_flow; // @[Math.scala 150:24:@90290.4]
  wire [31:0] x1250_sum_1_io_result; // @[Math.scala 150:24:@90290.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@90300.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@90300.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@90300.4]
  wire [31:0] RetimeWrapper_134_io_in; // @[package.scala 93:22:@90300.4]
  wire [31:0] RetimeWrapper_134_io_out; // @[package.scala 93:22:@90300.4]
  wire  x998_sum_1_clock; // @[Math.scala 150:24:@90311.4]
  wire  x998_sum_1_reset; // @[Math.scala 150:24:@90311.4]
  wire [31:0] x998_sum_1_io_a; // @[Math.scala 150:24:@90311.4]
  wire [31:0] x998_sum_1_io_b; // @[Math.scala 150:24:@90311.4]
  wire  x998_sum_1_io_flow; // @[Math.scala 150:24:@90311.4]
  wire [31:0] x998_sum_1_io_result; // @[Math.scala 150:24:@90311.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@90321.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@90321.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@90321.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@90321.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@90321.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@90330.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@90330.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@90330.4]
  wire [31:0] RetimeWrapper_136_io_in; // @[package.scala 93:22:@90330.4]
  wire [31:0] RetimeWrapper_136_io_out; // @[package.scala 93:22:@90330.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@90342.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@90342.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@90342.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@90342.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@90342.4]
  wire  x1003_sum_1_clock; // @[Math.scala 150:24:@90369.4]
  wire  x1003_sum_1_reset; // @[Math.scala 150:24:@90369.4]
  wire [31:0] x1003_sum_1_io_a; // @[Math.scala 150:24:@90369.4]
  wire [31:0] x1003_sum_1_io_b; // @[Math.scala 150:24:@90369.4]
  wire  x1003_sum_1_io_flow; // @[Math.scala 150:24:@90369.4]
  wire [31:0] x1003_sum_1_io_result; // @[Math.scala 150:24:@90369.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@90379.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@90379.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@90379.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@90379.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@90379.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@90391.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@90391.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@90391.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@90391.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@90391.4]
  wire  x1008_sum_1_clock; // @[Math.scala 150:24:@90418.4]
  wire  x1008_sum_1_reset; // @[Math.scala 150:24:@90418.4]
  wire [31:0] x1008_sum_1_io_a; // @[Math.scala 150:24:@90418.4]
  wire [31:0] x1008_sum_1_io_b; // @[Math.scala 150:24:@90418.4]
  wire  x1008_sum_1_io_flow; // @[Math.scala 150:24:@90418.4]
  wire [31:0] x1008_sum_1_io_result; // @[Math.scala 150:24:@90418.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@90428.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@90428.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@90428.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@90428.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@90428.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@90440.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@90440.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@90440.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@90440.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@90440.4]
  wire  x1013_sum_1_clock; // @[Math.scala 150:24:@90467.4]
  wire  x1013_sum_1_reset; // @[Math.scala 150:24:@90467.4]
  wire [31:0] x1013_sum_1_io_a; // @[Math.scala 150:24:@90467.4]
  wire [31:0] x1013_sum_1_io_b; // @[Math.scala 150:24:@90467.4]
  wire  x1013_sum_1_io_flow; // @[Math.scala 150:24:@90467.4]
  wire [31:0] x1013_sum_1_io_result; // @[Math.scala 150:24:@90467.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@90477.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@90477.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@90477.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@90477.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@90477.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@90489.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@90489.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@90489.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@90489.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@90489.4]
  wire  x1018_sum_1_clock; // @[Math.scala 150:24:@90516.4]
  wire  x1018_sum_1_reset; // @[Math.scala 150:24:@90516.4]
  wire [31:0] x1018_sum_1_io_a; // @[Math.scala 150:24:@90516.4]
  wire [31:0] x1018_sum_1_io_b; // @[Math.scala 150:24:@90516.4]
  wire  x1018_sum_1_io_flow; // @[Math.scala 150:24:@90516.4]
  wire [31:0] x1018_sum_1_io_result; // @[Math.scala 150:24:@90516.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@90526.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@90526.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@90526.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@90526.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@90526.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@90538.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@90538.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@90538.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@90538.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@90538.4]
  wire  x1023_sum_1_clock; // @[Math.scala 150:24:@90565.4]
  wire  x1023_sum_1_reset; // @[Math.scala 150:24:@90565.4]
  wire [31:0] x1023_sum_1_io_a; // @[Math.scala 150:24:@90565.4]
  wire [31:0] x1023_sum_1_io_b; // @[Math.scala 150:24:@90565.4]
  wire  x1023_sum_1_io_flow; // @[Math.scala 150:24:@90565.4]
  wire [31:0] x1023_sum_1_io_result; // @[Math.scala 150:24:@90565.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@90575.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@90575.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@90575.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@90575.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@90575.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@90587.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@90587.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@90587.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@90587.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@90587.4]
  wire  x1028_sum_1_clock; // @[Math.scala 150:24:@90614.4]
  wire  x1028_sum_1_reset; // @[Math.scala 150:24:@90614.4]
  wire [31:0] x1028_sum_1_io_a; // @[Math.scala 150:24:@90614.4]
  wire [31:0] x1028_sum_1_io_b; // @[Math.scala 150:24:@90614.4]
  wire  x1028_sum_1_io_flow; // @[Math.scala 150:24:@90614.4]
  wire [31:0] x1028_sum_1_io_result; // @[Math.scala 150:24:@90614.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@90624.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@90624.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@90624.4]
  wire  RetimeWrapper_148_io_in; // @[package.scala 93:22:@90624.4]
  wire  RetimeWrapper_148_io_out; // @[package.scala 93:22:@90624.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@90636.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@90636.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@90636.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@90636.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@90636.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@90663.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@90663.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@90663.4]
  wire [31:0] RetimeWrapper_150_io_in; // @[package.scala 93:22:@90663.4]
  wire [31:0] RetimeWrapper_150_io_out; // @[package.scala 93:22:@90663.4]
  wire  x1033_sum_1_clock; // @[Math.scala 150:24:@90672.4]
  wire  x1033_sum_1_reset; // @[Math.scala 150:24:@90672.4]
  wire [31:0] x1033_sum_1_io_a; // @[Math.scala 150:24:@90672.4]
  wire [31:0] x1033_sum_1_io_b; // @[Math.scala 150:24:@90672.4]
  wire  x1033_sum_1_io_flow; // @[Math.scala 150:24:@90672.4]
  wire [31:0] x1033_sum_1_io_result; // @[Math.scala 150:24:@90672.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@90682.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@90682.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@90682.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@90682.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@90682.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@90691.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@90691.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@90691.4]
  wire [31:0] RetimeWrapper_152_io_in; // @[package.scala 93:22:@90691.4]
  wire [31:0] RetimeWrapper_152_io_out; // @[package.scala 93:22:@90691.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@90703.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@90703.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@90703.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@90703.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@90703.4]
  wire  x1038_sum_1_clock; // @[Math.scala 150:24:@90732.4]
  wire  x1038_sum_1_reset; // @[Math.scala 150:24:@90732.4]
  wire [31:0] x1038_sum_1_io_a; // @[Math.scala 150:24:@90732.4]
  wire [31:0] x1038_sum_1_io_b; // @[Math.scala 150:24:@90732.4]
  wire  x1038_sum_1_io_flow; // @[Math.scala 150:24:@90732.4]
  wire [31:0] x1038_sum_1_io_result; // @[Math.scala 150:24:@90732.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@90742.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@90742.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@90742.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@90742.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@90742.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@90754.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@90754.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@90754.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@90754.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@90754.4]
  wire  x1043_sum_1_clock; // @[Math.scala 150:24:@90781.4]
  wire  x1043_sum_1_reset; // @[Math.scala 150:24:@90781.4]
  wire [31:0] x1043_sum_1_io_a; // @[Math.scala 150:24:@90781.4]
  wire [31:0] x1043_sum_1_io_b; // @[Math.scala 150:24:@90781.4]
  wire  x1043_sum_1_io_flow; // @[Math.scala 150:24:@90781.4]
  wire [31:0] x1043_sum_1_io_result; // @[Math.scala 150:24:@90781.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@90791.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@90791.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@90791.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@90791.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@90791.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@90803.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@90803.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@90803.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@90803.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@90803.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@90826.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@90826.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@90826.4]
  wire [8:0] RetimeWrapper_158_io_in; // @[package.scala 93:22:@90826.4]
  wire [8:0] RetimeWrapper_158_io_out; // @[package.scala 93:22:@90826.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@90838.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@90838.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@90838.4]
  wire [8:0] RetimeWrapper_159_io_in; // @[package.scala 93:22:@90838.4]
  wire [8:0] RetimeWrapper_159_io_out; // @[package.scala 93:22:@90838.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@90850.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@90850.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@90850.4]
  wire [9:0] RetimeWrapper_160_io_in; // @[package.scala 93:22:@90850.4]
  wire [9:0] RetimeWrapper_160_io_out; // @[package.scala 93:22:@90850.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@90862.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@90862.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@90862.4]
  wire [8:0] RetimeWrapper_161_io_in; // @[package.scala 93:22:@90862.4]
  wire [8:0] RetimeWrapper_161_io_out; // @[package.scala 93:22:@90862.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@90874.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@90874.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@90874.4]
  wire [8:0] RetimeWrapper_162_io_in; // @[package.scala 93:22:@90874.4]
  wire [8:0] RetimeWrapper_162_io_out; // @[package.scala 93:22:@90874.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@90884.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@90884.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@90884.4]
  wire [7:0] RetimeWrapper_163_io_in; // @[package.scala 93:22:@90884.4]
  wire [7:0] RetimeWrapper_163_io_out; // @[package.scala 93:22:@90884.4]
  wire [7:0] x1051_x15_1_io_a; // @[Math.scala 150:24:@90893.4]
  wire [7:0] x1051_x15_1_io_b; // @[Math.scala 150:24:@90893.4]
  wire [7:0] x1051_x15_1_io_result; // @[Math.scala 150:24:@90893.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@90903.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@90903.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@90903.4]
  wire [7:0] RetimeWrapper_164_io_in; // @[package.scala 93:22:@90903.4]
  wire [7:0] RetimeWrapper_164_io_out; // @[package.scala 93:22:@90903.4]
  wire [7:0] x1052_x16_1_io_a; // @[Math.scala 150:24:@90912.4]
  wire [7:0] x1052_x16_1_io_b; // @[Math.scala 150:24:@90912.4]
  wire [7:0] x1052_x16_1_io_result; // @[Math.scala 150:24:@90912.4]
  wire [7:0] x1053_x15_1_io_a; // @[Math.scala 150:24:@90922.4]
  wire [7:0] x1053_x15_1_io_b; // @[Math.scala 150:24:@90922.4]
  wire [7:0] x1053_x15_1_io_result; // @[Math.scala 150:24:@90922.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@90932.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@90932.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@90932.4]
  wire [7:0] RetimeWrapper_165_io_in; // @[package.scala 93:22:@90932.4]
  wire [7:0] RetimeWrapper_165_io_out; // @[package.scala 93:22:@90932.4]
  wire [7:0] x1054_x16_1_io_a; // @[Math.scala 150:24:@90941.4]
  wire [7:0] x1054_x16_1_io_b; // @[Math.scala 150:24:@90941.4]
  wire [7:0] x1054_x16_1_io_result; // @[Math.scala 150:24:@90941.4]
  wire [7:0] x1055_x15_1_io_a; // @[Math.scala 150:24:@90951.4]
  wire [7:0] x1055_x15_1_io_b; // @[Math.scala 150:24:@90951.4]
  wire [7:0] x1055_x15_1_io_result; // @[Math.scala 150:24:@90951.4]
  wire [7:0] x1056_x16_1_io_a; // @[Math.scala 150:24:@90961.4]
  wire [7:0] x1056_x16_1_io_b; // @[Math.scala 150:24:@90961.4]
  wire [7:0] x1056_x16_1_io_result; // @[Math.scala 150:24:@90961.4]
  wire [7:0] x1057_x15_1_io_a; // @[Math.scala 150:24:@90971.4]
  wire [7:0] x1057_x15_1_io_b; // @[Math.scala 150:24:@90971.4]
  wire [7:0] x1057_x15_1_io_result; // @[Math.scala 150:24:@90971.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@90981.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@90981.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@90981.4]
  wire [7:0] RetimeWrapper_166_io_in; // @[package.scala 93:22:@90981.4]
  wire [7:0] RetimeWrapper_166_io_out; // @[package.scala 93:22:@90981.4]
  wire  x1058_sum_1_clock; // @[Math.scala 150:24:@90990.4]
  wire  x1058_sum_1_reset; // @[Math.scala 150:24:@90990.4]
  wire [7:0] x1058_sum_1_io_a; // @[Math.scala 150:24:@90990.4]
  wire [7:0] x1058_sum_1_io_b; // @[Math.scala 150:24:@90990.4]
  wire  x1058_sum_1_io_flow; // @[Math.scala 150:24:@90990.4]
  wire [7:0] x1058_sum_1_io_result; // @[Math.scala 150:24:@90990.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@91009.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@91009.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@91009.4]
  wire [8:0] RetimeWrapper_167_io_in; // @[package.scala 93:22:@91009.4]
  wire [8:0] RetimeWrapper_167_io_out; // @[package.scala 93:22:@91009.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@91021.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@91021.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@91021.4]
  wire [8:0] RetimeWrapper_168_io_in; // @[package.scala 93:22:@91021.4]
  wire [8:0] RetimeWrapper_168_io_out; // @[package.scala 93:22:@91021.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@91033.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@91033.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@91033.4]
  wire [9:0] RetimeWrapper_169_io_in; // @[package.scala 93:22:@91033.4]
  wire [9:0] RetimeWrapper_169_io_out; // @[package.scala 93:22:@91033.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@91045.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@91045.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@91045.4]
  wire [8:0] RetimeWrapper_170_io_in; // @[package.scala 93:22:@91045.4]
  wire [8:0] RetimeWrapper_170_io_out; // @[package.scala 93:22:@91045.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@91057.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@91057.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@91057.4]
  wire [8:0] RetimeWrapper_171_io_in; // @[package.scala 93:22:@91057.4]
  wire [8:0] RetimeWrapper_171_io_out; // @[package.scala 93:22:@91057.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@91067.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@91067.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@91067.4]
  wire [7:0] RetimeWrapper_172_io_in; // @[package.scala 93:22:@91067.4]
  wire [7:0] RetimeWrapper_172_io_out; // @[package.scala 93:22:@91067.4]
  wire [7:0] x1065_x15_1_io_a; // @[Math.scala 150:24:@91076.4]
  wire [7:0] x1065_x15_1_io_b; // @[Math.scala 150:24:@91076.4]
  wire [7:0] x1065_x15_1_io_result; // @[Math.scala 150:24:@91076.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@91086.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@91086.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@91086.4]
  wire [7:0] RetimeWrapper_173_io_in; // @[package.scala 93:22:@91086.4]
  wire [7:0] RetimeWrapper_173_io_out; // @[package.scala 93:22:@91086.4]
  wire [7:0] x1066_x16_1_io_a; // @[Math.scala 150:24:@91095.4]
  wire [7:0] x1066_x16_1_io_b; // @[Math.scala 150:24:@91095.4]
  wire [7:0] x1066_x16_1_io_result; // @[Math.scala 150:24:@91095.4]
  wire [7:0] x1067_x15_1_io_a; // @[Math.scala 150:24:@91105.4]
  wire [7:0] x1067_x15_1_io_b; // @[Math.scala 150:24:@91105.4]
  wire [7:0] x1067_x15_1_io_result; // @[Math.scala 150:24:@91105.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@91115.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@91115.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@91115.4]
  wire [7:0] RetimeWrapper_174_io_in; // @[package.scala 93:22:@91115.4]
  wire [7:0] RetimeWrapper_174_io_out; // @[package.scala 93:22:@91115.4]
  wire [7:0] x1068_x16_1_io_a; // @[Math.scala 150:24:@91124.4]
  wire [7:0] x1068_x16_1_io_b; // @[Math.scala 150:24:@91124.4]
  wire [7:0] x1068_x16_1_io_result; // @[Math.scala 150:24:@91124.4]
  wire [7:0] x1069_x15_1_io_a; // @[Math.scala 150:24:@91134.4]
  wire [7:0] x1069_x15_1_io_b; // @[Math.scala 150:24:@91134.4]
  wire [7:0] x1069_x15_1_io_result; // @[Math.scala 150:24:@91134.4]
  wire [7:0] x1070_x16_1_io_a; // @[Math.scala 150:24:@91144.4]
  wire [7:0] x1070_x16_1_io_b; // @[Math.scala 150:24:@91144.4]
  wire [7:0] x1070_x16_1_io_result; // @[Math.scala 150:24:@91144.4]
  wire [7:0] x1071_x15_1_io_a; // @[Math.scala 150:24:@91154.4]
  wire [7:0] x1071_x15_1_io_b; // @[Math.scala 150:24:@91154.4]
  wire [7:0] x1071_x15_1_io_result; // @[Math.scala 150:24:@91154.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@91164.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@91164.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@91164.4]
  wire [7:0] RetimeWrapper_175_io_in; // @[package.scala 93:22:@91164.4]
  wire [7:0] RetimeWrapper_175_io_out; // @[package.scala 93:22:@91164.4]
  wire  x1072_sum_1_clock; // @[Math.scala 150:24:@91173.4]
  wire  x1072_sum_1_reset; // @[Math.scala 150:24:@91173.4]
  wire [7:0] x1072_sum_1_io_a; // @[Math.scala 150:24:@91173.4]
  wire [7:0] x1072_sum_1_io_b; // @[Math.scala 150:24:@91173.4]
  wire  x1072_sum_1_io_flow; // @[Math.scala 150:24:@91173.4]
  wire [7:0] x1072_sum_1_io_result; // @[Math.scala 150:24:@91173.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@91192.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@91192.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@91192.4]
  wire [8:0] RetimeWrapper_176_io_in; // @[package.scala 93:22:@91192.4]
  wire [8:0] RetimeWrapper_176_io_out; // @[package.scala 93:22:@91192.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@91206.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@91206.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@91206.4]
  wire [9:0] RetimeWrapper_177_io_in; // @[package.scala 93:22:@91206.4]
  wire [9:0] RetimeWrapper_177_io_out; // @[package.scala 93:22:@91206.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@91218.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@91218.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@91218.4]
  wire [8:0] RetimeWrapper_178_io_in; // @[package.scala 93:22:@91218.4]
  wire [8:0] RetimeWrapper_178_io_out; // @[package.scala 93:22:@91218.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@91230.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@91230.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@91230.4]
  wire [8:0] RetimeWrapper_179_io_in; // @[package.scala 93:22:@91230.4]
  wire [8:0] RetimeWrapper_179_io_out; // @[package.scala 93:22:@91230.4]
  wire [7:0] x1078_x15_1_io_a; // @[Math.scala 150:24:@91240.4]
  wire [7:0] x1078_x15_1_io_b; // @[Math.scala 150:24:@91240.4]
  wire [7:0] x1078_x15_1_io_result; // @[Math.scala 150:24:@91240.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@91250.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@91250.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@91250.4]
  wire [7:0] RetimeWrapper_180_io_in; // @[package.scala 93:22:@91250.4]
  wire [7:0] RetimeWrapper_180_io_out; // @[package.scala 93:22:@91250.4]
  wire [7:0] x1079_x16_1_io_a; // @[Math.scala 150:24:@91259.4]
  wire [7:0] x1079_x16_1_io_b; // @[Math.scala 150:24:@91259.4]
  wire [7:0] x1079_x16_1_io_result; // @[Math.scala 150:24:@91259.4]
  wire [7:0] x1080_x15_1_io_a; // @[Math.scala 150:24:@91269.4]
  wire [7:0] x1080_x15_1_io_b; // @[Math.scala 150:24:@91269.4]
  wire [7:0] x1080_x15_1_io_result; // @[Math.scala 150:24:@91269.4]
  wire [7:0] x1081_x16_1_io_a; // @[Math.scala 150:24:@91279.4]
  wire [7:0] x1081_x16_1_io_b; // @[Math.scala 150:24:@91279.4]
  wire [7:0] x1081_x16_1_io_result; // @[Math.scala 150:24:@91279.4]
  wire [7:0] x1082_x15_1_io_a; // @[Math.scala 150:24:@91289.4]
  wire [7:0] x1082_x15_1_io_b; // @[Math.scala 150:24:@91289.4]
  wire [7:0] x1082_x15_1_io_result; // @[Math.scala 150:24:@91289.4]
  wire [7:0] x1083_x16_1_io_a; // @[Math.scala 150:24:@91299.4]
  wire [7:0] x1083_x16_1_io_b; // @[Math.scala 150:24:@91299.4]
  wire [7:0] x1083_x16_1_io_result; // @[Math.scala 150:24:@91299.4]
  wire [7:0] x1084_x15_1_io_a; // @[Math.scala 150:24:@91309.4]
  wire [7:0] x1084_x15_1_io_b; // @[Math.scala 150:24:@91309.4]
  wire [7:0] x1084_x15_1_io_result; // @[Math.scala 150:24:@91309.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@91319.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@91319.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@91319.4]
  wire [7:0] RetimeWrapper_181_io_in; // @[package.scala 93:22:@91319.4]
  wire [7:0] RetimeWrapper_181_io_out; // @[package.scala 93:22:@91319.4]
  wire  x1085_sum_1_clock; // @[Math.scala 150:24:@91328.4]
  wire  x1085_sum_1_reset; // @[Math.scala 150:24:@91328.4]
  wire [7:0] x1085_sum_1_io_a; // @[Math.scala 150:24:@91328.4]
  wire [7:0] x1085_sum_1_io_b; // @[Math.scala 150:24:@91328.4]
  wire  x1085_sum_1_io_flow; // @[Math.scala 150:24:@91328.4]
  wire [7:0] x1085_sum_1_io_result; // @[Math.scala 150:24:@91328.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@91347.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@91347.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@91347.4]
  wire [8:0] RetimeWrapper_182_io_in; // @[package.scala 93:22:@91347.4]
  wire [8:0] RetimeWrapper_182_io_out; // @[package.scala 93:22:@91347.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@91359.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@91359.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@91359.4]
  wire [9:0] RetimeWrapper_183_io_in; // @[package.scala 93:22:@91359.4]
  wire [9:0] RetimeWrapper_183_io_out; // @[package.scala 93:22:@91359.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@91371.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@91371.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@91371.4]
  wire [8:0] RetimeWrapper_184_io_in; // @[package.scala 93:22:@91371.4]
  wire [8:0] RetimeWrapper_184_io_out; // @[package.scala 93:22:@91371.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@91383.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@91383.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@91383.4]
  wire [8:0] RetimeWrapper_185_io_in; // @[package.scala 93:22:@91383.4]
  wire [8:0] RetimeWrapper_185_io_out; // @[package.scala 93:22:@91383.4]
  wire [7:0] x1091_x15_1_io_a; // @[Math.scala 150:24:@91393.4]
  wire [7:0] x1091_x15_1_io_b; // @[Math.scala 150:24:@91393.4]
  wire [7:0] x1091_x15_1_io_result; // @[Math.scala 150:24:@91393.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@91403.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@91403.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@91403.4]
  wire [7:0] RetimeWrapper_186_io_in; // @[package.scala 93:22:@91403.4]
  wire [7:0] RetimeWrapper_186_io_out; // @[package.scala 93:22:@91403.4]
  wire [7:0] x1092_x16_1_io_a; // @[Math.scala 150:24:@91412.4]
  wire [7:0] x1092_x16_1_io_b; // @[Math.scala 150:24:@91412.4]
  wire [7:0] x1092_x16_1_io_result; // @[Math.scala 150:24:@91412.4]
  wire [7:0] x1093_x15_1_io_a; // @[Math.scala 150:24:@91422.4]
  wire [7:0] x1093_x15_1_io_b; // @[Math.scala 150:24:@91422.4]
  wire [7:0] x1093_x15_1_io_result; // @[Math.scala 150:24:@91422.4]
  wire [7:0] x1094_x16_1_io_a; // @[Math.scala 150:24:@91432.4]
  wire [7:0] x1094_x16_1_io_b; // @[Math.scala 150:24:@91432.4]
  wire [7:0] x1094_x16_1_io_result; // @[Math.scala 150:24:@91432.4]
  wire [7:0] x1095_x15_1_io_a; // @[Math.scala 150:24:@91442.4]
  wire [7:0] x1095_x15_1_io_b; // @[Math.scala 150:24:@91442.4]
  wire [7:0] x1095_x15_1_io_result; // @[Math.scala 150:24:@91442.4]
  wire [7:0] x1096_x16_1_io_a; // @[Math.scala 150:24:@91452.4]
  wire [7:0] x1096_x16_1_io_b; // @[Math.scala 150:24:@91452.4]
  wire [7:0] x1096_x16_1_io_result; // @[Math.scala 150:24:@91452.4]
  wire [7:0] x1097_x15_1_io_a; // @[Math.scala 150:24:@91462.4]
  wire [7:0] x1097_x15_1_io_b; // @[Math.scala 150:24:@91462.4]
  wire [7:0] x1097_x15_1_io_result; // @[Math.scala 150:24:@91462.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@91472.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@91472.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@91472.4]
  wire [7:0] RetimeWrapper_187_io_in; // @[package.scala 93:22:@91472.4]
  wire [7:0] RetimeWrapper_187_io_out; // @[package.scala 93:22:@91472.4]
  wire  x1098_sum_1_clock; // @[Math.scala 150:24:@91481.4]
  wire  x1098_sum_1_reset; // @[Math.scala 150:24:@91481.4]
  wire [7:0] x1098_sum_1_io_a; // @[Math.scala 150:24:@91481.4]
  wire [7:0] x1098_sum_1_io_b; // @[Math.scala 150:24:@91481.4]
  wire  x1098_sum_1_io_flow; // @[Math.scala 150:24:@91481.4]
  wire [7:0] x1098_sum_1_io_result; // @[Math.scala 150:24:@91481.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@91500.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@91500.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@91500.4]
  wire [8:0] RetimeWrapper_188_io_in; // @[package.scala 93:22:@91500.4]
  wire [8:0] RetimeWrapper_188_io_out; // @[package.scala 93:22:@91500.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@91512.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@91512.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@91512.4]
  wire [9:0] RetimeWrapper_189_io_in; // @[package.scala 93:22:@91512.4]
  wire [9:0] RetimeWrapper_189_io_out; // @[package.scala 93:22:@91512.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@91524.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@91524.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@91524.4]
  wire [8:0] RetimeWrapper_190_io_in; // @[package.scala 93:22:@91524.4]
  wire [8:0] RetimeWrapper_190_io_out; // @[package.scala 93:22:@91524.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@91536.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@91536.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@91536.4]
  wire [8:0] RetimeWrapper_191_io_in; // @[package.scala 93:22:@91536.4]
  wire [8:0] RetimeWrapper_191_io_out; // @[package.scala 93:22:@91536.4]
  wire [7:0] x1104_x15_1_io_a; // @[Math.scala 150:24:@91546.4]
  wire [7:0] x1104_x15_1_io_b; // @[Math.scala 150:24:@91546.4]
  wire [7:0] x1104_x15_1_io_result; // @[Math.scala 150:24:@91546.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@91556.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@91556.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@91556.4]
  wire [7:0] RetimeWrapper_192_io_in; // @[package.scala 93:22:@91556.4]
  wire [7:0] RetimeWrapper_192_io_out; // @[package.scala 93:22:@91556.4]
  wire [7:0] x1105_x16_1_io_a; // @[Math.scala 150:24:@91565.4]
  wire [7:0] x1105_x16_1_io_b; // @[Math.scala 150:24:@91565.4]
  wire [7:0] x1105_x16_1_io_result; // @[Math.scala 150:24:@91565.4]
  wire [7:0] x1106_x15_1_io_a; // @[Math.scala 150:24:@91575.4]
  wire [7:0] x1106_x15_1_io_b; // @[Math.scala 150:24:@91575.4]
  wire [7:0] x1106_x15_1_io_result; // @[Math.scala 150:24:@91575.4]
  wire [7:0] x1107_x16_1_io_a; // @[Math.scala 150:24:@91585.4]
  wire [7:0] x1107_x16_1_io_b; // @[Math.scala 150:24:@91585.4]
  wire [7:0] x1107_x16_1_io_result; // @[Math.scala 150:24:@91585.4]
  wire [7:0] x1108_x15_1_io_a; // @[Math.scala 150:24:@91595.4]
  wire [7:0] x1108_x15_1_io_b; // @[Math.scala 150:24:@91595.4]
  wire [7:0] x1108_x15_1_io_result; // @[Math.scala 150:24:@91595.4]
  wire [7:0] x1109_x16_1_io_a; // @[Math.scala 150:24:@91605.4]
  wire [7:0] x1109_x16_1_io_b; // @[Math.scala 150:24:@91605.4]
  wire [7:0] x1109_x16_1_io_result; // @[Math.scala 150:24:@91605.4]
  wire [7:0] x1110_x15_1_io_a; // @[Math.scala 150:24:@91615.4]
  wire [7:0] x1110_x15_1_io_b; // @[Math.scala 150:24:@91615.4]
  wire [7:0] x1110_x15_1_io_result; // @[Math.scala 150:24:@91615.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@91625.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@91625.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@91625.4]
  wire [7:0] RetimeWrapper_193_io_in; // @[package.scala 93:22:@91625.4]
  wire [7:0] RetimeWrapper_193_io_out; // @[package.scala 93:22:@91625.4]
  wire  x1111_sum_1_clock; // @[Math.scala 150:24:@91634.4]
  wire  x1111_sum_1_reset; // @[Math.scala 150:24:@91634.4]
  wire [7:0] x1111_sum_1_io_a; // @[Math.scala 150:24:@91634.4]
  wire [7:0] x1111_sum_1_io_b; // @[Math.scala 150:24:@91634.4]
  wire  x1111_sum_1_io_flow; // @[Math.scala 150:24:@91634.4]
  wire [7:0] x1111_sum_1_io_result; // @[Math.scala 150:24:@91634.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@91653.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@91653.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@91653.4]
  wire [8:0] RetimeWrapper_194_io_in; // @[package.scala 93:22:@91653.4]
  wire [8:0] RetimeWrapper_194_io_out; // @[package.scala 93:22:@91653.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@91665.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@91665.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@91665.4]
  wire [9:0] RetimeWrapper_195_io_in; // @[package.scala 93:22:@91665.4]
  wire [9:0] RetimeWrapper_195_io_out; // @[package.scala 93:22:@91665.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@91677.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@91677.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@91677.4]
  wire [8:0] RetimeWrapper_196_io_in; // @[package.scala 93:22:@91677.4]
  wire [8:0] RetimeWrapper_196_io_out; // @[package.scala 93:22:@91677.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@91689.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@91689.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@91689.4]
  wire [8:0] RetimeWrapper_197_io_in; // @[package.scala 93:22:@91689.4]
  wire [8:0] RetimeWrapper_197_io_out; // @[package.scala 93:22:@91689.4]
  wire [7:0] x1117_x15_1_io_a; // @[Math.scala 150:24:@91699.4]
  wire [7:0] x1117_x15_1_io_b; // @[Math.scala 150:24:@91699.4]
  wire [7:0] x1117_x15_1_io_result; // @[Math.scala 150:24:@91699.4]
  wire  RetimeWrapper_198_clock; // @[package.scala 93:22:@91709.4]
  wire  RetimeWrapper_198_reset; // @[package.scala 93:22:@91709.4]
  wire  RetimeWrapper_198_io_flow; // @[package.scala 93:22:@91709.4]
  wire [7:0] RetimeWrapper_198_io_in; // @[package.scala 93:22:@91709.4]
  wire [7:0] RetimeWrapper_198_io_out; // @[package.scala 93:22:@91709.4]
  wire [7:0] x1118_x16_1_io_a; // @[Math.scala 150:24:@91720.4]
  wire [7:0] x1118_x16_1_io_b; // @[Math.scala 150:24:@91720.4]
  wire [7:0] x1118_x16_1_io_result; // @[Math.scala 150:24:@91720.4]
  wire [7:0] x1119_x15_1_io_a; // @[Math.scala 150:24:@91730.4]
  wire [7:0] x1119_x15_1_io_b; // @[Math.scala 150:24:@91730.4]
  wire [7:0] x1119_x15_1_io_result; // @[Math.scala 150:24:@91730.4]
  wire [7:0] x1120_x16_1_io_a; // @[Math.scala 150:24:@91740.4]
  wire [7:0] x1120_x16_1_io_b; // @[Math.scala 150:24:@91740.4]
  wire [7:0] x1120_x16_1_io_result; // @[Math.scala 150:24:@91740.4]
  wire [7:0] x1121_x15_1_io_a; // @[Math.scala 150:24:@91750.4]
  wire [7:0] x1121_x15_1_io_b; // @[Math.scala 150:24:@91750.4]
  wire [7:0] x1121_x15_1_io_result; // @[Math.scala 150:24:@91750.4]
  wire [7:0] x1122_x16_1_io_a; // @[Math.scala 150:24:@91760.4]
  wire [7:0] x1122_x16_1_io_b; // @[Math.scala 150:24:@91760.4]
  wire [7:0] x1122_x16_1_io_result; // @[Math.scala 150:24:@91760.4]
  wire [7:0] x1123_x15_1_io_a; // @[Math.scala 150:24:@91770.4]
  wire [7:0] x1123_x15_1_io_b; // @[Math.scala 150:24:@91770.4]
  wire [7:0] x1123_x15_1_io_result; // @[Math.scala 150:24:@91770.4]
  wire  RetimeWrapper_199_clock; // @[package.scala 93:22:@91780.4]
  wire  RetimeWrapper_199_reset; // @[package.scala 93:22:@91780.4]
  wire  RetimeWrapper_199_io_flow; // @[package.scala 93:22:@91780.4]
  wire [7:0] RetimeWrapper_199_io_in; // @[package.scala 93:22:@91780.4]
  wire [7:0] RetimeWrapper_199_io_out; // @[package.scala 93:22:@91780.4]
  wire  x1124_sum_1_clock; // @[Math.scala 150:24:@91789.4]
  wire  x1124_sum_1_reset; // @[Math.scala 150:24:@91789.4]
  wire [7:0] x1124_sum_1_io_a; // @[Math.scala 150:24:@91789.4]
  wire [7:0] x1124_sum_1_io_b; // @[Math.scala 150:24:@91789.4]
  wire  x1124_sum_1_io_flow; // @[Math.scala 150:24:@91789.4]
  wire [7:0] x1124_sum_1_io_result; // @[Math.scala 150:24:@91789.4]
  wire  RetimeWrapper_200_clock; // @[package.scala 93:22:@91808.4]
  wire  RetimeWrapper_200_reset; // @[package.scala 93:22:@91808.4]
  wire  RetimeWrapper_200_io_flow; // @[package.scala 93:22:@91808.4]
  wire [8:0] RetimeWrapper_200_io_in; // @[package.scala 93:22:@91808.4]
  wire [8:0] RetimeWrapper_200_io_out; // @[package.scala 93:22:@91808.4]
  wire  RetimeWrapper_201_clock; // @[package.scala 93:22:@91820.4]
  wire  RetimeWrapper_201_reset; // @[package.scala 93:22:@91820.4]
  wire  RetimeWrapper_201_io_flow; // @[package.scala 93:22:@91820.4]
  wire [9:0] RetimeWrapper_201_io_in; // @[package.scala 93:22:@91820.4]
  wire [9:0] RetimeWrapper_201_io_out; // @[package.scala 93:22:@91820.4]
  wire  RetimeWrapper_202_clock; // @[package.scala 93:22:@91832.4]
  wire  RetimeWrapper_202_reset; // @[package.scala 93:22:@91832.4]
  wire  RetimeWrapper_202_io_flow; // @[package.scala 93:22:@91832.4]
  wire [8:0] RetimeWrapper_202_io_in; // @[package.scala 93:22:@91832.4]
  wire [8:0] RetimeWrapper_202_io_out; // @[package.scala 93:22:@91832.4]
  wire  RetimeWrapper_203_clock; // @[package.scala 93:22:@91844.4]
  wire  RetimeWrapper_203_reset; // @[package.scala 93:22:@91844.4]
  wire  RetimeWrapper_203_io_flow; // @[package.scala 93:22:@91844.4]
  wire [8:0] RetimeWrapper_203_io_in; // @[package.scala 93:22:@91844.4]
  wire [8:0] RetimeWrapper_203_io_out; // @[package.scala 93:22:@91844.4]
  wire [7:0] x1130_x15_1_io_a; // @[Math.scala 150:24:@91854.4]
  wire [7:0] x1130_x15_1_io_b; // @[Math.scala 150:24:@91854.4]
  wire [7:0] x1130_x15_1_io_result; // @[Math.scala 150:24:@91854.4]
  wire  RetimeWrapper_204_clock; // @[package.scala 93:22:@91864.4]
  wire  RetimeWrapper_204_reset; // @[package.scala 93:22:@91864.4]
  wire  RetimeWrapper_204_io_flow; // @[package.scala 93:22:@91864.4]
  wire [7:0] RetimeWrapper_204_io_in; // @[package.scala 93:22:@91864.4]
  wire [7:0] RetimeWrapper_204_io_out; // @[package.scala 93:22:@91864.4]
  wire [7:0] x1131_x16_1_io_a; // @[Math.scala 150:24:@91873.4]
  wire [7:0] x1131_x16_1_io_b; // @[Math.scala 150:24:@91873.4]
  wire [7:0] x1131_x16_1_io_result; // @[Math.scala 150:24:@91873.4]
  wire [7:0] x1132_x15_1_io_a; // @[Math.scala 150:24:@91883.4]
  wire [7:0] x1132_x15_1_io_b; // @[Math.scala 150:24:@91883.4]
  wire [7:0] x1132_x15_1_io_result; // @[Math.scala 150:24:@91883.4]
  wire [7:0] x1133_x16_1_io_a; // @[Math.scala 150:24:@91893.4]
  wire [7:0] x1133_x16_1_io_b; // @[Math.scala 150:24:@91893.4]
  wire [7:0] x1133_x16_1_io_result; // @[Math.scala 150:24:@91893.4]
  wire [7:0] x1134_x15_1_io_a; // @[Math.scala 150:24:@91903.4]
  wire [7:0] x1134_x15_1_io_b; // @[Math.scala 150:24:@91903.4]
  wire [7:0] x1134_x15_1_io_result; // @[Math.scala 150:24:@91903.4]
  wire [7:0] x1135_x16_1_io_a; // @[Math.scala 150:24:@91913.4]
  wire [7:0] x1135_x16_1_io_b; // @[Math.scala 150:24:@91913.4]
  wire [7:0] x1135_x16_1_io_result; // @[Math.scala 150:24:@91913.4]
  wire [7:0] x1136_x15_1_io_a; // @[Math.scala 150:24:@91923.4]
  wire [7:0] x1136_x15_1_io_b; // @[Math.scala 150:24:@91923.4]
  wire [7:0] x1136_x15_1_io_result; // @[Math.scala 150:24:@91923.4]
  wire  RetimeWrapper_205_clock; // @[package.scala 93:22:@91933.4]
  wire  RetimeWrapper_205_reset; // @[package.scala 93:22:@91933.4]
  wire  RetimeWrapper_205_io_flow; // @[package.scala 93:22:@91933.4]
  wire [7:0] RetimeWrapper_205_io_in; // @[package.scala 93:22:@91933.4]
  wire [7:0] RetimeWrapper_205_io_out; // @[package.scala 93:22:@91933.4]
  wire  x1137_sum_1_clock; // @[Math.scala 150:24:@91942.4]
  wire  x1137_sum_1_reset; // @[Math.scala 150:24:@91942.4]
  wire [7:0] x1137_sum_1_io_a; // @[Math.scala 150:24:@91942.4]
  wire [7:0] x1137_sum_1_io_b; // @[Math.scala 150:24:@91942.4]
  wire  x1137_sum_1_io_flow; // @[Math.scala 150:24:@91942.4]
  wire [7:0] x1137_sum_1_io_result; // @[Math.scala 150:24:@91942.4]
  wire  RetimeWrapper_206_clock; // @[package.scala 93:22:@91961.4]
  wire  RetimeWrapper_206_reset; // @[package.scala 93:22:@91961.4]
  wire  RetimeWrapper_206_io_flow; // @[package.scala 93:22:@91961.4]
  wire [8:0] RetimeWrapper_206_io_in; // @[package.scala 93:22:@91961.4]
  wire [8:0] RetimeWrapper_206_io_out; // @[package.scala 93:22:@91961.4]
  wire  RetimeWrapper_207_clock; // @[package.scala 93:22:@91973.4]
  wire  RetimeWrapper_207_reset; // @[package.scala 93:22:@91973.4]
  wire  RetimeWrapper_207_io_flow; // @[package.scala 93:22:@91973.4]
  wire [9:0] RetimeWrapper_207_io_in; // @[package.scala 93:22:@91973.4]
  wire [9:0] RetimeWrapper_207_io_out; // @[package.scala 93:22:@91973.4]
  wire  RetimeWrapper_208_clock; // @[package.scala 93:22:@91985.4]
  wire  RetimeWrapper_208_reset; // @[package.scala 93:22:@91985.4]
  wire  RetimeWrapper_208_io_flow; // @[package.scala 93:22:@91985.4]
  wire [8:0] RetimeWrapper_208_io_in; // @[package.scala 93:22:@91985.4]
  wire [8:0] RetimeWrapper_208_io_out; // @[package.scala 93:22:@91985.4]
  wire  RetimeWrapper_209_clock; // @[package.scala 93:22:@91997.4]
  wire  RetimeWrapper_209_reset; // @[package.scala 93:22:@91997.4]
  wire  RetimeWrapper_209_io_flow; // @[package.scala 93:22:@91997.4]
  wire [8:0] RetimeWrapper_209_io_in; // @[package.scala 93:22:@91997.4]
  wire [8:0] RetimeWrapper_209_io_out; // @[package.scala 93:22:@91997.4]
  wire [7:0] x1143_x15_1_io_a; // @[Math.scala 150:24:@92007.4]
  wire [7:0] x1143_x15_1_io_b; // @[Math.scala 150:24:@92007.4]
  wire [7:0] x1143_x15_1_io_result; // @[Math.scala 150:24:@92007.4]
  wire  RetimeWrapper_210_clock; // @[package.scala 93:22:@92017.4]
  wire  RetimeWrapper_210_reset; // @[package.scala 93:22:@92017.4]
  wire  RetimeWrapper_210_io_flow; // @[package.scala 93:22:@92017.4]
  wire [7:0] RetimeWrapper_210_io_in; // @[package.scala 93:22:@92017.4]
  wire [7:0] RetimeWrapper_210_io_out; // @[package.scala 93:22:@92017.4]
  wire [7:0] x1144_x16_1_io_a; // @[Math.scala 150:24:@92026.4]
  wire [7:0] x1144_x16_1_io_b; // @[Math.scala 150:24:@92026.4]
  wire [7:0] x1144_x16_1_io_result; // @[Math.scala 150:24:@92026.4]
  wire [7:0] x1145_x15_1_io_a; // @[Math.scala 150:24:@92036.4]
  wire [7:0] x1145_x15_1_io_b; // @[Math.scala 150:24:@92036.4]
  wire [7:0] x1145_x15_1_io_result; // @[Math.scala 150:24:@92036.4]
  wire [7:0] x1146_x16_1_io_a; // @[Math.scala 150:24:@92046.4]
  wire [7:0] x1146_x16_1_io_b; // @[Math.scala 150:24:@92046.4]
  wire [7:0] x1146_x16_1_io_result; // @[Math.scala 150:24:@92046.4]
  wire [7:0] x1147_x15_1_io_a; // @[Math.scala 150:24:@92056.4]
  wire [7:0] x1147_x15_1_io_b; // @[Math.scala 150:24:@92056.4]
  wire [7:0] x1147_x15_1_io_result; // @[Math.scala 150:24:@92056.4]
  wire [7:0] x1148_x16_1_io_a; // @[Math.scala 150:24:@92066.4]
  wire [7:0] x1148_x16_1_io_b; // @[Math.scala 150:24:@92066.4]
  wire [7:0] x1148_x16_1_io_result; // @[Math.scala 150:24:@92066.4]
  wire [7:0] x1149_x15_1_io_a; // @[Math.scala 150:24:@92076.4]
  wire [7:0] x1149_x15_1_io_b; // @[Math.scala 150:24:@92076.4]
  wire [7:0] x1149_x15_1_io_result; // @[Math.scala 150:24:@92076.4]
  wire  RetimeWrapper_211_clock; // @[package.scala 93:22:@92086.4]
  wire  RetimeWrapper_211_reset; // @[package.scala 93:22:@92086.4]
  wire  RetimeWrapper_211_io_flow; // @[package.scala 93:22:@92086.4]
  wire [7:0] RetimeWrapper_211_io_in; // @[package.scala 93:22:@92086.4]
  wire [7:0] RetimeWrapper_211_io_out; // @[package.scala 93:22:@92086.4]
  wire  x1150_sum_1_clock; // @[Math.scala 150:24:@92095.4]
  wire  x1150_sum_1_reset; // @[Math.scala 150:24:@92095.4]
  wire [7:0] x1150_sum_1_io_a; // @[Math.scala 150:24:@92095.4]
  wire [7:0] x1150_sum_1_io_b; // @[Math.scala 150:24:@92095.4]
  wire  x1150_sum_1_io_flow; // @[Math.scala 150:24:@92095.4]
  wire [7:0] x1150_sum_1_io_result; // @[Math.scala 150:24:@92095.4]
  wire  RetimeWrapper_212_clock; // @[package.scala 93:22:@92130.4]
  wire  RetimeWrapper_212_reset; // @[package.scala 93:22:@92130.4]
  wire  RetimeWrapper_212_io_flow; // @[package.scala 93:22:@92130.4]
  wire [63:0] RetimeWrapper_212_io_in; // @[package.scala 93:22:@92130.4]
  wire [63:0] RetimeWrapper_212_io_out; // @[package.scala 93:22:@92130.4]
  wire  RetimeWrapper_213_clock; // @[package.scala 93:22:@92139.4]
  wire  RetimeWrapper_213_reset; // @[package.scala 93:22:@92139.4]
  wire  RetimeWrapper_213_io_flow; // @[package.scala 93:22:@92139.4]
  wire  RetimeWrapper_213_io_in; // @[package.scala 93:22:@92139.4]
  wire  RetimeWrapper_213_io_out; // @[package.scala 93:22:@92139.4]
  wire  RetimeWrapper_214_clock; // @[package.scala 93:22:@92148.4]
  wire  RetimeWrapper_214_reset; // @[package.scala 93:22:@92148.4]
  wire  RetimeWrapper_214_io_flow; // @[package.scala 93:22:@92148.4]
  wire  RetimeWrapper_214_io_in; // @[package.scala 93:22:@92148.4]
  wire  RetimeWrapper_214_io_out; // @[package.scala 93:22:@92148.4]
  wire  RetimeWrapper_215_clock; // @[package.scala 93:22:@92157.4]
  wire  RetimeWrapper_215_reset; // @[package.scala 93:22:@92157.4]
  wire  RetimeWrapper_215_io_flow; // @[package.scala 93:22:@92157.4]
  wire  RetimeWrapper_215_io_in; // @[package.scala 93:22:@92157.4]
  wire  RetimeWrapper_215_io_out; // @[package.scala 93:22:@92157.4]
  wire  b801; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 62:18:@87288.4]
  wire  b802; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 63:18:@87289.4]
  wire  _T_205; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 67:30:@87291.4]
  wire  _T_206; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 67:37:@87292.4]
  wire  _T_210; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 69:76:@87297.4]
  wire  _T_211; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 69:62:@87298.4]
  wire  _T_213; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 69:101:@87299.4]
  wire [63:0] x1256_x803_D1_0_number; // @[package.scala 96:25:@87308.4 package.scala 96:25:@87309.4]
  wire [31:0] b799_number; // @[Math.scala 712:22:@87273.4 Math.scala 713:14:@87274.4]
  wire [31:0] _T_254; // @[Math.scala 499:52:@87585.4]
  wire  x808; // @[Math.scala 499:44:@87593.4]
  wire  x809; // @[Math.scala 499:44:@87600.4]
  wire  x810; // @[Math.scala 499:44:@87607.4]
  wire [31:0] _T_301; // @[Mux.scala 19:72:@87619.4]
  wire [31:0] _T_303; // @[Mux.scala 19:72:@87620.4]
  wire [31:0] _T_305; // @[Mux.scala 19:72:@87621.4]
  wire [31:0] _T_307; // @[Mux.scala 19:72:@87623.4]
  wire [31:0] x1257_x811_D2_number; // @[package.scala 96:25:@87636.4 package.scala 96:25:@87637.4]
  wire [31:0] _T_322; // @[Math.scala 406:49:@87643.4]
  wire [31:0] _T_324; // @[Math.scala 406:56:@87645.4]
  wire [31:0] _T_325; // @[Math.scala 406:56:@87646.4]
  wire  _T_337; // @[FixedPoint.scala 50:25:@87664.4]
  wire [1:0] _T_341; // @[Bitwise.scala 72:12:@87666.4]
  wire [29:0] _T_342; // @[FixedPoint.scala 18:52:@87667.4]
  wire [31:0] x815_number; // @[Cat.scala 30:58:@87668.4]
  wire [38:0] _GEN_0; // @[Math.scala 450:32:@87673.4]
  wire [38:0] _T_347; // @[Math.scala 450:32:@87673.4]
  wire [37:0] _GEN_1; // @[Math.scala 450:32:@87678.4]
  wire [37:0] _T_351; // @[Math.scala 450:32:@87678.4]
  wire  _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:101:@87776.4]
  wire  _T_391; // @[package.scala 96:25:@87784.4 package.scala 96:25:@87785.4]
  wire  _T_393; // @[implicits.scala 55:10:@87786.4]
  wire  _T_394; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:118:@87787.4]
  wire  _T_396; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:207:@87789.4]
  wire  _T_397; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:226:@87790.4]
  wire  x1264_b801_D28; // @[package.scala 96:25:@87773.4 package.scala 96:25:@87774.4]
  wire  _T_398; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:252:@87791.4]
  wire  x1260_b802_D28; // @[package.scala 96:25:@87737.4 package.scala 96:25:@87738.4]
  wire  _T_442; // @[package.scala 96:25:@87891.4 package.scala 96:25:@87892.4]
  wire  _T_444; // @[implicits.scala 55:10:@87893.4]
  wire  _T_445; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:118:@87894.4]
  wire  _T_447; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:207:@87896.4]
  wire  _T_448; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:226:@87897.4]
  wire  _T_449; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:252:@87898.4]
  wire  _T_490; // @[package.scala 96:25:@87989.4 package.scala 96:25:@87990.4]
  wire  _T_492; // @[implicits.scala 55:10:@87991.4]
  wire  _T_493; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:118:@87992.4]
  wire  _T_495; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:207:@87994.4]
  wire  _T_496; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:226:@87995.4]
  wire  _T_497; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:252:@87996.4]
  wire  _T_540; // @[package.scala 96:25:@88089.4 package.scala 96:25:@88090.4]
  wire  _T_542; // @[implicits.scala 55:10:@88091.4]
  wire  _T_543; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:166:@88092.4]
  wire  _T_545; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:255:@88094.4]
  wire  _T_546; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:274:@88095.4]
  wire  _T_547; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:300:@88096.4]
  wire  _T_588; // @[package.scala 96:25:@88187.4 package.scala 96:25:@88188.4]
  wire  _T_590; // @[implicits.scala 55:10:@88189.4]
  wire  _T_591; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:166:@88190.4]
  wire  _T_593; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:255:@88192.4]
  wire  _T_594; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:274:@88193.4]
  wire  _T_595; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:300:@88194.4]
  wire  _T_636; // @[package.scala 96:25:@88285.4 package.scala 96:25:@88286.4]
  wire  _T_638; // @[implicits.scala 55:10:@88287.4]
  wire  _T_639; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:166:@88288.4]
  wire  _T_641; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:255:@88290.4]
  wire  _T_642; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:274:@88291.4]
  wire  _T_643; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:300:@88292.4]
  wire  _T_684; // @[package.scala 96:25:@88383.4 package.scala 96:25:@88384.4]
  wire  _T_686; // @[implicits.scala 55:10:@88385.4]
  wire  _T_687; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:166:@88386.4]
  wire  _T_689; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:255:@88388.4]
  wire  _T_690; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:274:@88389.4]
  wire  _T_691; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:300:@88390.4]
  wire  _T_732; // @[package.scala 96:25:@88481.4 package.scala 96:25:@88482.4]
  wire  _T_734; // @[implicits.scala 55:10:@88483.4]
  wire  _T_735; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:166:@88484.4]
  wire  _T_737; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:255:@88486.4]
  wire  _T_738; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:274:@88487.4]
  wire  _T_739; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:300:@88488.4]
  wire [31:0] x1287_b799_D30_number; // @[package.scala 96:25:@88502.4 package.scala 96:25:@88503.4]
  wire [31:0] _T_751; // @[Math.scala 406:49:@88509.4]
  wire [31:0] _T_753; // @[Math.scala 406:56:@88511.4]
  wire [31:0] _T_754; // @[Math.scala 406:56:@88512.4]
  wire [31:0] _T_758; // @[package.scala 96:25:@88520.4]
  wire [31:0] x1236_number; // @[implicits.scala 133:21:@88522.4]
  wire [31:0] x1288_x856_rdcol_D30_number; // @[package.scala 96:25:@88545.4 package.scala 96:25:@88546.4]
  wire [31:0] _T_778; // @[Math.scala 465:37:@88551.4]
  wire  x1289_x864_D1; // @[package.scala 96:25:@88568.4 package.scala 96:25:@88569.4]
  wire  x865; // @[package.scala 96:25:@88559.4 package.scala 96:25:@88560.4]
  wire  x866; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 305:25:@88572.4]
  wire [31:0] _T_799; // @[Math.scala 406:49:@88583.4]
  wire [31:0] _T_801; // @[Math.scala 406:56:@88585.4]
  wire [31:0] _T_802; // @[Math.scala 406:56:@88586.4]
  wire  _T_807; // @[FixedPoint.scala 50:25:@88592.4]
  wire [1:0] _T_811; // @[Bitwise.scala 72:12:@88594.4]
  wire [29:0] _T_812; // @[FixedPoint.scala 18:52:@88595.4]
  wire [31:0] x869_number; // @[Cat.scala 30:58:@88596.4]
  wire [38:0] _GEN_2; // @[Math.scala 450:32:@88601.4]
  wire [38:0] _T_817; // @[Math.scala 450:32:@88601.4]
  wire [37:0] _GEN_3; // @[Math.scala 450:32:@88606.4]
  wire [37:0] _T_821; // @[Math.scala 450:32:@88606.4]
  wire  _T_860; // @[package.scala 96:25:@88701.4 package.scala 96:25:@88702.4]
  wire  _T_862; // @[implicits.scala 55:10:@88703.4]
  wire  _T_863; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 340:194:@88704.4]
  wire  x1295_x867_D20; // @[package.scala 96:25:@88680.4 package.scala 96:25:@88681.4]
  wire  _T_864; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 340:283:@88705.4]
  wire  x1296_b801_D52; // @[package.scala 96:25:@88689.4 package.scala 96:25:@88690.4]
  wire  _T_865; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 340:292:@88706.4]
  wire  x1293_b802_D52; // @[package.scala 96:25:@88662.4 package.scala 96:25:@88663.4]
  wire [31:0] x1297_x850_rdcol_D30_number; // @[package.scala 96:25:@88722.4 package.scala 96:25:@88723.4]
  wire [31:0] _T_876; // @[Math.scala 465:37:@88728.4]
  wire  x874; // @[package.scala 96:25:@88736.4 package.scala 96:25:@88737.4]
  wire  x875; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 348:25:@88740.4]
  wire  _T_908; // @[package.scala 96:25:@88791.4 package.scala 96:25:@88792.4]
  wire  _T_910; // @[implicits.scala 55:10:@88793.4]
  wire  _T_911; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:194:@88794.4]
  wire  x1300_x876_D20; // @[package.scala 96:25:@88779.4 package.scala 96:25:@88780.4]
  wire  _T_912; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:283:@88795.4]
  wire  _T_913; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:292:@88796.4]
  wire [31:0] x1301_x844_rdcol_D30_number; // @[package.scala 96:25:@88812.4 package.scala 96:25:@88813.4]
  wire [31:0] _T_924; // @[Math.scala 465:37:@88818.4]
  wire  x880; // @[package.scala 96:25:@88826.4 package.scala 96:25:@88827.4]
  wire  x881; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 371:25:@88830.4]
  wire  _T_956; // @[package.scala 96:25:@88881.4 package.scala 96:25:@88882.4]
  wire  _T_958; // @[implicits.scala 55:10:@88883.4]
  wire  _T_959; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:194:@88884.4]
  wire  x1304_x882_D20; // @[package.scala 96:25:@88869.4 package.scala 96:25:@88870.4]
  wire  _T_960; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:283:@88885.4]
  wire  _T_961; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:292:@88886.4]
  wire [31:0] x1305_x838_rdcol_D30_number; // @[package.scala 96:25:@88902.4 package.scala 96:25:@88903.4]
  wire [31:0] _T_972; // @[Math.scala 465:37:@88908.4]
  wire  x886; // @[package.scala 96:25:@88916.4 package.scala 96:25:@88917.4]
  wire  x887; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 394:25:@88920.4]
  wire  _T_1004; // @[package.scala 96:25:@88971.4 package.scala 96:25:@88972.4]
  wire  _T_1006; // @[implicits.scala 55:10:@88973.4]
  wire  _T_1007; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:194:@88974.4]
  wire  x1307_x888_D20; // @[package.scala 96:25:@88950.4 package.scala 96:25:@88951.4]
  wire  _T_1008; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:283:@88975.4]
  wire  _T_1009; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:292:@88976.4]
  wire [31:0] x1309_x832_rdcol_D30_number; // @[package.scala 96:25:@88992.4 package.scala 96:25:@88993.4]
  wire [31:0] _T_1022; // @[Math.scala 465:37:@89000.4]
  wire  x892; // @[package.scala 96:25:@89008.4 package.scala 96:25:@89009.4]
  wire  x893; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 425:60:@89012.4]
  wire  _T_1054; // @[package.scala 96:25:@89063.4 package.scala 96:25:@89064.4]
  wire  _T_1056; // @[implicits.scala 55:10:@89065.4]
  wire  _T_1057; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:194:@89066.4]
  wire  x1312_x894_D20; // @[package.scala 96:25:@89051.4 package.scala 96:25:@89052.4]
  wire  _T_1058; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:283:@89067.4]
  wire  _T_1059; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:292:@89068.4]
  wire [31:0] x1313_x826_rdcol_D30_number; // @[package.scala 96:25:@89084.4 package.scala 96:25:@89085.4]
  wire [31:0] _T_1070; // @[Math.scala 465:37:@89090.4]
  wire  x898; // @[package.scala 96:25:@89098.4 package.scala 96:25:@89099.4]
  wire  x899; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 448:60:@89102.4]
  wire  _T_1102; // @[package.scala 96:25:@89153.4 package.scala 96:25:@89154.4]
  wire  _T_1104; // @[implicits.scala 55:10:@89155.4]
  wire  _T_1105; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:194:@89156.4]
  wire  x1315_x900_D20; // @[package.scala 96:25:@89132.4 package.scala 96:25:@89133.4]
  wire  _T_1106; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:283:@89157.4]
  wire  _T_1107; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:292:@89158.4]
  wire [31:0] x1317_x820_rdcol_D30_number; // @[package.scala 96:25:@89174.4 package.scala 96:25:@89175.4]
  wire [31:0] _T_1118; // @[Math.scala 465:37:@89180.4]
  wire  x904; // @[package.scala 96:25:@89188.4 package.scala 96:25:@89189.4]
  wire  x905; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 471:60:@89192.4]
  wire  _T_1150; // @[package.scala 96:25:@89243.4 package.scala 96:25:@89244.4]
  wire  _T_1152; // @[implicits.scala 55:10:@89245.4]
  wire  _T_1153; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:194:@89246.4]
  wire  x1319_x906_D20; // @[package.scala 96:25:@89222.4 package.scala 96:25:@89223.4]
  wire  _T_1154; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:283:@89247.4]
  wire  _T_1155; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:292:@89248.4]
  wire [31:0] x1321_b800_D30_number; // @[package.scala 96:25:@89264.4 package.scala 96:25:@89265.4]
  wire [31:0] _T_1166; // @[Math.scala 465:37:@89270.4]
  wire  x864; // @[package.scala 96:25:@88536.4 package.scala 96:25:@88537.4]
  wire  x910; // @[package.scala 96:25:@89278.4 package.scala 96:25:@89279.4]
  wire  x911; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 494:59:@89282.4]
  wire  _T_1204; // @[package.scala 96:25:@89351.4 package.scala 96:25:@89352.4]
  wire  _T_1206; // @[implicits.scala 55:10:@89353.4]
  wire  _T_1207; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:194:@89354.4]
  wire  x1326_x912_D21; // @[package.scala 96:25:@89339.4 package.scala 96:25:@89340.4]
  wire  _T_1208; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:283:@89355.4]
  wire  _T_1209; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:292:@89356.4]
  wire [31:0] x916_rdcol_number; // @[Math.scala 154:22:@89375.4 Math.scala 155:14:@89376.4]
  wire [31:0] _T_1224; // @[Math.scala 465:37:@89381.4]
  wire  x917; // @[package.scala 96:25:@89389.4 package.scala 96:25:@89390.4]
  wire  x918; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 521:60:@89393.4]
  wire  _T_1267; // @[package.scala 96:25:@89459.4 package.scala 96:25:@89460.4]
  wire  _T_1269; // @[implicits.scala 55:10:@89461.4]
  wire  _T_1270; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:194:@89462.4]
  wire  x1328_x919_D20; // @[package.scala 96:25:@89447.4 package.scala 96:25:@89448.4]
  wire  _T_1271; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:283:@89463.4]
  wire  _T_1272; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:292:@89464.4]
  wire [31:0] x925_rdcol_number; // @[Math.scala 154:22:@89485.4 Math.scala 155:14:@89486.4]
  wire [31:0] _T_1289; // @[Math.scala 465:37:@89491.4]
  wire  x926; // @[package.scala 96:25:@89499.4 package.scala 96:25:@89500.4]
  wire  x927; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 554:60:@89503.4]
  wire  _T_1332; // @[package.scala 96:25:@89569.4 package.scala 96:25:@89570.4]
  wire  _T_1334; // @[implicits.scala 55:10:@89571.4]
  wire  _T_1335; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 571:194:@89572.4]
  wire  x1330_x928_D20; // @[package.scala 96:25:@89557.4 package.scala 96:25:@89558.4]
  wire  _T_1336; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 571:283:@89573.4]
  wire  _T_1337; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 571:292:@89574.4]
  wire [31:0] x934_rdrow_number; // @[Math.scala 195:22:@89593.4 Math.scala 196:14:@89594.4]
  wire [31:0] _T_1354; // @[Math.scala 406:49:@89600.4]
  wire [31:0] _T_1356; // @[Math.scala 406:56:@89602.4]
  wire [31:0] _T_1357; // @[Math.scala 406:56:@89603.4]
  wire [31:0] _T_1361; // @[package.scala 96:25:@89611.4]
  wire [31:0] x1241_number; // @[implicits.scala 133:21:@89613.4]
  wire  x936; // @[package.scala 96:25:@89627.4 package.scala 96:25:@89628.4]
  wire  x937; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 581:24:@89631.4]
  wire [31:0] _T_1384; // @[Math.scala 406:49:@89640.4]
  wire [31:0] _T_1386; // @[Math.scala 406:56:@89642.4]
  wire [31:0] _T_1387; // @[Math.scala 406:56:@89643.4]
  wire  _T_1392; // @[FixedPoint.scala 50:25:@89649.4]
  wire [1:0] _T_1396; // @[Bitwise.scala 72:12:@89651.4]
  wire [29:0] _T_1397; // @[FixedPoint.scala 18:52:@89652.4]
  wire [31:0] x940_number; // @[Cat.scala 30:58:@89653.4]
  wire [38:0] _GEN_4; // @[Math.scala 450:32:@89658.4]
  wire [38:0] _T_1402; // @[Math.scala 450:32:@89658.4]
  wire [37:0] _GEN_5; // @[Math.scala 450:32:@89663.4]
  wire [37:0] _T_1406; // @[Math.scala 450:32:@89663.4]
  wire  _T_1433; // @[package.scala 96:25:@89722.4 package.scala 96:25:@89723.4]
  wire  _T_1435; // @[implicits.scala 55:10:@89724.4]
  wire  _T_1436; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:194:@89725.4]
  wire  x1333_x938_D20; // @[package.scala 96:25:@89710.4 package.scala 96:25:@89711.4]
  wire  _T_1437; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:283:@89726.4]
  wire  _T_1438; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:292:@89727.4]
  wire  x945; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 610:24:@89738.4]
  wire  _T_1462; // @[package.scala 96:25:@89771.4 package.scala 96:25:@89772.4]
  wire  _T_1464; // @[implicits.scala 55:10:@89773.4]
  wire  _T_1465; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:194:@89774.4]
  wire  x1334_x946_D20; // @[package.scala 96:25:@89759.4 package.scala 96:25:@89760.4]
  wire  _T_1466; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:283:@89775.4]
  wire  _T_1467; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:292:@89776.4]
  wire  x950; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 625:24:@89787.4]
  wire  _T_1491; // @[package.scala 96:25:@89820.4 package.scala 96:25:@89821.4]
  wire  _T_1493; // @[implicits.scala 55:10:@89822.4]
  wire  _T_1494; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:194:@89823.4]
  wire  x1335_x951_D20; // @[package.scala 96:25:@89808.4 package.scala 96:25:@89809.4]
  wire  _T_1495; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:283:@89824.4]
  wire  _T_1496; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:292:@89825.4]
  wire  x955; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 640:24:@89836.4]
  wire  _T_1520; // @[package.scala 96:25:@89869.4 package.scala 96:25:@89870.4]
  wire  _T_1522; // @[implicits.scala 55:10:@89871.4]
  wire  _T_1523; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:194:@89872.4]
  wire  x1336_x956_D20; // @[package.scala 96:25:@89857.4 package.scala 96:25:@89858.4]
  wire  _T_1524; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:283:@89873.4]
  wire  _T_1525; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:292:@89874.4]
  wire  x960; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 655:24:@89885.4]
  wire  _T_1551; // @[package.scala 96:25:@89920.4 package.scala 96:25:@89921.4]
  wire  _T_1553; // @[implicits.scala 55:10:@89922.4]
  wire  _T_1554; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:194:@89923.4]
  wire  x1337_x961_D20; // @[package.scala 96:25:@89908.4 package.scala 96:25:@89909.4]
  wire  _T_1555; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:283:@89924.4]
  wire  _T_1556; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:292:@89925.4]
  wire  x965; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 678:59:@89936.4]
  wire  _T_1580; // @[package.scala 96:25:@89969.4 package.scala 96:25:@89970.4]
  wire  _T_1582; // @[implicits.scala 55:10:@89971.4]
  wire  _T_1583; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:194:@89972.4]
  wire  x1338_x966_D20; // @[package.scala 96:25:@89957.4 package.scala 96:25:@89958.4]
  wire  _T_1584; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:283:@89973.4]
  wire  _T_1585; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:292:@89974.4]
  wire  x970; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 693:59:@89985.4]
  wire  _T_1609; // @[package.scala 96:25:@90018.4 package.scala 96:25:@90019.4]
  wire  _T_1611; // @[implicits.scala 55:10:@90020.4]
  wire  _T_1612; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:194:@90021.4]
  wire  x1339_x971_D20; // @[package.scala 96:25:@90006.4 package.scala 96:25:@90007.4]
  wire  _T_1613; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:283:@90022.4]
  wire  _T_1614; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:292:@90023.4]
  wire  x1340_x910_D1; // @[package.scala 96:25:@90039.4 package.scala 96:25:@90040.4]
  wire  x975; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 710:59:@90043.4]
  wire  _T_1647; // @[package.scala 96:25:@90094.4 package.scala 96:25:@90095.4]
  wire  _T_1649; // @[implicits.scala 55:10:@90096.4]
  wire  _T_1650; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:194:@90097.4]
  wire  x1343_x976_D20; // @[package.scala 96:25:@90082.4 package.scala 96:25:@90083.4]
  wire  _T_1651; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:283:@90098.4]
  wire  _T_1652; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:292:@90099.4]
  wire  x980; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 729:59:@90110.4]
  wire  _T_1676; // @[package.scala 96:25:@90143.4 package.scala 96:25:@90144.4]
  wire  _T_1678; // @[implicits.scala 55:10:@90145.4]
  wire  _T_1679; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:194:@90146.4]
  wire  x1344_x981_D20; // @[package.scala 96:25:@90131.4 package.scala 96:25:@90132.4]
  wire  _T_1680; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:283:@90147.4]
  wire  _T_1681; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:292:@90148.4]
  wire  x985; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 744:59:@90159.4]
  wire  _T_1705; // @[package.scala 96:25:@90192.4 package.scala 96:25:@90193.4]
  wire  _T_1707; // @[implicits.scala 55:10:@90194.4]
  wire  _T_1708; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:194:@90195.4]
  wire  x1345_x986_D20; // @[package.scala 96:25:@90180.4 package.scala 96:25:@90181.4]
  wire  _T_1709; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:283:@90196.4]
  wire  _T_1710; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:292:@90197.4]
  wire [31:0] x990_rdrow_number; // @[Math.scala 195:22:@90216.4 Math.scala 196:14:@90217.4]
  wire [31:0] _T_1727; // @[Math.scala 406:49:@90223.4]
  wire [31:0] _T_1729; // @[Math.scala 406:56:@90225.4]
  wire [31:0] _T_1730; // @[Math.scala 406:56:@90226.4]
  wire [31:0] _T_1734; // @[package.scala 96:25:@90234.4]
  wire [31:0] x1246_number; // @[implicits.scala 133:21:@90236.4]
  wire  x992; // @[package.scala 96:25:@90250.4 package.scala 96:25:@90251.4]
  wire  x993; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 765:24:@90254.4]
  wire [31:0] _T_1757; // @[Math.scala 406:49:@90263.4]
  wire [31:0] _T_1759; // @[Math.scala 406:56:@90265.4]
  wire [31:0] _T_1760; // @[Math.scala 406:56:@90266.4]
  wire  _T_1765; // @[FixedPoint.scala 50:25:@90272.4]
  wire [1:0] _T_1769; // @[Bitwise.scala 72:12:@90274.4]
  wire [29:0] _T_1770; // @[FixedPoint.scala 18:52:@90275.4]
  wire [31:0] x996_number; // @[Cat.scala 30:58:@90276.4]
  wire [38:0] _GEN_6; // @[Math.scala 450:32:@90281.4]
  wire [38:0] _T_1775; // @[Math.scala 450:32:@90281.4]
  wire [37:0] _GEN_7; // @[Math.scala 450:32:@90286.4]
  wire [37:0] _T_1779; // @[Math.scala 450:32:@90286.4]
  wire  _T_1808; // @[package.scala 96:25:@90347.4 package.scala 96:25:@90348.4]
  wire  _T_1810; // @[implicits.scala 55:10:@90349.4]
  wire  _T_1811; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 798:194:@90350.4]
  wire  x1347_x994_D20; // @[package.scala 96:25:@90326.4 package.scala 96:25:@90327.4]
  wire  _T_1812; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 798:283:@90351.4]
  wire  _T_1813; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 798:292:@90352.4]
  wire  x1001; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 802:60:@90363.4]
  wire  _T_1837; // @[package.scala 96:25:@90396.4 package.scala 96:25:@90397.4]
  wire  _T_1839; // @[implicits.scala 55:10:@90398.4]
  wire  _T_1840; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:199:@90399.4]
  wire  x1349_x1002_D20; // @[package.scala 96:25:@90384.4 package.scala 96:25:@90385.4]
  wire  _T_1841; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:288:@90400.4]
  wire  _T_1842; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:297:@90401.4]
  wire  x1006; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 817:60:@90412.4]
  wire  _T_1866; // @[package.scala 96:25:@90445.4 package.scala 96:25:@90446.4]
  wire  _T_1868; // @[implicits.scala 55:10:@90447.4]
  wire  _T_1869; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:199:@90448.4]
  wire  x1350_x1007_D20; // @[package.scala 96:25:@90433.4 package.scala 96:25:@90434.4]
  wire  _T_1870; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:288:@90449.4]
  wire  _T_1871; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:297:@90450.4]
  wire  x1011; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 832:60:@90461.4]
  wire  _T_1895; // @[package.scala 96:25:@90494.4 package.scala 96:25:@90495.4]
  wire  _T_1897; // @[implicits.scala 55:10:@90496.4]
  wire  _T_1898; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:199:@90497.4]
  wire  x1351_x1012_D20; // @[package.scala 96:25:@90482.4 package.scala 96:25:@90483.4]
  wire  _T_1899; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:288:@90498.4]
  wire  _T_1900; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:297:@90499.4]
  wire  x1016; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 847:60:@90510.4]
  wire  _T_1924; // @[package.scala 96:25:@90543.4 package.scala 96:25:@90544.4]
  wire  _T_1926; // @[implicits.scala 55:10:@90545.4]
  wire  _T_1927; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:199:@90546.4]
  wire  x1352_x1017_D20; // @[package.scala 96:25:@90531.4 package.scala 96:25:@90532.4]
  wire  _T_1928; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:288:@90547.4]
  wire  _T_1929; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:297:@90548.4]
  wire  x1021; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 862:60:@90559.4]
  wire  _T_1953; // @[package.scala 96:25:@90592.4 package.scala 96:25:@90593.4]
  wire  _T_1955; // @[implicits.scala 55:10:@90594.4]
  wire  _T_1956; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:199:@90595.4]
  wire  x1353_x1022_D20; // @[package.scala 96:25:@90580.4 package.scala 96:25:@90581.4]
  wire  _T_1957; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:288:@90596.4]
  wire  _T_1958; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:297:@90597.4]
  wire  x1026; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 877:60:@90608.4]
  wire  _T_1982; // @[package.scala 96:25:@90641.4 package.scala 96:25:@90642.4]
  wire  _T_1984; // @[implicits.scala 55:10:@90643.4]
  wire  _T_1985; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:199:@90644.4]
  wire  x1354_x1027_D20; // @[package.scala 96:25:@90629.4 package.scala 96:25:@90630.4]
  wire  _T_1986; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:288:@90645.4]
  wire  _T_1987; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:297:@90646.4]
  wire  x1031; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 892:60:@90657.4]
  wire  _T_2017; // @[package.scala 96:25:@90708.4 package.scala 96:25:@90709.4]
  wire  _T_2019; // @[implicits.scala 55:10:@90710.4]
  wire  _T_2020; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:199:@90711.4]
  wire  x1356_x1032_D20; // @[package.scala 96:25:@90687.4 package.scala 96:25:@90688.4]
  wire  _T_2021; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:288:@90712.4]
  wire  _T_2022; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:297:@90713.4]
  wire  x1036; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 917:60:@90724.4]
  wire  _T_2048; // @[package.scala 96:25:@90759.4 package.scala 96:25:@90760.4]
  wire  _T_2050; // @[implicits.scala 55:10:@90761.4]
  wire  _T_2051; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:199:@90762.4]
  wire  x1358_x1037_D20; // @[package.scala 96:25:@90747.4 package.scala 96:25:@90748.4]
  wire  _T_2052; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:288:@90763.4]
  wire  _T_2053; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:297:@90764.4]
  wire  x1041; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 934:60:@90775.4]
  wire  _T_2077; // @[package.scala 96:25:@90808.4 package.scala 96:25:@90809.4]
  wire  _T_2079; // @[implicits.scala 55:10:@90810.4]
  wire  _T_2080; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 945:199:@90811.4]
  wire  x1359_x1042_D20; // @[package.scala 96:25:@90796.4 package.scala 96:25:@90797.4]
  wire  _T_2081; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 945:288:@90812.4]
  wire  _T_2082; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 945:297:@90813.4]
  wire [7:0] x878_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 359:29:@88782.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:341:@88803.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@90825.4]
  wire [7:0] x943_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 602:29:@89713.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:411:@89734.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@90837.4]
  wire [7:0] x948_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 617:29:@89762.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:411:@89783.4]
  wire [9:0] _GEN_10; // @[Math.scala 450:32:@90849.4]
  wire [7:0] x953_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 632:29:@89811.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:411:@89832.4]
  wire [8:0] _GEN_11; // @[Math.scala 450:32:@90861.4]
  wire [7:0] x1004_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 809:30:@90387.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:416:@90408.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@90873.4]
  wire [7:0] x1058_sum_number; // @[Math.scala 154:22:@90996.4 Math.scala 155:14:@90997.4]
  wire [3:0] _T_2159; // @[FixedPoint.scala 18:52:@91002.4]
  wire [7:0] x884_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 382:29:@88872.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:341:@88893.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@91008.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@91020.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@91032.4]
  wire [7:0] x958_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 647:29:@89860.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:411:@89881.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@91044.4]
  wire [7:0] x1009_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 824:30:@90436.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:416:@90457.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@91056.4]
  wire [7:0] x1072_sum_number; // @[Math.scala 154:22:@91179.4 Math.scala 155:14:@91180.4]
  wire [3:0] _T_2235; // @[FixedPoint.scala 18:52:@91185.4]
  wire [7:0] x890_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 405:29:@88962.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:341:@88983.4]
  wire [8:0] _GEN_18; // @[Math.scala 450:32:@91191.4]
  wire [9:0] _GEN_19; // @[Math.scala 450:32:@91205.4]
  wire [7:0] x963_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 670:29:@89911.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:411:@89932.4]
  wire [8:0] _GEN_20; // @[Math.scala 450:32:@91217.4]
  wire [7:0] x1014_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 839:30:@90485.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:416:@90506.4]
  wire [8:0] _GEN_21; // @[Math.scala 450:32:@91229.4]
  wire [7:0] x1085_sum_number; // @[Math.scala 154:22:@91334.4 Math.scala 155:14:@91335.4]
  wire [3:0] _T_2301; // @[FixedPoint.scala 18:52:@91340.4]
  wire [7:0] x896_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 436:29:@89054.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:411:@89075.4]
  wire [8:0] _GEN_22; // @[Math.scala 450:32:@91346.4]
  wire [9:0] _GEN_23; // @[Math.scala 450:32:@91358.4]
  wire [7:0] x968_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 685:29:@89960.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:411:@89981.4]
  wire [8:0] _GEN_24; // @[Math.scala 450:32:@91370.4]
  wire [7:0] x1019_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 854:30:@90534.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:416:@90555.4]
  wire [8:0] _GEN_25; // @[Math.scala 450:32:@91382.4]
  wire [7:0] x1098_sum_number; // @[Math.scala 154:22:@91487.4 Math.scala 155:14:@91488.4]
  wire [3:0] _T_2365; // @[FixedPoint.scala 18:52:@91493.4]
  wire [7:0] x902_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 459:29:@89144.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:411:@89165.4]
  wire [8:0] _GEN_26; // @[Math.scala 450:32:@91499.4]
  wire [9:0] _GEN_27; // @[Math.scala 450:32:@91511.4]
  wire [7:0] x973_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 700:29:@90009.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:411:@90030.4]
  wire [8:0] _GEN_28; // @[Math.scala 450:32:@91523.4]
  wire [7:0] x1024_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 869:30:@90583.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:416:@90604.4]
  wire [8:0] _GEN_29; // @[Math.scala 450:32:@91535.4]
  wire [7:0] x1111_sum_number; // @[Math.scala 154:22:@91640.4 Math.scala 155:14:@91641.4]
  wire [3:0] _T_2429; // @[FixedPoint.scala 18:52:@91646.4]
  wire [7:0] x908_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 482:29:@89234.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:411:@89255.4]
  wire [8:0] _GEN_30; // @[Math.scala 450:32:@91652.4]
  wire [9:0] _GEN_31; // @[Math.scala 450:32:@91664.4]
  wire [7:0] x978_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 721:29:@90085.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:411:@90106.4]
  wire [8:0] _GEN_32; // @[Math.scala 450:32:@91676.4]
  wire [7:0] x1029_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 884:30:@90632.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:416:@90653.4]
  wire [8:0] _GEN_33; // @[Math.scala 450:32:@91688.4]
  wire [7:0] x1124_sum_number; // @[Math.scala 154:22:@91795.4 Math.scala 155:14:@91796.4]
  wire [3:0] _T_2495; // @[FixedPoint.scala 18:52:@91801.4]
  wire [7:0] x914_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 509:29:@89342.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:411:@89363.4]
  wire [8:0] _GEN_34; // @[Math.scala 450:32:@91807.4]
  wire [9:0] _GEN_35; // @[Math.scala 450:32:@91819.4]
  wire [7:0] x983_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 736:29:@90134.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:411:@90155.4]
  wire [8:0] _GEN_36; // @[Math.scala 450:32:@91831.4]
  wire [7:0] x1034_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 903:30:@90699.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:416:@90720.4]
  wire [8:0] _GEN_37; // @[Math.scala 450:32:@91843.4]
  wire [7:0] x1137_sum_number; // @[Math.scala 154:22:@91948.4 Math.scala 155:14:@91949.4]
  wire [3:0] _T_2559; // @[FixedPoint.scala 18:52:@91954.4]
  wire [7:0] x923_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 540:29:@89450.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:411:@89471.4]
  wire [8:0] _GEN_38; // @[Math.scala 450:32:@91960.4]
  wire [9:0] _GEN_39; // @[Math.scala 450:32:@91972.4]
  wire [7:0] x988_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 751:29:@90183.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:411:@90204.4]
  wire [8:0] _GEN_40; // @[Math.scala 450:32:@91984.4]
  wire [7:0] x1039_rd_0_number; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 926:30:@90750.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:416:@90771.4]
  wire [8:0] _GEN_41; // @[Math.scala 450:32:@91996.4]
  wire [7:0] x1150_sum_number; // @[Math.scala 154:22:@92101.4 Math.scala 155:14:@92102.4]
  wire [3:0] _T_2623; // @[FixedPoint.scala 18:52:@92107.4]
  wire [31:0] _T_2642; // @[Cat.scala 30:58:@92123.4]
  wire [31:0] _T_2645; // @[Cat.scala 30:58:@92126.4]
  wire  _T_2658; // @[package.scala 96:25:@92162.4 package.scala 96:25:@92163.4]
  wire  _T_2660; // @[implicits.scala 55:10:@92164.4]
  wire  x1380_b801_D59; // @[package.scala 96:25:@92144.4 package.scala 96:25:@92145.4]
  wire  _T_2661; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1225:117:@92165.4]
  wire  x1381_b802_D59; // @[package.scala 96:25:@92153.4 package.scala 96:25:@92154.4]
  wire  _T_2662; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1225:124:@92166.4]
  wire [31:0] x1259_x814_D12_number; // @[package.scala 96:25:@87728.4 package.scala 96:25:@87729.4]
  wire [31:0] x1261_x1232_D26_number; // @[package.scala 96:25:@87746.4 package.scala 96:25:@87747.4]
  wire [31:0] x1263_x818_sum_D7_number; // @[package.scala 96:25:@87764.4 package.scala 96:25:@87765.4]
  wire [31:0] x1267_x824_sum_D6_number; // @[package.scala 96:25:@87871.4 package.scala 96:25:@87872.4]
  wire [31:0] x1268_x822_D11_number; // @[package.scala 96:25:@87880.4 package.scala 96:25:@87881.4]
  wire [31:0] x1269_x830_sum_D6_number; // @[package.scala 96:25:@87960.4 package.scala 96:25:@87961.4]
  wire [31:0] x1271_x828_D11_number; // @[package.scala 96:25:@87978.4 package.scala 96:25:@87979.4]
  wire [31:0] x1272_x834_D11_number; // @[package.scala 96:25:@88060.4 package.scala 96:25:@88061.4]
  wire [31:0] x1273_x836_sum_D6_number; // @[package.scala 96:25:@88069.4 package.scala 96:25:@88070.4]
  wire [31:0] x1275_x842_sum_D6_number; // @[package.scala 96:25:@88158.4 package.scala 96:25:@88159.4]
  wire [31:0] x1276_x840_D11_number; // @[package.scala 96:25:@88167.4 package.scala 96:25:@88168.4]
  wire [31:0] x1278_x846_D11_number; // @[package.scala 96:25:@88256.4 package.scala 96:25:@88257.4]
  wire [31:0] x1279_x848_sum_D6_number; // @[package.scala 96:25:@88265.4 package.scala 96:25:@88266.4]
  wire [31:0] x1281_x852_D11_number; // @[package.scala 96:25:@88354.4 package.scala 96:25:@88355.4]
  wire [31:0] x1283_x854_sum_D6_number; // @[package.scala 96:25:@88372.4 package.scala 96:25:@88373.4]
  wire [31:0] x1285_x858_D11_number; // @[package.scala 96:25:@88461.4 package.scala 96:25:@88462.4]
  wire [31:0] x1286_x860_sum_D6_number; // @[package.scala 96:25:@88470.4 package.scala 96:25:@88471.4]
  wire [31:0] x871_sum_number; // @[Math.scala 154:22:@88644.4 Math.scala 155:14:@88645.4]
  wire [31:0] x1292_x1237_D21_number; // @[package.scala 96:25:@88653.4 package.scala 96:25:@88654.4]
  wire [31:0] x1294_x858_D35_number; // @[package.scala 96:25:@88671.4 package.scala 96:25:@88672.4]
  wire [31:0] x877_sum_number; // @[Math.scala 154:22:@88761.4 Math.scala 155:14:@88762.4]
  wire [31:0] x1299_x852_D35_number; // @[package.scala 96:25:@88770.4 package.scala 96:25:@88771.4]
  wire [31:0] x883_sum_number; // @[Math.scala 154:22:@88851.4 Math.scala 155:14:@88852.4]
  wire [31:0] x1303_x846_D35_number; // @[package.scala 96:25:@88860.4 package.scala 96:25:@88861.4]
  wire [31:0] x889_sum_number; // @[Math.scala 154:22:@88941.4 Math.scala 155:14:@88942.4]
  wire [31:0] x1308_x840_D35_number; // @[package.scala 96:25:@88959.4 package.scala 96:25:@88960.4]
  wire [31:0] x895_sum_number; // @[Math.scala 154:22:@89033.4 Math.scala 155:14:@89034.4]
  wire [31:0] x1311_x834_D35_number; // @[package.scala 96:25:@89042.4 package.scala 96:25:@89043.4]
  wire [31:0] x901_sum_number; // @[Math.scala 154:22:@89123.4 Math.scala 155:14:@89124.4]
  wire [31:0] x1316_x828_D35_number; // @[package.scala 96:25:@89141.4 package.scala 96:25:@89142.4]
  wire [31:0] x907_sum_number; // @[Math.scala 154:22:@89213.4 Math.scala 155:14:@89214.4]
  wire [31:0] x1320_x822_D35_number; // @[package.scala 96:25:@89231.4 package.scala 96:25:@89232.4]
  wire [31:0] x1324_x814_D36_number; // @[package.scala 96:25:@89321.4 package.scala 96:25:@89322.4]
  wire [31:0] x1325_x913_sum_D1_number; // @[package.scala 96:25:@89330.4 package.scala 96:25:@89331.4]
  wire [31:0] x922_sum_number; // @[Math.scala 154:22:@89429.4 Math.scala 155:14:@89430.4]
  wire [31:0] x1327_x920_D5_number; // @[package.scala 96:25:@89438.4 package.scala 96:25:@89439.4]
  wire [31:0] x931_sum_number; // @[Math.scala 154:22:@89539.4 Math.scala 155:14:@89540.4]
  wire [31:0] x1329_x929_D5_number; // @[package.scala 96:25:@89548.4 package.scala 96:25:@89549.4]
  wire [31:0] x942_sum_number; // @[Math.scala 154:22:@89692.4 Math.scala 155:14:@89693.4]
  wire [31:0] x1332_x1242_D20_number; // @[package.scala 96:25:@89701.4 package.scala 96:25:@89702.4]
  wire [31:0] x947_sum_number; // @[Math.scala 154:22:@89750.4 Math.scala 155:14:@89751.4]
  wire [31:0] x952_sum_number; // @[Math.scala 154:22:@89799.4 Math.scala 155:14:@89800.4]
  wire [31:0] x957_sum_number; // @[Math.scala 154:22:@89848.4 Math.scala 155:14:@89849.4]
  wire [31:0] x962_sum_number; // @[Math.scala 154:22:@89899.4 Math.scala 155:14:@89900.4]
  wire [31:0] x967_sum_number; // @[Math.scala 154:22:@89948.4 Math.scala 155:14:@89949.4]
  wire [31:0] x972_sum_number; // @[Math.scala 154:22:@89997.4 Math.scala 155:14:@89998.4]
  wire [31:0] x1342_x977_sum_D1_number; // @[package.scala 96:25:@90073.4 package.scala 96:25:@90074.4]
  wire [31:0] x982_sum_number; // @[Math.scala 154:22:@90122.4 Math.scala 155:14:@90123.4]
  wire [31:0] x987_sum_number; // @[Math.scala 154:22:@90171.4 Math.scala 155:14:@90172.4]
  wire [31:0] x998_sum_number; // @[Math.scala 154:22:@90317.4 Math.scala 155:14:@90318.4]
  wire [31:0] x1348_x1247_D20_number; // @[package.scala 96:25:@90335.4 package.scala 96:25:@90336.4]
  wire [31:0] x1003_sum_number; // @[Math.scala 154:22:@90375.4 Math.scala 155:14:@90376.4]
  wire [31:0] x1008_sum_number; // @[Math.scala 154:22:@90424.4 Math.scala 155:14:@90425.4]
  wire [31:0] x1013_sum_number; // @[Math.scala 154:22:@90473.4 Math.scala 155:14:@90474.4]
  wire [31:0] x1018_sum_number; // @[Math.scala 154:22:@90522.4 Math.scala 155:14:@90523.4]
  wire [31:0] x1023_sum_number; // @[Math.scala 154:22:@90571.4 Math.scala 155:14:@90572.4]
  wire [31:0] x1028_sum_number; // @[Math.scala 154:22:@90620.4 Math.scala 155:14:@90621.4]
  wire [31:0] x1357_x1033_sum_D1_number; // @[package.scala 96:25:@90696.4 package.scala 96:25:@90697.4]
  wire [31:0] x1038_sum_number; // @[Math.scala 154:22:@90738.4 Math.scala 155:14:@90739.4]
  wire [31:0] x1043_sum_number; // @[Math.scala 154:22:@90787.4 Math.scala 155:14:@90788.4]
  wire [8:0] _T_2090; // @[package.scala 96:25:@90831.4 package.scala 96:25:@90832.4]
  wire [8:0] _T_2096; // @[package.scala 96:25:@90843.4 package.scala 96:25:@90844.4]
  wire [9:0] _T_2102; // @[package.scala 96:25:@90855.4 package.scala 96:25:@90856.4]
  wire [8:0] _T_2108; // @[package.scala 96:25:@90867.4 package.scala 96:25:@90868.4]
  wire [8:0] _T_2114; // @[package.scala 96:25:@90879.4 package.scala 96:25:@90880.4]
  wire [8:0] _T_2166; // @[package.scala 96:25:@91014.4 package.scala 96:25:@91015.4]
  wire [8:0] _T_2172; // @[package.scala 96:25:@91026.4 package.scala 96:25:@91027.4]
  wire [9:0] _T_2178; // @[package.scala 96:25:@91038.4 package.scala 96:25:@91039.4]
  wire [8:0] _T_2184; // @[package.scala 96:25:@91050.4 package.scala 96:25:@91051.4]
  wire [8:0] _T_2190; // @[package.scala 96:25:@91062.4 package.scala 96:25:@91063.4]
  wire [8:0] _T_2242; // @[package.scala 96:25:@91197.4 package.scala 96:25:@91198.4]
  wire [9:0] _T_2250; // @[package.scala 96:25:@91211.4 package.scala 96:25:@91212.4]
  wire [8:0] _T_2256; // @[package.scala 96:25:@91223.4 package.scala 96:25:@91224.4]
  wire [8:0] _T_2262; // @[package.scala 96:25:@91235.4 package.scala 96:25:@91236.4]
  wire [8:0] _T_2308; // @[package.scala 96:25:@91352.4 package.scala 96:25:@91353.4]
  wire [9:0] _T_2314; // @[package.scala 96:25:@91364.4 package.scala 96:25:@91365.4]
  wire [8:0] _T_2320; // @[package.scala 96:25:@91376.4 package.scala 96:25:@91377.4]
  wire [8:0] _T_2326; // @[package.scala 96:25:@91388.4 package.scala 96:25:@91389.4]
  wire [8:0] _T_2372; // @[package.scala 96:25:@91505.4 package.scala 96:25:@91506.4]
  wire [9:0] _T_2378; // @[package.scala 96:25:@91517.4 package.scala 96:25:@91518.4]
  wire [8:0] _T_2384; // @[package.scala 96:25:@91529.4 package.scala 96:25:@91530.4]
  wire [8:0] _T_2390; // @[package.scala 96:25:@91541.4 package.scala 96:25:@91542.4]
  wire [8:0] _T_2436; // @[package.scala 96:25:@91658.4 package.scala 96:25:@91659.4]
  wire [9:0] _T_2442; // @[package.scala 96:25:@91670.4 package.scala 96:25:@91671.4]
  wire [8:0] _T_2448; // @[package.scala 96:25:@91682.4 package.scala 96:25:@91683.4]
  wire [8:0] _T_2454; // @[package.scala 96:25:@91694.4 package.scala 96:25:@91695.4]
  wire [8:0] _T_2502; // @[package.scala 96:25:@91813.4 package.scala 96:25:@91814.4]
  wire [9:0] _T_2508; // @[package.scala 96:25:@91825.4 package.scala 96:25:@91826.4]
  wire [8:0] _T_2514; // @[package.scala 96:25:@91837.4 package.scala 96:25:@91838.4]
  wire [8:0] _T_2520; // @[package.scala 96:25:@91849.4 package.scala 96:25:@91850.4]
  wire [8:0] _T_2566; // @[package.scala 96:25:@91966.4 package.scala 96:25:@91967.4]
  wire [9:0] _T_2572; // @[package.scala 96:25:@91978.4 package.scala 96:25:@91979.4]
  wire [8:0] _T_2578; // @[package.scala 96:25:@91990.4 package.scala 96:25:@91991.4]
  wire [8:0] _T_2584; // @[package.scala 96:25:@92002.4 package.scala 96:25:@92003.4]
  _ _ ( // @[Math.scala 709:24:@87268.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@87280.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_64 RetimeWrapper ( // @[package.scala 93:22:@87303.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x805_lb_0 x805_lb_0 ( // @[m_x805_lb_0.scala 63:17:@87313.4]
    .clock(x805_lb_0_clock),
    .reset(x805_lb_0_reset),
    .io_rPort_29_banks_1(x805_lb_0_io_rPort_29_banks_1),
    .io_rPort_29_banks_0(x805_lb_0_io_rPort_29_banks_0),
    .io_rPort_29_ofs_0(x805_lb_0_io_rPort_29_ofs_0),
    .io_rPort_29_en_0(x805_lb_0_io_rPort_29_en_0),
    .io_rPort_29_backpressure(x805_lb_0_io_rPort_29_backpressure),
    .io_rPort_29_output_0(x805_lb_0_io_rPort_29_output_0),
    .io_rPort_28_banks_1(x805_lb_0_io_rPort_28_banks_1),
    .io_rPort_28_banks_0(x805_lb_0_io_rPort_28_banks_0),
    .io_rPort_28_ofs_0(x805_lb_0_io_rPort_28_ofs_0),
    .io_rPort_28_en_0(x805_lb_0_io_rPort_28_en_0),
    .io_rPort_28_backpressure(x805_lb_0_io_rPort_28_backpressure),
    .io_rPort_28_output_0(x805_lb_0_io_rPort_28_output_0),
    .io_rPort_27_banks_1(x805_lb_0_io_rPort_27_banks_1),
    .io_rPort_27_banks_0(x805_lb_0_io_rPort_27_banks_0),
    .io_rPort_27_ofs_0(x805_lb_0_io_rPort_27_ofs_0),
    .io_rPort_27_en_0(x805_lb_0_io_rPort_27_en_0),
    .io_rPort_27_backpressure(x805_lb_0_io_rPort_27_backpressure),
    .io_rPort_27_output_0(x805_lb_0_io_rPort_27_output_0),
    .io_rPort_26_banks_1(x805_lb_0_io_rPort_26_banks_1),
    .io_rPort_26_banks_0(x805_lb_0_io_rPort_26_banks_0),
    .io_rPort_26_ofs_0(x805_lb_0_io_rPort_26_ofs_0),
    .io_rPort_26_en_0(x805_lb_0_io_rPort_26_en_0),
    .io_rPort_26_backpressure(x805_lb_0_io_rPort_26_backpressure),
    .io_rPort_26_output_0(x805_lb_0_io_rPort_26_output_0),
    .io_rPort_25_banks_1(x805_lb_0_io_rPort_25_banks_1),
    .io_rPort_25_banks_0(x805_lb_0_io_rPort_25_banks_0),
    .io_rPort_25_ofs_0(x805_lb_0_io_rPort_25_ofs_0),
    .io_rPort_25_en_0(x805_lb_0_io_rPort_25_en_0),
    .io_rPort_25_backpressure(x805_lb_0_io_rPort_25_backpressure),
    .io_rPort_25_output_0(x805_lb_0_io_rPort_25_output_0),
    .io_rPort_24_banks_1(x805_lb_0_io_rPort_24_banks_1),
    .io_rPort_24_banks_0(x805_lb_0_io_rPort_24_banks_0),
    .io_rPort_24_ofs_0(x805_lb_0_io_rPort_24_ofs_0),
    .io_rPort_24_en_0(x805_lb_0_io_rPort_24_en_0),
    .io_rPort_24_backpressure(x805_lb_0_io_rPort_24_backpressure),
    .io_rPort_24_output_0(x805_lb_0_io_rPort_24_output_0),
    .io_rPort_23_banks_1(x805_lb_0_io_rPort_23_banks_1),
    .io_rPort_23_banks_0(x805_lb_0_io_rPort_23_banks_0),
    .io_rPort_23_ofs_0(x805_lb_0_io_rPort_23_ofs_0),
    .io_rPort_23_en_0(x805_lb_0_io_rPort_23_en_0),
    .io_rPort_23_backpressure(x805_lb_0_io_rPort_23_backpressure),
    .io_rPort_23_output_0(x805_lb_0_io_rPort_23_output_0),
    .io_rPort_22_banks_1(x805_lb_0_io_rPort_22_banks_1),
    .io_rPort_22_banks_0(x805_lb_0_io_rPort_22_banks_0),
    .io_rPort_22_ofs_0(x805_lb_0_io_rPort_22_ofs_0),
    .io_rPort_22_en_0(x805_lb_0_io_rPort_22_en_0),
    .io_rPort_22_backpressure(x805_lb_0_io_rPort_22_backpressure),
    .io_rPort_22_output_0(x805_lb_0_io_rPort_22_output_0),
    .io_rPort_21_banks_1(x805_lb_0_io_rPort_21_banks_1),
    .io_rPort_21_banks_0(x805_lb_0_io_rPort_21_banks_0),
    .io_rPort_21_ofs_0(x805_lb_0_io_rPort_21_ofs_0),
    .io_rPort_21_en_0(x805_lb_0_io_rPort_21_en_0),
    .io_rPort_21_backpressure(x805_lb_0_io_rPort_21_backpressure),
    .io_rPort_21_output_0(x805_lb_0_io_rPort_21_output_0),
    .io_rPort_20_banks_1(x805_lb_0_io_rPort_20_banks_1),
    .io_rPort_20_banks_0(x805_lb_0_io_rPort_20_banks_0),
    .io_rPort_20_ofs_0(x805_lb_0_io_rPort_20_ofs_0),
    .io_rPort_20_en_0(x805_lb_0_io_rPort_20_en_0),
    .io_rPort_20_backpressure(x805_lb_0_io_rPort_20_backpressure),
    .io_rPort_20_output_0(x805_lb_0_io_rPort_20_output_0),
    .io_rPort_19_banks_1(x805_lb_0_io_rPort_19_banks_1),
    .io_rPort_19_banks_0(x805_lb_0_io_rPort_19_banks_0),
    .io_rPort_19_ofs_0(x805_lb_0_io_rPort_19_ofs_0),
    .io_rPort_19_en_0(x805_lb_0_io_rPort_19_en_0),
    .io_rPort_19_backpressure(x805_lb_0_io_rPort_19_backpressure),
    .io_rPort_19_output_0(x805_lb_0_io_rPort_19_output_0),
    .io_rPort_18_banks_1(x805_lb_0_io_rPort_18_banks_1),
    .io_rPort_18_banks_0(x805_lb_0_io_rPort_18_banks_0),
    .io_rPort_18_ofs_0(x805_lb_0_io_rPort_18_ofs_0),
    .io_rPort_18_en_0(x805_lb_0_io_rPort_18_en_0),
    .io_rPort_18_backpressure(x805_lb_0_io_rPort_18_backpressure),
    .io_rPort_18_output_0(x805_lb_0_io_rPort_18_output_0),
    .io_rPort_17_banks_1(x805_lb_0_io_rPort_17_banks_1),
    .io_rPort_17_banks_0(x805_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x805_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x805_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x805_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x805_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_1(x805_lb_0_io_rPort_16_banks_1),
    .io_rPort_16_banks_0(x805_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x805_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x805_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x805_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x805_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_1(x805_lb_0_io_rPort_15_banks_1),
    .io_rPort_15_banks_0(x805_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x805_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x805_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x805_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x805_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_1(x805_lb_0_io_rPort_14_banks_1),
    .io_rPort_14_banks_0(x805_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x805_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x805_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x805_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x805_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_1(x805_lb_0_io_rPort_13_banks_1),
    .io_rPort_13_banks_0(x805_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x805_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x805_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x805_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x805_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_1(x805_lb_0_io_rPort_12_banks_1),
    .io_rPort_12_banks_0(x805_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x805_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x805_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x805_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x805_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_1(x805_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x805_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x805_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x805_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x805_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x805_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x805_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x805_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x805_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x805_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x805_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x805_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x805_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x805_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x805_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x805_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x805_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x805_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x805_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x805_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x805_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x805_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x805_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x805_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x805_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x805_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x805_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x805_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x805_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x805_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x805_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x805_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x805_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x805_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x805_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x805_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x805_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x805_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x805_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x805_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x805_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x805_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x805_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x805_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x805_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x805_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x805_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x805_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x805_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x805_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x805_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x805_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x805_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x805_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x805_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x805_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x805_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x805_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x805_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x805_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x805_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x805_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x805_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x805_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x805_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x805_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x805_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x805_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x805_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x805_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x805_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x805_lb_0_io_rPort_0_output_0),
    .io_wPort_7_banks_1(x805_lb_0_io_wPort_7_banks_1),
    .io_wPort_7_banks_0(x805_lb_0_io_wPort_7_banks_0),
    .io_wPort_7_ofs_0(x805_lb_0_io_wPort_7_ofs_0),
    .io_wPort_7_data_0(x805_lb_0_io_wPort_7_data_0),
    .io_wPort_7_en_0(x805_lb_0_io_wPort_7_en_0),
    .io_wPort_6_banks_1(x805_lb_0_io_wPort_6_banks_1),
    .io_wPort_6_banks_0(x805_lb_0_io_wPort_6_banks_0),
    .io_wPort_6_ofs_0(x805_lb_0_io_wPort_6_ofs_0),
    .io_wPort_6_data_0(x805_lb_0_io_wPort_6_data_0),
    .io_wPort_6_en_0(x805_lb_0_io_wPort_6_en_0),
    .io_wPort_5_banks_1(x805_lb_0_io_wPort_5_banks_1),
    .io_wPort_5_banks_0(x805_lb_0_io_wPort_5_banks_0),
    .io_wPort_5_ofs_0(x805_lb_0_io_wPort_5_ofs_0),
    .io_wPort_5_data_0(x805_lb_0_io_wPort_5_data_0),
    .io_wPort_5_en_0(x805_lb_0_io_wPort_5_en_0),
    .io_wPort_4_banks_1(x805_lb_0_io_wPort_4_banks_1),
    .io_wPort_4_banks_0(x805_lb_0_io_wPort_4_banks_0),
    .io_wPort_4_ofs_0(x805_lb_0_io_wPort_4_ofs_0),
    .io_wPort_4_data_0(x805_lb_0_io_wPort_4_data_0),
    .io_wPort_4_en_0(x805_lb_0_io_wPort_4_en_0),
    .io_wPort_3_banks_1(x805_lb_0_io_wPort_3_banks_1),
    .io_wPort_3_banks_0(x805_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x805_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x805_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x805_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_1(x805_lb_0_io_wPort_2_banks_1),
    .io_wPort_2_banks_0(x805_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x805_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x805_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x805_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_1(x805_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x805_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x805_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x805_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x805_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x805_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x805_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x805_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x805_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x805_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_705 RetimeWrapper_1 ( // @[package.scala 93:22:@87631.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x814 x814_1 ( // @[Math.scala 366:24:@87653.4]
    .clock(x814_1_clock),
    .reset(x814_1_reset),
    .io_a(x814_1_io_a),
    .io_flow(x814_1_io_flow),
    .io_result(x814_1_io_result)
  );
  x758_sum x1235_sum_1 ( // @[Math.scala 150:24:@87682.4]
    .clock(x1235_sum_1_clock),
    .reset(x1235_sum_1_reset),
    .io_a(x1235_sum_1_io_a),
    .io_b(x1235_sum_1_io_b),
    .io_flow(x1235_sum_1_io_flow),
    .io_result(x1235_sum_1_io_result)
  );
  x817_div x817_div_1 ( // @[Math.scala 327:24:@87694.4]
    .clock(x817_div_1_clock),
    .reset(x817_div_1_reset),
    .io_a(x817_div_1_io_a),
    .io_flow(x817_div_1_io_flow),
    .io_result(x817_div_1_io_result)
  );
  RetimeWrapper_709 RetimeWrapper_2 ( // @[package.scala 93:22:@87704.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x758_sum x818_sum_1 ( // @[Math.scala 150:24:@87713.4]
    .clock(x818_sum_1_clock),
    .reset(x818_sum_1_reset),
    .io_a(x818_sum_1_io_a),
    .io_b(x818_sum_1_io_b),
    .io_flow(x818_sum_1_io_flow),
    .io_result(x818_sum_1_io_result)
  );
  RetimeWrapper_711 RetimeWrapper_3 ( // @[package.scala 93:22:@87723.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_4 ( // @[package.scala 93:22:@87732.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_713 RetimeWrapper_5 ( // @[package.scala 93:22:@87741.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_714 RetimeWrapper_6 ( // @[package.scala 93:22:@87750.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_715 RetimeWrapper_7 ( // @[package.scala 93:22:@87759.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_8 ( // @[package.scala 93:22:@87768.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_9 ( // @[package.scala 93:22:@87779.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  x758_sum x820_rdcol_1 ( // @[Math.scala 150:24:@87802.4]
    .clock(x820_rdcol_1_clock),
    .reset(x820_rdcol_1_reset),
    .io_a(x820_rdcol_1_io_a),
    .io_b(x820_rdcol_1_io_b),
    .io_flow(x820_rdcol_1_io_flow),
    .io_result(x820_rdcol_1_io_result)
  );
  x814 x822_1 ( // @[Math.scala 366:24:@87816.4]
    .clock(x822_1_clock),
    .reset(x822_1_reset),
    .io_a(x822_1_io_a),
    .io_flow(x822_1_io_flow),
    .io_result(x822_1_io_result)
  );
  x817_div x823_div_1 ( // @[Math.scala 327:24:@87828.4]
    .clock(x823_div_1_clock),
    .reset(x823_div_1_reset),
    .io_a(x823_div_1_io_a),
    .io_flow(x823_div_1_io_flow),
    .io_result(x823_div_1_io_result)
  );
  RetimeWrapper_721 RetimeWrapper_10 ( // @[package.scala 93:22:@87838.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x758_sum x824_sum_1 ( // @[Math.scala 150:24:@87847.4]
    .clock(x824_sum_1_clock),
    .reset(x824_sum_1_reset),
    .io_a(x824_sum_1_io_a),
    .io_b(x824_sum_1_io_b),
    .io_flow(x824_sum_1_io_flow),
    .io_result(x824_sum_1_io_result)
  );
  RetimeWrapper_714 RetimeWrapper_11 ( // @[package.scala 93:22:@87857.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_724 RetimeWrapper_12 ( // @[package.scala 93:22:@87866.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_725 RetimeWrapper_13 ( // @[package.scala 93:22:@87875.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_14 ( // @[package.scala 93:22:@87886.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  x758_sum x826_rdcol_1 ( // @[Math.scala 150:24:@87909.4]
    .clock(x826_rdcol_1_clock),
    .reset(x826_rdcol_1_reset),
    .io_a(x826_rdcol_1_io_a),
    .io_b(x826_rdcol_1_io_b),
    .io_flow(x826_rdcol_1_io_flow),
    .io_result(x826_rdcol_1_io_result)
  );
  x814 x828_1 ( // @[Math.scala 366:24:@87923.4]
    .clock(x828_1_clock),
    .reset(x828_1_reset),
    .io_a(x828_1_io_a),
    .io_flow(x828_1_io_flow),
    .io_result(x828_1_io_result)
  );
  x817_div x829_div_1 ( // @[Math.scala 327:24:@87935.4]
    .clock(x829_div_1_clock),
    .reset(x829_div_1_reset),
    .io_a(x829_div_1_io_a),
    .io_flow(x829_div_1_io_flow),
    .io_result(x829_div_1_io_result)
  );
  x758_sum x830_sum_1 ( // @[Math.scala 150:24:@87945.4]
    .clock(x830_sum_1_clock),
    .reset(x830_sum_1_reset),
    .io_a(x830_sum_1_io_a),
    .io_b(x830_sum_1_io_b),
    .io_flow(x830_sum_1_io_flow),
    .io_result(x830_sum_1_io_result)
  );
  RetimeWrapper_724 RetimeWrapper_15 ( // @[package.scala 93:22:@87955.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_714 RetimeWrapper_16 ( // @[package.scala 93:22:@87964.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_725 RetimeWrapper_17 ( // @[package.scala 93:22:@87973.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_18 ( // @[package.scala 93:22:@87984.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  x758_sum x832_rdcol_1 ( // @[Math.scala 150:24:@88007.4]
    .clock(x832_rdcol_1_clock),
    .reset(x832_rdcol_1_reset),
    .io_a(x832_rdcol_1_io_a),
    .io_b(x832_rdcol_1_io_b),
    .io_flow(x832_rdcol_1_io_flow),
    .io_result(x832_rdcol_1_io_result)
  );
  x814 x834_1 ( // @[Math.scala 366:24:@88023.4]
    .clock(x834_1_clock),
    .reset(x834_1_reset),
    .io_a(x834_1_io_a),
    .io_flow(x834_1_io_flow),
    .io_result(x834_1_io_result)
  );
  x817_div x835_div_1 ( // @[Math.scala 327:24:@88035.4]
    .clock(x835_div_1_clock),
    .reset(x835_div_1_reset),
    .io_a(x835_div_1_io_a),
    .io_flow(x835_div_1_io_flow),
    .io_result(x835_div_1_io_result)
  );
  x758_sum x836_sum_1 ( // @[Math.scala 150:24:@88045.4]
    .clock(x836_sum_1_clock),
    .reset(x836_sum_1_reset),
    .io_a(x836_sum_1_io_a),
    .io_b(x836_sum_1_io_b),
    .io_flow(x836_sum_1_io_flow),
    .io_result(x836_sum_1_io_result)
  );
  RetimeWrapper_725 RetimeWrapper_19 ( // @[package.scala 93:22:@88055.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_724 RetimeWrapper_20 ( // @[package.scala 93:22:@88064.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_714 RetimeWrapper_21 ( // @[package.scala 93:22:@88073.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_22 ( // @[package.scala 93:22:@88084.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  x758_sum x838_rdcol_1 ( // @[Math.scala 150:24:@88107.4]
    .clock(x838_rdcol_1_clock),
    .reset(x838_rdcol_1_reset),
    .io_a(x838_rdcol_1_io_a),
    .io_b(x838_rdcol_1_io_b),
    .io_flow(x838_rdcol_1_io_flow),
    .io_result(x838_rdcol_1_io_result)
  );
  x814 x840_1 ( // @[Math.scala 366:24:@88121.4]
    .clock(x840_1_clock),
    .reset(x840_1_reset),
    .io_a(x840_1_io_a),
    .io_flow(x840_1_io_flow),
    .io_result(x840_1_io_result)
  );
  x817_div x841_div_1 ( // @[Math.scala 327:24:@88133.4]
    .clock(x841_div_1_clock),
    .reset(x841_div_1_reset),
    .io_a(x841_div_1_io_a),
    .io_flow(x841_div_1_io_flow),
    .io_result(x841_div_1_io_result)
  );
  x758_sum x842_sum_1 ( // @[Math.scala 150:24:@88143.4]
    .clock(x842_sum_1_clock),
    .reset(x842_sum_1_reset),
    .io_a(x842_sum_1_io_a),
    .io_b(x842_sum_1_io_b),
    .io_flow(x842_sum_1_io_flow),
    .io_result(x842_sum_1_io_result)
  );
  RetimeWrapper_724 RetimeWrapper_23 ( // @[package.scala 93:22:@88153.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_725 RetimeWrapper_24 ( // @[package.scala 93:22:@88162.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_714 RetimeWrapper_25 ( // @[package.scala 93:22:@88171.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_26 ( // @[package.scala 93:22:@88182.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  x758_sum x844_rdcol_1 ( // @[Math.scala 150:24:@88205.4]
    .clock(x844_rdcol_1_clock),
    .reset(x844_rdcol_1_reset),
    .io_a(x844_rdcol_1_io_a),
    .io_b(x844_rdcol_1_io_b),
    .io_flow(x844_rdcol_1_io_flow),
    .io_result(x844_rdcol_1_io_result)
  );
  x814 x846_1 ( // @[Math.scala 366:24:@88219.4]
    .clock(x846_1_clock),
    .reset(x846_1_reset),
    .io_a(x846_1_io_a),
    .io_flow(x846_1_io_flow),
    .io_result(x846_1_io_result)
  );
  x817_div x847_div_1 ( // @[Math.scala 327:24:@88231.4]
    .clock(x847_div_1_clock),
    .reset(x847_div_1_reset),
    .io_a(x847_div_1_io_a),
    .io_flow(x847_div_1_io_flow),
    .io_result(x847_div_1_io_result)
  );
  x758_sum x848_sum_1 ( // @[Math.scala 150:24:@88241.4]
    .clock(x848_sum_1_clock),
    .reset(x848_sum_1_reset),
    .io_a(x848_sum_1_io_a),
    .io_b(x848_sum_1_io_b),
    .io_flow(x848_sum_1_io_flow),
    .io_result(x848_sum_1_io_result)
  );
  RetimeWrapper_725 RetimeWrapper_27 ( // @[package.scala 93:22:@88251.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_724 RetimeWrapper_28 ( // @[package.scala 93:22:@88260.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_714 RetimeWrapper_29 ( // @[package.scala 93:22:@88269.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_30 ( // @[package.scala 93:22:@88280.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x758_sum x850_rdcol_1 ( // @[Math.scala 150:24:@88303.4]
    .clock(x850_rdcol_1_clock),
    .reset(x850_rdcol_1_reset),
    .io_a(x850_rdcol_1_io_a),
    .io_b(x850_rdcol_1_io_b),
    .io_flow(x850_rdcol_1_io_flow),
    .io_result(x850_rdcol_1_io_result)
  );
  x814 x852_1 ( // @[Math.scala 366:24:@88317.4]
    .clock(x852_1_clock),
    .reset(x852_1_reset),
    .io_a(x852_1_io_a),
    .io_flow(x852_1_io_flow),
    .io_result(x852_1_io_result)
  );
  x817_div x853_div_1 ( // @[Math.scala 327:24:@88329.4]
    .clock(x853_div_1_clock),
    .reset(x853_div_1_reset),
    .io_a(x853_div_1_io_a),
    .io_flow(x853_div_1_io_flow),
    .io_result(x853_div_1_io_result)
  );
  x758_sum x854_sum_1 ( // @[Math.scala 150:24:@88339.4]
    .clock(x854_sum_1_clock),
    .reset(x854_sum_1_reset),
    .io_a(x854_sum_1_io_a),
    .io_b(x854_sum_1_io_b),
    .io_flow(x854_sum_1_io_flow),
    .io_result(x854_sum_1_io_result)
  );
  RetimeWrapper_725 RetimeWrapper_31 ( // @[package.scala 93:22:@88349.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_714 RetimeWrapper_32 ( // @[package.scala 93:22:@88358.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_724 RetimeWrapper_33 ( // @[package.scala 93:22:@88367.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_34 ( // @[package.scala 93:22:@88378.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x758_sum x856_rdcol_1 ( // @[Math.scala 150:24:@88401.4]
    .clock(x856_rdcol_1_clock),
    .reset(x856_rdcol_1_reset),
    .io_a(x856_rdcol_1_io_a),
    .io_b(x856_rdcol_1_io_b),
    .io_flow(x856_rdcol_1_io_flow),
    .io_result(x856_rdcol_1_io_result)
  );
  x814 x858_1 ( // @[Math.scala 366:24:@88415.4]
    .clock(x858_1_clock),
    .reset(x858_1_reset),
    .io_a(x858_1_io_a),
    .io_flow(x858_1_io_flow),
    .io_result(x858_1_io_result)
  );
  x817_div x859_div_1 ( // @[Math.scala 327:24:@88427.4]
    .clock(x859_div_1_clock),
    .reset(x859_div_1_reset),
    .io_a(x859_div_1_io_a),
    .io_flow(x859_div_1_io_flow),
    .io_result(x859_div_1_io_result)
  );
  x758_sum x860_sum_1 ( // @[Math.scala 150:24:@88437.4]
    .clock(x860_sum_1_clock),
    .reset(x860_sum_1_reset),
    .io_a(x860_sum_1_io_a),
    .io_b(x860_sum_1_io_b),
    .io_flow(x860_sum_1_io_flow),
    .io_result(x860_sum_1_io_result)
  );
  RetimeWrapper_714 RetimeWrapper_35 ( // @[package.scala 93:22:@88447.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_725 RetimeWrapper_36 ( // @[package.scala 93:22:@88456.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_724 RetimeWrapper_37 ( // @[package.scala 93:22:@88465.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_712 RetimeWrapper_38 ( // @[package.scala 93:22:@88476.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_39 ( // @[package.scala 93:22:@88497.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_40 ( // @[package.scala 93:22:@88513.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@88531.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_42 ( // @[package.scala 93:22:@88540.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper RetimeWrapper_43 ( // @[package.scala 93:22:@88554.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@88563.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  x758_sum x1240_sum_1 ( // @[Math.scala 150:24:@88610.4]
    .clock(x1240_sum_1_clock),
    .reset(x1240_sum_1_reset),
    .io_a(x1240_sum_1_io_a),
    .io_b(x1240_sum_1_io_b),
    .io_flow(x1240_sum_1_io_flow),
    .io_result(x1240_sum_1_io_result)
  );
  RetimeWrapper_782 RetimeWrapper_45 ( // @[package.scala 93:22:@88620.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_46 ( // @[package.scala 93:22:@88629.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  x758_sum x871_sum_1 ( // @[Math.scala 150:24:@88638.4]
    .clock(x871_sum_1_clock),
    .reset(x871_sum_1_reset),
    .io_a(x871_sum_1_io_a),
    .io_b(x871_sum_1_io_b),
    .io_flow(x871_sum_1_io_flow),
    .io_result(x871_sum_1_io_result)
  );
  RetimeWrapper_785 RetimeWrapper_47 ( // @[package.scala 93:22:@88648.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_48 ( // @[package.scala 93:22:@88657.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_787 RetimeWrapper_49 ( // @[package.scala 93:22:@88666.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_50 ( // @[package.scala 93:22:@88675.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_51 ( // @[package.scala 93:22:@88684.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_52 ( // @[package.scala 93:22:@88696.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_53 ( // @[package.scala 93:22:@88717.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper RetimeWrapper_54 ( // @[package.scala 93:22:@88731.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_55 ( // @[package.scala 93:22:@88746.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x758_sum x877_sum_1 ( // @[Math.scala 150:24:@88755.4]
    .clock(x877_sum_1_clock),
    .reset(x877_sum_1_reset),
    .io_a(x877_sum_1_io_a),
    .io_b(x877_sum_1_io_b),
    .io_flow(x877_sum_1_io_flow),
    .io_result(x877_sum_1_io_result)
  );
  RetimeWrapper_787 RetimeWrapper_56 ( // @[package.scala 93:22:@88765.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_57 ( // @[package.scala 93:22:@88774.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_58 ( // @[package.scala 93:22:@88786.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_59 ( // @[package.scala 93:22:@88807.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper RetimeWrapper_60 ( // @[package.scala 93:22:@88821.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_61 ( // @[package.scala 93:22:@88836.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x758_sum x883_sum_1 ( // @[Math.scala 150:24:@88845.4]
    .clock(x883_sum_1_clock),
    .reset(x883_sum_1_reset),
    .io_a(x883_sum_1_io_a),
    .io_b(x883_sum_1_io_b),
    .io_flow(x883_sum_1_io_flow),
    .io_result(x883_sum_1_io_result)
  );
  RetimeWrapper_787 RetimeWrapper_62 ( // @[package.scala 93:22:@88855.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_63 ( // @[package.scala 93:22:@88864.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_64 ( // @[package.scala 93:22:@88876.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_65 ( // @[package.scala 93:22:@88897.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper RetimeWrapper_66 ( // @[package.scala 93:22:@88911.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_67 ( // @[package.scala 93:22:@88926.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x758_sum x889_sum_1 ( // @[Math.scala 150:24:@88935.4]
    .clock(x889_sum_1_clock),
    .reset(x889_sum_1_reset),
    .io_a(x889_sum_1_io_a),
    .io_b(x889_sum_1_io_b),
    .io_flow(x889_sum_1_io_flow),
    .io_result(x889_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_68 ( // @[package.scala 93:22:@88945.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_787 RetimeWrapper_69 ( // @[package.scala 93:22:@88954.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_70 ( // @[package.scala 93:22:@88966.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_71 ( // @[package.scala 93:22:@88987.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper RetimeWrapper_72 ( // @[package.scala 93:22:@89003.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_73 ( // @[package.scala 93:22:@89018.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x758_sum x895_sum_1 ( // @[Math.scala 150:24:@89027.4]
    .clock(x895_sum_1_clock),
    .reset(x895_sum_1_reset),
    .io_a(x895_sum_1_io_a),
    .io_b(x895_sum_1_io_b),
    .io_flow(x895_sum_1_io_flow),
    .io_result(x895_sum_1_io_result)
  );
  RetimeWrapper_787 RetimeWrapper_74 ( // @[package.scala 93:22:@89037.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_75 ( // @[package.scala 93:22:@89046.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_76 ( // @[package.scala 93:22:@89058.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_77 ( // @[package.scala 93:22:@89079.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper RetimeWrapper_78 ( // @[package.scala 93:22:@89093.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_79 ( // @[package.scala 93:22:@89108.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  x758_sum x901_sum_1 ( // @[Math.scala 150:24:@89117.4]
    .clock(x901_sum_1_clock),
    .reset(x901_sum_1_reset),
    .io_a(x901_sum_1_io_a),
    .io_b(x901_sum_1_io_b),
    .io_flow(x901_sum_1_io_flow),
    .io_result(x901_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_80 ( // @[package.scala 93:22:@89127.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_787 RetimeWrapper_81 ( // @[package.scala 93:22:@89136.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_82 ( // @[package.scala 93:22:@89148.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_83 ( // @[package.scala 93:22:@89169.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper RetimeWrapper_84 ( // @[package.scala 93:22:@89183.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_85 ( // @[package.scala 93:22:@89198.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  x758_sum x907_sum_1 ( // @[Math.scala 150:24:@89207.4]
    .clock(x907_sum_1_clock),
    .reset(x907_sum_1_reset),
    .io_a(x907_sum_1_io_a),
    .io_b(x907_sum_1_io_b),
    .io_flow(x907_sum_1_io_flow),
    .io_result(x907_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_86 ( // @[package.scala 93:22:@89217.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_787 RetimeWrapper_87 ( // @[package.scala 93:22:@89226.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_88 ( // @[package.scala 93:22:@89238.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_89 ( // @[package.scala 93:22:@89259.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper RetimeWrapper_90 ( // @[package.scala 93:22:@89273.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_721 RetimeWrapper_91 ( // @[package.scala 93:22:@89288.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_775 RetimeWrapper_92 ( // @[package.scala 93:22:@89297.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  x758_sum x913_sum_1 ( // @[Math.scala 150:24:@89306.4]
    .clock(x913_sum_1_clock),
    .reset(x913_sum_1_reset),
    .io_a(x913_sum_1_io_a),
    .io_b(x913_sum_1_io_b),
    .io_flow(x913_sum_1_io_flow),
    .io_result(x913_sum_1_io_result)
  );
  RetimeWrapper_838 RetimeWrapper_93 ( // @[package.scala 93:22:@89316.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_94 ( // @[package.scala 93:22:@89325.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_840 RetimeWrapper_95 ( // @[package.scala 93:22:@89334.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_96 ( // @[package.scala 93:22:@89346.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  x758_sum x916_rdcol_1 ( // @[Math.scala 150:24:@89369.4]
    .clock(x916_rdcol_1_clock),
    .reset(x916_rdcol_1_reset),
    .io_a(x916_rdcol_1_io_a),
    .io_b(x916_rdcol_1_io_b),
    .io_flow(x916_rdcol_1_io_flow),
    .io_result(x916_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_97 ( // @[package.scala 93:22:@89384.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  x814 x920_1 ( // @[Math.scala 366:24:@89401.4]
    .clock(x920_1_clock),
    .reset(x920_1_reset),
    .io_a(x920_1_io_a),
    .io_flow(x920_1_io_flow),
    .io_result(x920_1_io_result)
  );
  x817_div x921_div_1 ( // @[Math.scala 327:24:@89413.4]
    .clock(x921_div_1_clock),
    .reset(x921_div_1_reset),
    .io_a(x921_div_1_io_a),
    .io_flow(x921_div_1_io_flow),
    .io_result(x921_div_1_io_result)
  );
  x758_sum x922_sum_1 ( // @[Math.scala 150:24:@89423.4]
    .clock(x922_sum_1_clock),
    .reset(x922_sum_1_reset),
    .io_a(x922_sum_1_io_a),
    .io_b(x922_sum_1_io_b),
    .io_flow(x922_sum_1_io_flow),
    .io_result(x922_sum_1_io_result)
  );
  RetimeWrapper_847 RetimeWrapper_98 ( // @[package.scala 93:22:@89433.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_99 ( // @[package.scala 93:22:@89442.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_100 ( // @[package.scala 93:22:@89454.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  x758_sum x925_rdcol_1 ( // @[Math.scala 150:24:@89479.4]
    .clock(x925_rdcol_1_clock),
    .reset(x925_rdcol_1_reset),
    .io_a(x925_rdcol_1_io_a),
    .io_b(x925_rdcol_1_io_b),
    .io_flow(x925_rdcol_1_io_flow),
    .io_result(x925_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_101 ( // @[package.scala 93:22:@89494.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  x814 x929_1 ( // @[Math.scala 366:24:@89511.4]
    .clock(x929_1_clock),
    .reset(x929_1_reset),
    .io_a(x929_1_io_a),
    .io_flow(x929_1_io_flow),
    .io_result(x929_1_io_result)
  );
  x817_div x930_div_1 ( // @[Math.scala 327:24:@89523.4]
    .clock(x930_div_1_clock),
    .reset(x930_div_1_reset),
    .io_a(x930_div_1_io_a),
    .io_flow(x930_div_1_io_flow),
    .io_result(x930_div_1_io_result)
  );
  x758_sum x931_sum_1 ( // @[Math.scala 150:24:@89533.4]
    .clock(x931_sum_1_clock),
    .reset(x931_sum_1_reset),
    .io_a(x931_sum_1_io_a),
    .io_b(x931_sum_1_io_b),
    .io_flow(x931_sum_1_io_flow),
    .io_result(x931_sum_1_io_result)
  );
  RetimeWrapper_847 RetimeWrapper_102 ( // @[package.scala 93:22:@89543.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_103 ( // @[package.scala 93:22:@89552.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_104 ( // @[package.scala 93:22:@89564.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  x1207_sub x934_rdrow_1 ( // @[Math.scala 191:24:@89587.4]
    .clock(x934_rdrow_1_clock),
    .reset(x934_rdrow_1_reset),
    .io_a(x934_rdrow_1_io_a),
    .io_b(x934_rdrow_1_io_b),
    .io_flow(x934_rdrow_1_io_flow),
    .io_result(x934_rdrow_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_105 ( // @[package.scala 93:22:@89604.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper RetimeWrapper_106 ( // @[package.scala 93:22:@89622.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  x758_sum x1245_sum_1 ( // @[Math.scala 150:24:@89667.4]
    .clock(x1245_sum_1_clock),
    .reset(x1245_sum_1_reset),
    .io_a(x1245_sum_1_io_a),
    .io_b(x1245_sum_1_io_b),
    .io_flow(x1245_sum_1_io_flow),
    .io_result(x1245_sum_1_io_result)
  );
  RetimeWrapper_721 RetimeWrapper_107 ( // @[package.scala 93:22:@89677.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  x758_sum x942_sum_1 ( // @[Math.scala 150:24:@89686.4]
    .clock(x942_sum_1_clock),
    .reset(x942_sum_1_reset),
    .io_a(x942_sum_1_io_a),
    .io_b(x942_sum_1_io_b),
    .io_flow(x942_sum_1_io_flow),
    .io_result(x942_sum_1_io_result)
  );
  RetimeWrapper_708 RetimeWrapper_108 ( // @[package.scala 93:22:@89696.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_109 ( // @[package.scala 93:22:@89705.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_110 ( // @[package.scala 93:22:@89717.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  x758_sum x947_sum_1 ( // @[Math.scala 150:24:@89744.4]
    .clock(x947_sum_1_clock),
    .reset(x947_sum_1_reset),
    .io_a(x947_sum_1_io_a),
    .io_b(x947_sum_1_io_b),
    .io_flow(x947_sum_1_io_flow),
    .io_result(x947_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_111 ( // @[package.scala 93:22:@89754.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_112 ( // @[package.scala 93:22:@89766.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  x758_sum x952_sum_1 ( // @[Math.scala 150:24:@89793.4]
    .clock(x952_sum_1_clock),
    .reset(x952_sum_1_reset),
    .io_a(x952_sum_1_io_a),
    .io_b(x952_sum_1_io_b),
    .io_flow(x952_sum_1_io_flow),
    .io_result(x952_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_113 ( // @[package.scala 93:22:@89803.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_114 ( // @[package.scala 93:22:@89815.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  x758_sum x957_sum_1 ( // @[Math.scala 150:24:@89842.4]
    .clock(x957_sum_1_clock),
    .reset(x957_sum_1_reset),
    .io_a(x957_sum_1_io_a),
    .io_b(x957_sum_1_io_b),
    .io_flow(x957_sum_1_io_flow),
    .io_result(x957_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_115 ( // @[package.scala 93:22:@89852.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_116 ( // @[package.scala 93:22:@89864.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  x758_sum x962_sum_1 ( // @[Math.scala 150:24:@89893.4]
    .clock(x962_sum_1_clock),
    .reset(x962_sum_1_reset),
    .io_a(x962_sum_1_io_a),
    .io_b(x962_sum_1_io_b),
    .io_flow(x962_sum_1_io_flow),
    .io_result(x962_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_117 ( // @[package.scala 93:22:@89903.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_118 ( // @[package.scala 93:22:@89915.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  x758_sum x967_sum_1 ( // @[Math.scala 150:24:@89942.4]
    .clock(x967_sum_1_clock),
    .reset(x967_sum_1_reset),
    .io_a(x967_sum_1_io_a),
    .io_b(x967_sum_1_io_b),
    .io_flow(x967_sum_1_io_flow),
    .io_result(x967_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_119 ( // @[package.scala 93:22:@89952.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_120 ( // @[package.scala 93:22:@89964.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  x758_sum x972_sum_1 ( // @[Math.scala 150:24:@89991.4]
    .clock(x972_sum_1_clock),
    .reset(x972_sum_1_reset),
    .io_a(x972_sum_1_io_a),
    .io_b(x972_sum_1_io_b),
    .io_flow(x972_sum_1_io_flow),
    .io_result(x972_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_121 ( // @[package.scala 93:22:@90001.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_122 ( // @[package.scala 93:22:@90013.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper RetimeWrapper_123 ( // @[package.scala 93:22:@90034.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_709 RetimeWrapper_124 ( // @[package.scala 93:22:@90049.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  x758_sum x977_sum_1 ( // @[Math.scala 150:24:@90058.4]
    .clock(x977_sum_1_clock),
    .reset(x977_sum_1_reset),
    .io_a(x977_sum_1_io_a),
    .io_b(x977_sum_1_io_b),
    .io_flow(x977_sum_1_io_flow),
    .io_result(x977_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_125 ( // @[package.scala 93:22:@90068.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_788 RetimeWrapper_126 ( // @[package.scala 93:22:@90077.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_127 ( // @[package.scala 93:22:@90089.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  x758_sum x982_sum_1 ( // @[Math.scala 150:24:@90116.4]
    .clock(x982_sum_1_clock),
    .reset(x982_sum_1_reset),
    .io_a(x982_sum_1_io_a),
    .io_b(x982_sum_1_io_b),
    .io_flow(x982_sum_1_io_flow),
    .io_result(x982_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_128 ( // @[package.scala 93:22:@90126.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_129 ( // @[package.scala 93:22:@90138.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  x758_sum x987_sum_1 ( // @[Math.scala 150:24:@90165.4]
    .clock(x987_sum_1_clock),
    .reset(x987_sum_1_reset),
    .io_a(x987_sum_1_io_a),
    .io_b(x987_sum_1_io_b),
    .io_flow(x987_sum_1_io_flow),
    .io_result(x987_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_130 ( // @[package.scala 93:22:@90175.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_131 ( // @[package.scala 93:22:@90187.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  x1207_sub x990_rdrow_1 ( // @[Math.scala 191:24:@90210.4]
    .clock(x990_rdrow_1_clock),
    .reset(x990_rdrow_1_reset),
    .io_a(x990_rdrow_1_io_a),
    .io_b(x990_rdrow_1_io_b),
    .io_flow(x990_rdrow_1_io_flow),
    .io_result(x990_rdrow_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_132 ( // @[package.scala 93:22:@90227.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper RetimeWrapper_133 ( // @[package.scala 93:22:@90245.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  x758_sum x1250_sum_1 ( // @[Math.scala 150:24:@90290.4]
    .clock(x1250_sum_1_clock),
    .reset(x1250_sum_1_reset),
    .io_a(x1250_sum_1_io_a),
    .io_b(x1250_sum_1_io_b),
    .io_flow(x1250_sum_1_io_flow),
    .io_result(x1250_sum_1_io_result)
  );
  RetimeWrapper_721 RetimeWrapper_134 ( // @[package.scala 93:22:@90300.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  x758_sum x998_sum_1 ( // @[Math.scala 150:24:@90311.4]
    .clock(x998_sum_1_clock),
    .reset(x998_sum_1_reset),
    .io_a(x998_sum_1_io_a),
    .io_b(x998_sum_1_io_b),
    .io_flow(x998_sum_1_io_flow),
    .io_result(x998_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_135 ( // @[package.scala 93:22:@90321.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_708 RetimeWrapper_136 ( // @[package.scala 93:22:@90330.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_137 ( // @[package.scala 93:22:@90342.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  x758_sum x1003_sum_1 ( // @[Math.scala 150:24:@90369.4]
    .clock(x1003_sum_1_clock),
    .reset(x1003_sum_1_reset),
    .io_a(x1003_sum_1_io_a),
    .io_b(x1003_sum_1_io_b),
    .io_flow(x1003_sum_1_io_flow),
    .io_result(x1003_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_138 ( // @[package.scala 93:22:@90379.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_139 ( // @[package.scala 93:22:@90391.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  x758_sum x1008_sum_1 ( // @[Math.scala 150:24:@90418.4]
    .clock(x1008_sum_1_clock),
    .reset(x1008_sum_1_reset),
    .io_a(x1008_sum_1_io_a),
    .io_b(x1008_sum_1_io_b),
    .io_flow(x1008_sum_1_io_flow),
    .io_result(x1008_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_140 ( // @[package.scala 93:22:@90428.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_141 ( // @[package.scala 93:22:@90440.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  x758_sum x1013_sum_1 ( // @[Math.scala 150:24:@90467.4]
    .clock(x1013_sum_1_clock),
    .reset(x1013_sum_1_reset),
    .io_a(x1013_sum_1_io_a),
    .io_b(x1013_sum_1_io_b),
    .io_flow(x1013_sum_1_io_flow),
    .io_result(x1013_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_142 ( // @[package.scala 93:22:@90477.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_143 ( // @[package.scala 93:22:@90489.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  x758_sum x1018_sum_1 ( // @[Math.scala 150:24:@90516.4]
    .clock(x1018_sum_1_clock),
    .reset(x1018_sum_1_reset),
    .io_a(x1018_sum_1_io_a),
    .io_b(x1018_sum_1_io_b),
    .io_flow(x1018_sum_1_io_flow),
    .io_result(x1018_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_144 ( // @[package.scala 93:22:@90526.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_145 ( // @[package.scala 93:22:@90538.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  x758_sum x1023_sum_1 ( // @[Math.scala 150:24:@90565.4]
    .clock(x1023_sum_1_clock),
    .reset(x1023_sum_1_reset),
    .io_a(x1023_sum_1_io_a),
    .io_b(x1023_sum_1_io_b),
    .io_flow(x1023_sum_1_io_flow),
    .io_result(x1023_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_146 ( // @[package.scala 93:22:@90575.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_147 ( // @[package.scala 93:22:@90587.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  x758_sum x1028_sum_1 ( // @[Math.scala 150:24:@90614.4]
    .clock(x1028_sum_1_clock),
    .reset(x1028_sum_1_reset),
    .io_a(x1028_sum_1_io_a),
    .io_b(x1028_sum_1_io_b),
    .io_flow(x1028_sum_1_io_flow),
    .io_result(x1028_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_148 ( // @[package.scala 93:22:@90624.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_149 ( // @[package.scala 93:22:@90636.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_709 RetimeWrapper_150 ( // @[package.scala 93:22:@90663.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  x758_sum x1033_sum_1 ( // @[Math.scala 150:24:@90672.4]
    .clock(x1033_sum_1_clock),
    .reset(x1033_sum_1_reset),
    .io_a(x1033_sum_1_io_a),
    .io_b(x1033_sum_1_io_b),
    .io_flow(x1033_sum_1_io_flow),
    .io_result(x1033_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_151 ( // @[package.scala 93:22:@90682.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_152 ( // @[package.scala 93:22:@90691.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_153 ( // @[package.scala 93:22:@90703.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  x758_sum x1038_sum_1 ( // @[Math.scala 150:24:@90732.4]
    .clock(x1038_sum_1_clock),
    .reset(x1038_sum_1_reset),
    .io_a(x1038_sum_1_io_a),
    .io_b(x1038_sum_1_io_b),
    .io_flow(x1038_sum_1_io_flow),
    .io_result(x1038_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_154 ( // @[package.scala 93:22:@90742.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_155 ( // @[package.scala 93:22:@90754.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  x758_sum x1043_sum_1 ( // @[Math.scala 150:24:@90781.4]
    .clock(x1043_sum_1_clock),
    .reset(x1043_sum_1_reset),
    .io_a(x1043_sum_1_io_a),
    .io_b(x1043_sum_1_io_b),
    .io_flow(x1043_sum_1_io_flow),
    .io_result(x1043_sum_1_io_result)
  );
  RetimeWrapper_788 RetimeWrapper_156 ( // @[package.scala 93:22:@90791.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_786 RetimeWrapper_157 ( // @[package.scala 93:22:@90803.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_158 ( // @[package.scala 93:22:@90826.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_159 ( // @[package.scala 93:22:@90838.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_160 ( // @[package.scala 93:22:@90850.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_161 ( // @[package.scala 93:22:@90862.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_162 ( // @[package.scala 93:22:@90874.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_65 RetimeWrapper_163 ( // @[package.scala 93:22:@90884.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  x1051_x15 x1051_x15_1 ( // @[Math.scala 150:24:@90893.4]
    .io_a(x1051_x15_1_io_a),
    .io_b(x1051_x15_1_io_b),
    .io_result(x1051_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_164 ( // @[package.scala 93:22:@90903.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  x1051_x15 x1052_x16_1 ( // @[Math.scala 150:24:@90912.4]
    .io_a(x1052_x16_1_io_a),
    .io_b(x1052_x16_1_io_b),
    .io_result(x1052_x16_1_io_result)
  );
  x1051_x15 x1053_x15_1 ( // @[Math.scala 150:24:@90922.4]
    .io_a(x1053_x15_1_io_a),
    .io_b(x1053_x15_1_io_b),
    .io_result(x1053_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_165 ( // @[package.scala 93:22:@90932.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  x1051_x15 x1054_x16_1 ( // @[Math.scala 150:24:@90941.4]
    .io_a(x1054_x16_1_io_a),
    .io_b(x1054_x16_1_io_b),
    .io_result(x1054_x16_1_io_result)
  );
  x1051_x15 x1055_x15_1 ( // @[Math.scala 150:24:@90951.4]
    .io_a(x1055_x15_1_io_a),
    .io_b(x1055_x15_1_io_b),
    .io_result(x1055_x15_1_io_result)
  );
  x1051_x15 x1056_x16_1 ( // @[Math.scala 150:24:@90961.4]
    .io_a(x1056_x16_1_io_a),
    .io_b(x1056_x16_1_io_b),
    .io_result(x1056_x16_1_io_result)
  );
  x1051_x15 x1057_x15_1 ( // @[Math.scala 150:24:@90971.4]
    .io_a(x1057_x15_1_io_a),
    .io_b(x1057_x15_1_io_b),
    .io_result(x1057_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_166 ( // @[package.scala 93:22:@90981.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  x1058_sum x1058_sum_1 ( // @[Math.scala 150:24:@90990.4]
    .clock(x1058_sum_1_clock),
    .reset(x1058_sum_1_reset),
    .io_a(x1058_sum_1_io_a),
    .io_b(x1058_sum_1_io_b),
    .io_flow(x1058_sum_1_io_flow),
    .io_result(x1058_sum_1_io_result)
  );
  RetimeWrapper_935 RetimeWrapper_167 ( // @[package.scala 93:22:@91009.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_168 ( // @[package.scala 93:22:@91021.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_169 ( // @[package.scala 93:22:@91033.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_170 ( // @[package.scala 93:22:@91045.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_171 ( // @[package.scala 93:22:@91057.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_65 RetimeWrapper_172 ( // @[package.scala 93:22:@91067.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  x1051_x15 x1065_x15_1 ( // @[Math.scala 150:24:@91076.4]
    .io_a(x1065_x15_1_io_a),
    .io_b(x1065_x15_1_io_b),
    .io_result(x1065_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_173 ( // @[package.scala 93:22:@91086.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  x1051_x15 x1066_x16_1 ( // @[Math.scala 150:24:@91095.4]
    .io_a(x1066_x16_1_io_a),
    .io_b(x1066_x16_1_io_b),
    .io_result(x1066_x16_1_io_result)
  );
  x1051_x15 x1067_x15_1 ( // @[Math.scala 150:24:@91105.4]
    .io_a(x1067_x15_1_io_a),
    .io_b(x1067_x15_1_io_b),
    .io_result(x1067_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_174 ( // @[package.scala 93:22:@91115.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  x1051_x15 x1068_x16_1 ( // @[Math.scala 150:24:@91124.4]
    .io_a(x1068_x16_1_io_a),
    .io_b(x1068_x16_1_io_b),
    .io_result(x1068_x16_1_io_result)
  );
  x1051_x15 x1069_x15_1 ( // @[Math.scala 150:24:@91134.4]
    .io_a(x1069_x15_1_io_a),
    .io_b(x1069_x15_1_io_b),
    .io_result(x1069_x15_1_io_result)
  );
  x1051_x15 x1070_x16_1 ( // @[Math.scala 150:24:@91144.4]
    .io_a(x1070_x16_1_io_a),
    .io_b(x1070_x16_1_io_b),
    .io_result(x1070_x16_1_io_result)
  );
  x1051_x15 x1071_x15_1 ( // @[Math.scala 150:24:@91154.4]
    .io_a(x1071_x15_1_io_a),
    .io_b(x1071_x15_1_io_b),
    .io_result(x1071_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_175 ( // @[package.scala 93:22:@91164.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  x1058_sum x1072_sum_1 ( // @[Math.scala 150:24:@91173.4]
    .clock(x1072_sum_1_clock),
    .reset(x1072_sum_1_reset),
    .io_a(x1072_sum_1_io_a),
    .io_b(x1072_sum_1_io_b),
    .io_flow(x1072_sum_1_io_flow),
    .io_result(x1072_sum_1_io_result)
  );
  RetimeWrapper_935 RetimeWrapper_176 ( // @[package.scala 93:22:@91192.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_177 ( // @[package.scala 93:22:@91206.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_178 ( // @[package.scala 93:22:@91218.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_179 ( // @[package.scala 93:22:@91230.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  x1051_x15 x1078_x15_1 ( // @[Math.scala 150:24:@91240.4]
    .io_a(x1078_x15_1_io_a),
    .io_b(x1078_x15_1_io_b),
    .io_result(x1078_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_180 ( // @[package.scala 93:22:@91250.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  x1051_x15 x1079_x16_1 ( // @[Math.scala 150:24:@91259.4]
    .io_a(x1079_x16_1_io_a),
    .io_b(x1079_x16_1_io_b),
    .io_result(x1079_x16_1_io_result)
  );
  x1051_x15 x1080_x15_1 ( // @[Math.scala 150:24:@91269.4]
    .io_a(x1080_x15_1_io_a),
    .io_b(x1080_x15_1_io_b),
    .io_result(x1080_x15_1_io_result)
  );
  x1051_x15 x1081_x16_1 ( // @[Math.scala 150:24:@91279.4]
    .io_a(x1081_x16_1_io_a),
    .io_b(x1081_x16_1_io_b),
    .io_result(x1081_x16_1_io_result)
  );
  x1051_x15 x1082_x15_1 ( // @[Math.scala 150:24:@91289.4]
    .io_a(x1082_x15_1_io_a),
    .io_b(x1082_x15_1_io_b),
    .io_result(x1082_x15_1_io_result)
  );
  x1051_x15 x1083_x16_1 ( // @[Math.scala 150:24:@91299.4]
    .io_a(x1083_x16_1_io_a),
    .io_b(x1083_x16_1_io_b),
    .io_result(x1083_x16_1_io_result)
  );
  x1051_x15 x1084_x15_1 ( // @[Math.scala 150:24:@91309.4]
    .io_a(x1084_x15_1_io_a),
    .io_b(x1084_x15_1_io_b),
    .io_result(x1084_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_181 ( // @[package.scala 93:22:@91319.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  x1058_sum x1085_sum_1 ( // @[Math.scala 150:24:@91328.4]
    .clock(x1085_sum_1_clock),
    .reset(x1085_sum_1_reset),
    .io_a(x1085_sum_1_io_a),
    .io_b(x1085_sum_1_io_b),
    .io_flow(x1085_sum_1_io_flow),
    .io_result(x1085_sum_1_io_result)
  );
  RetimeWrapper_935 RetimeWrapper_182 ( // @[package.scala 93:22:@91347.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_183 ( // @[package.scala 93:22:@91359.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_184 ( // @[package.scala 93:22:@91371.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_185 ( // @[package.scala 93:22:@91383.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  x1051_x15 x1091_x15_1 ( // @[Math.scala 150:24:@91393.4]
    .io_a(x1091_x15_1_io_a),
    .io_b(x1091_x15_1_io_b),
    .io_result(x1091_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_186 ( // @[package.scala 93:22:@91403.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  x1051_x15 x1092_x16_1 ( // @[Math.scala 150:24:@91412.4]
    .io_a(x1092_x16_1_io_a),
    .io_b(x1092_x16_1_io_b),
    .io_result(x1092_x16_1_io_result)
  );
  x1051_x15 x1093_x15_1 ( // @[Math.scala 150:24:@91422.4]
    .io_a(x1093_x15_1_io_a),
    .io_b(x1093_x15_1_io_b),
    .io_result(x1093_x15_1_io_result)
  );
  x1051_x15 x1094_x16_1 ( // @[Math.scala 150:24:@91432.4]
    .io_a(x1094_x16_1_io_a),
    .io_b(x1094_x16_1_io_b),
    .io_result(x1094_x16_1_io_result)
  );
  x1051_x15 x1095_x15_1 ( // @[Math.scala 150:24:@91442.4]
    .io_a(x1095_x15_1_io_a),
    .io_b(x1095_x15_1_io_b),
    .io_result(x1095_x15_1_io_result)
  );
  x1051_x15 x1096_x16_1 ( // @[Math.scala 150:24:@91452.4]
    .io_a(x1096_x16_1_io_a),
    .io_b(x1096_x16_1_io_b),
    .io_result(x1096_x16_1_io_result)
  );
  x1051_x15 x1097_x15_1 ( // @[Math.scala 150:24:@91462.4]
    .io_a(x1097_x15_1_io_a),
    .io_b(x1097_x15_1_io_b),
    .io_result(x1097_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_187 ( // @[package.scala 93:22:@91472.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  x1058_sum x1098_sum_1 ( // @[Math.scala 150:24:@91481.4]
    .clock(x1098_sum_1_clock),
    .reset(x1098_sum_1_reset),
    .io_a(x1098_sum_1_io_a),
    .io_b(x1098_sum_1_io_b),
    .io_flow(x1098_sum_1_io_flow),
    .io_result(x1098_sum_1_io_result)
  );
  RetimeWrapper_935 RetimeWrapper_188 ( // @[package.scala 93:22:@91500.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_189 ( // @[package.scala 93:22:@91512.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_190 ( // @[package.scala 93:22:@91524.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_191 ( // @[package.scala 93:22:@91536.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  x1051_x15 x1104_x15_1 ( // @[Math.scala 150:24:@91546.4]
    .io_a(x1104_x15_1_io_a),
    .io_b(x1104_x15_1_io_b),
    .io_result(x1104_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_192 ( // @[package.scala 93:22:@91556.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  x1051_x15 x1105_x16_1 ( // @[Math.scala 150:24:@91565.4]
    .io_a(x1105_x16_1_io_a),
    .io_b(x1105_x16_1_io_b),
    .io_result(x1105_x16_1_io_result)
  );
  x1051_x15 x1106_x15_1 ( // @[Math.scala 150:24:@91575.4]
    .io_a(x1106_x15_1_io_a),
    .io_b(x1106_x15_1_io_b),
    .io_result(x1106_x15_1_io_result)
  );
  x1051_x15 x1107_x16_1 ( // @[Math.scala 150:24:@91585.4]
    .io_a(x1107_x16_1_io_a),
    .io_b(x1107_x16_1_io_b),
    .io_result(x1107_x16_1_io_result)
  );
  x1051_x15 x1108_x15_1 ( // @[Math.scala 150:24:@91595.4]
    .io_a(x1108_x15_1_io_a),
    .io_b(x1108_x15_1_io_b),
    .io_result(x1108_x15_1_io_result)
  );
  x1051_x15 x1109_x16_1 ( // @[Math.scala 150:24:@91605.4]
    .io_a(x1109_x16_1_io_a),
    .io_b(x1109_x16_1_io_b),
    .io_result(x1109_x16_1_io_result)
  );
  x1051_x15 x1110_x15_1 ( // @[Math.scala 150:24:@91615.4]
    .io_a(x1110_x15_1_io_a),
    .io_b(x1110_x15_1_io_b),
    .io_result(x1110_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_193 ( // @[package.scala 93:22:@91625.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  x1058_sum x1111_sum_1 ( // @[Math.scala 150:24:@91634.4]
    .clock(x1111_sum_1_clock),
    .reset(x1111_sum_1_reset),
    .io_a(x1111_sum_1_io_a),
    .io_b(x1111_sum_1_io_b),
    .io_flow(x1111_sum_1_io_flow),
    .io_result(x1111_sum_1_io_result)
  );
  RetimeWrapper_935 RetimeWrapper_194 ( // @[package.scala 93:22:@91653.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_195 ( // @[package.scala 93:22:@91665.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_196 ( // @[package.scala 93:22:@91677.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_197 ( // @[package.scala 93:22:@91689.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  x1051_x15 x1117_x15_1 ( // @[Math.scala 150:24:@91699.4]
    .io_a(x1117_x15_1_io_a),
    .io_b(x1117_x15_1_io_b),
    .io_result(x1117_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_198 ( // @[package.scala 93:22:@91709.4]
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  x1051_x15 x1118_x16_1 ( // @[Math.scala 150:24:@91720.4]
    .io_a(x1118_x16_1_io_a),
    .io_b(x1118_x16_1_io_b),
    .io_result(x1118_x16_1_io_result)
  );
  x1051_x15 x1119_x15_1 ( // @[Math.scala 150:24:@91730.4]
    .io_a(x1119_x15_1_io_a),
    .io_b(x1119_x15_1_io_b),
    .io_result(x1119_x15_1_io_result)
  );
  x1051_x15 x1120_x16_1 ( // @[Math.scala 150:24:@91740.4]
    .io_a(x1120_x16_1_io_a),
    .io_b(x1120_x16_1_io_b),
    .io_result(x1120_x16_1_io_result)
  );
  x1051_x15 x1121_x15_1 ( // @[Math.scala 150:24:@91750.4]
    .io_a(x1121_x15_1_io_a),
    .io_b(x1121_x15_1_io_b),
    .io_result(x1121_x15_1_io_result)
  );
  x1051_x15 x1122_x16_1 ( // @[Math.scala 150:24:@91760.4]
    .io_a(x1122_x16_1_io_a),
    .io_b(x1122_x16_1_io_b),
    .io_result(x1122_x16_1_io_result)
  );
  x1051_x15 x1123_x15_1 ( // @[Math.scala 150:24:@91770.4]
    .io_a(x1123_x15_1_io_a),
    .io_b(x1123_x15_1_io_b),
    .io_result(x1123_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_199 ( // @[package.scala 93:22:@91780.4]
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  x1058_sum x1124_sum_1 ( // @[Math.scala 150:24:@91789.4]
    .clock(x1124_sum_1_clock),
    .reset(x1124_sum_1_reset),
    .io_a(x1124_sum_1_io_a),
    .io_b(x1124_sum_1_io_b),
    .io_flow(x1124_sum_1_io_flow),
    .io_result(x1124_sum_1_io_result)
  );
  RetimeWrapper_935 RetimeWrapper_200 ( // @[package.scala 93:22:@91808.4]
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_201 ( // @[package.scala 93:22:@91820.4]
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_202 ( // @[package.scala 93:22:@91832.4]
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_203 ( // @[package.scala 93:22:@91844.4]
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  x1051_x15 x1130_x15_1 ( // @[Math.scala 150:24:@91854.4]
    .io_a(x1130_x15_1_io_a),
    .io_b(x1130_x15_1_io_b),
    .io_result(x1130_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_204 ( // @[package.scala 93:22:@91864.4]
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  x1051_x15 x1131_x16_1 ( // @[Math.scala 150:24:@91873.4]
    .io_a(x1131_x16_1_io_a),
    .io_b(x1131_x16_1_io_b),
    .io_result(x1131_x16_1_io_result)
  );
  x1051_x15 x1132_x15_1 ( // @[Math.scala 150:24:@91883.4]
    .io_a(x1132_x15_1_io_a),
    .io_b(x1132_x15_1_io_b),
    .io_result(x1132_x15_1_io_result)
  );
  x1051_x15 x1133_x16_1 ( // @[Math.scala 150:24:@91893.4]
    .io_a(x1133_x16_1_io_a),
    .io_b(x1133_x16_1_io_b),
    .io_result(x1133_x16_1_io_result)
  );
  x1051_x15 x1134_x15_1 ( // @[Math.scala 150:24:@91903.4]
    .io_a(x1134_x15_1_io_a),
    .io_b(x1134_x15_1_io_b),
    .io_result(x1134_x15_1_io_result)
  );
  x1051_x15 x1135_x16_1 ( // @[Math.scala 150:24:@91913.4]
    .io_a(x1135_x16_1_io_a),
    .io_b(x1135_x16_1_io_b),
    .io_result(x1135_x16_1_io_result)
  );
  x1051_x15 x1136_x15_1 ( // @[Math.scala 150:24:@91923.4]
    .io_a(x1136_x15_1_io_a),
    .io_b(x1136_x15_1_io_b),
    .io_result(x1136_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_205 ( // @[package.scala 93:22:@91933.4]
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  x1058_sum x1137_sum_1 ( // @[Math.scala 150:24:@91942.4]
    .clock(x1137_sum_1_clock),
    .reset(x1137_sum_1_reset),
    .io_a(x1137_sum_1_io_a),
    .io_b(x1137_sum_1_io_b),
    .io_flow(x1137_sum_1_io_flow),
    .io_result(x1137_sum_1_io_result)
  );
  RetimeWrapper_935 RetimeWrapper_206 ( // @[package.scala 93:22:@91961.4]
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper_937 RetimeWrapper_207 ( // @[package.scala 93:22:@91973.4]
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_208 ( // @[package.scala 93:22:@91985.4]
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper_935 RetimeWrapper_209 ( // @[package.scala 93:22:@91997.4]
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  x1051_x15 x1143_x15_1 ( // @[Math.scala 150:24:@92007.4]
    .io_a(x1143_x15_1_io_a),
    .io_b(x1143_x15_1_io_b),
    .io_result(x1143_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_210 ( // @[package.scala 93:22:@92017.4]
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  x1051_x15 x1144_x16_1 ( // @[Math.scala 150:24:@92026.4]
    .io_a(x1144_x16_1_io_a),
    .io_b(x1144_x16_1_io_b),
    .io_result(x1144_x16_1_io_result)
  );
  x1051_x15 x1145_x15_1 ( // @[Math.scala 150:24:@92036.4]
    .io_a(x1145_x15_1_io_a),
    .io_b(x1145_x15_1_io_b),
    .io_result(x1145_x15_1_io_result)
  );
  x1051_x15 x1146_x16_1 ( // @[Math.scala 150:24:@92046.4]
    .io_a(x1146_x16_1_io_a),
    .io_b(x1146_x16_1_io_b),
    .io_result(x1146_x16_1_io_result)
  );
  x1051_x15 x1147_x15_1 ( // @[Math.scala 150:24:@92056.4]
    .io_a(x1147_x15_1_io_a),
    .io_b(x1147_x15_1_io_b),
    .io_result(x1147_x15_1_io_result)
  );
  x1051_x15 x1148_x16_1 ( // @[Math.scala 150:24:@92066.4]
    .io_a(x1148_x16_1_io_a),
    .io_b(x1148_x16_1_io_b),
    .io_result(x1148_x16_1_io_result)
  );
  x1051_x15 x1149_x15_1 ( // @[Math.scala 150:24:@92076.4]
    .io_a(x1149_x15_1_io_a),
    .io_b(x1149_x15_1_io_b),
    .io_result(x1149_x15_1_io_result)
  );
  RetimeWrapper_65 RetimeWrapper_211 ( // @[package.scala 93:22:@92086.4]
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  x1058_sum x1150_sum_1 ( // @[Math.scala 150:24:@92095.4]
    .clock(x1150_sum_1_clock),
    .reset(x1150_sum_1_reset),
    .io_a(x1150_sum_1_io_a),
    .io_b(x1150_sum_1_io_b),
    .io_flow(x1150_sum_1_io_flow),
    .io_result(x1150_sum_1_io_result)
  );
  RetimeWrapper_997 RetimeWrapper_212 ( // @[package.scala 93:22:@92130.4]
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  RetimeWrapper_56 RetimeWrapper_213 ( // @[package.scala 93:22:@92139.4]
    .clock(RetimeWrapper_213_clock),
    .reset(RetimeWrapper_213_reset),
    .io_flow(RetimeWrapper_213_io_flow),
    .io_in(RetimeWrapper_213_io_in),
    .io_out(RetimeWrapper_213_io_out)
  );
  RetimeWrapper_56 RetimeWrapper_214 ( // @[package.scala 93:22:@92148.4]
    .clock(RetimeWrapper_214_clock),
    .reset(RetimeWrapper_214_reset),
    .io_flow(RetimeWrapper_214_io_flow),
    .io_in(RetimeWrapper_214_io_in),
    .io_out(RetimeWrapper_214_io_out)
  );
  RetimeWrapper_56 RetimeWrapper_215 ( // @[package.scala 93:22:@92157.4]
    .clock(RetimeWrapper_215_clock),
    .reset(RetimeWrapper_215_reset),
    .io_flow(RetimeWrapper_215_io_flow),
    .io_in(RetimeWrapper_215_io_in),
    .io_out(RetimeWrapper_215_io_out)
  );
  assign b801 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 62:18:@87288.4]
  assign b802 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 63:18:@87289.4]
  assign _T_205 = b801 & b802; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 67:30:@87291.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 67:37:@87292.4]
  assign _T_210 = io_in_x744_TID == 8'h0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 69:76:@87297.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 69:62:@87298.4]
  assign _T_213 = io_in_x744_TDEST == 8'h0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 69:101:@87299.4]
  assign x1256_x803_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@87308.4 package.scala 96:25:@87309.4]
  assign b799_number = __io_result; // @[Math.scala 712:22:@87273.4 Math.scala 713:14:@87274.4]
  assign _T_254 = $signed(b799_number); // @[Math.scala 499:52:@87585.4]
  assign x808 = $signed(32'sh1) == $signed(_T_254); // @[Math.scala 499:44:@87593.4]
  assign x809 = $signed(32'sh2) == $signed(_T_254); // @[Math.scala 499:44:@87600.4]
  assign x810 = $signed(32'sh3) == $signed(_T_254); // @[Math.scala 499:44:@87607.4]
  assign _T_301 = x808 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@87619.4]
  assign _T_303 = x809 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@87620.4]
  assign _T_305 = x810 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@87621.4]
  assign _T_307 = _T_301 | _T_303; // @[Mux.scala 19:72:@87623.4]
  assign x1257_x811_D2_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@87636.4 package.scala 96:25:@87637.4]
  assign _T_322 = $signed(x1257_x811_D2_number); // @[Math.scala 406:49:@87643.4]
  assign _T_324 = $signed(_T_322) & $signed(32'sh3); // @[Math.scala 406:56:@87645.4]
  assign _T_325 = $signed(_T_324); // @[Math.scala 406:56:@87646.4]
  assign _T_337 = x1257_x811_D2_number[31]; // @[FixedPoint.scala 50:25:@87664.4]
  assign _T_341 = _T_337 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@87666.4]
  assign _T_342 = x1257_x811_D2_number[31:2]; // @[FixedPoint.scala 18:52:@87667.4]
  assign x815_number = {_T_341,_T_342}; // @[Cat.scala 30:58:@87668.4]
  assign _GEN_0 = {{7'd0}, x815_number}; // @[Math.scala 450:32:@87673.4]
  assign _T_347 = _GEN_0 << 7; // @[Math.scala 450:32:@87673.4]
  assign _GEN_1 = {{6'd0}, x815_number}; // @[Math.scala 450:32:@87678.4]
  assign _T_351 = _GEN_1 << 6; // @[Math.scala 450:32:@87678.4]
  assign _T_387 = ~ io_sigsIn_break; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:101:@87776.4]
  assign _T_391 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@87784.4 package.scala 96:25:@87785.4]
  assign _T_393 = io_rr ? _T_391 : 1'h0; // @[implicits.scala 55:10:@87786.4]
  assign _T_394 = _T_387 & _T_393; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:118:@87787.4]
  assign _T_396 = _T_394 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:207:@87789.4]
  assign _T_397 = _T_396 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:226:@87790.4]
  assign x1264_b801_D28 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@87773.4 package.scala 96:25:@87774.4]
  assign _T_398 = _T_397 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 127:252:@87791.4]
  assign x1260_b802_D28 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@87737.4 package.scala 96:25:@87738.4]
  assign _T_442 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@87891.4 package.scala 96:25:@87892.4]
  assign _T_444 = io_rr ? _T_442 : 1'h0; // @[implicits.scala 55:10:@87893.4]
  assign _T_445 = _T_387 & _T_444; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:118:@87894.4]
  assign _T_447 = _T_445 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:207:@87896.4]
  assign _T_448 = _T_447 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:226:@87897.4]
  assign _T_449 = _T_448 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 150:252:@87898.4]
  assign _T_490 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@87989.4 package.scala 96:25:@87990.4]
  assign _T_492 = io_rr ? _T_490 : 1'h0; // @[implicits.scala 55:10:@87991.4]
  assign _T_493 = _T_387 & _T_492; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:118:@87992.4]
  assign _T_495 = _T_493 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:207:@87994.4]
  assign _T_496 = _T_495 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:226:@87995.4]
  assign _T_497 = _T_496 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 171:252:@87996.4]
  assign _T_540 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@88089.4 package.scala 96:25:@88090.4]
  assign _T_542 = io_rr ? _T_540 : 1'h0; // @[implicits.scala 55:10:@88091.4]
  assign _T_543 = _T_387 & _T_542; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:166:@88092.4]
  assign _T_545 = _T_543 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:255:@88094.4]
  assign _T_546 = _T_545 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:274:@88095.4]
  assign _T_547 = _T_546 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 200:300:@88096.4]
  assign _T_588 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@88187.4 package.scala 96:25:@88188.4]
  assign _T_590 = io_rr ? _T_588 : 1'h0; // @[implicits.scala 55:10:@88189.4]
  assign _T_591 = _T_387 & _T_590; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:166:@88190.4]
  assign _T_593 = _T_591 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:255:@88192.4]
  assign _T_594 = _T_593 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:274:@88193.4]
  assign _T_595 = _T_594 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 221:300:@88194.4]
  assign _T_636 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@88285.4 package.scala 96:25:@88286.4]
  assign _T_638 = io_rr ? _T_636 : 1'h0; // @[implicits.scala 55:10:@88287.4]
  assign _T_639 = _T_387 & _T_638; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:166:@88288.4]
  assign _T_641 = _T_639 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:255:@88290.4]
  assign _T_642 = _T_641 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:274:@88291.4]
  assign _T_643 = _T_642 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 242:300:@88292.4]
  assign _T_684 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@88383.4 package.scala 96:25:@88384.4]
  assign _T_686 = io_rr ? _T_684 : 1'h0; // @[implicits.scala 55:10:@88385.4]
  assign _T_687 = _T_387 & _T_686; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:166:@88386.4]
  assign _T_689 = _T_687 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:255:@88388.4]
  assign _T_690 = _T_689 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:274:@88389.4]
  assign _T_691 = _T_690 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 263:300:@88390.4]
  assign _T_732 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@88481.4 package.scala 96:25:@88482.4]
  assign _T_734 = io_rr ? _T_732 : 1'h0; // @[implicits.scala 55:10:@88483.4]
  assign _T_735 = _T_387 & _T_734; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:166:@88484.4]
  assign _T_737 = _T_735 & _T_387; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:255:@88486.4]
  assign _T_738 = _T_737 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:274:@88487.4]
  assign _T_739 = _T_738 & x1264_b801_D28; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 284:300:@88488.4]
  assign x1287_b799_D30_number = RetimeWrapper_39_io_out; // @[package.scala 96:25:@88502.4 package.scala 96:25:@88503.4]
  assign _T_751 = $signed(x1287_b799_D30_number); // @[Math.scala 406:49:@88509.4]
  assign _T_753 = $signed(_T_751) & $signed(32'sh3); // @[Math.scala 406:56:@88511.4]
  assign _T_754 = $signed(_T_753); // @[Math.scala 406:56:@88512.4]
  assign _T_758 = $signed(RetimeWrapper_40_io_out); // @[package.scala 96:25:@88520.4]
  assign x1236_number = $unsigned(_T_758); // @[implicits.scala 133:21:@88522.4]
  assign x1288_x856_rdcol_D30_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@88545.4 package.scala 96:25:@88546.4]
  assign _T_778 = $signed(x1288_x856_rdcol_D30_number); // @[Math.scala 465:37:@88551.4]
  assign x1289_x864_D1 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@88568.4 package.scala 96:25:@88569.4]
  assign x865 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@88559.4 package.scala 96:25:@88560.4]
  assign x866 = x1289_x864_D1 | x865; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 305:25:@88572.4]
  assign _T_799 = $signed(x1236_number); // @[Math.scala 406:49:@88583.4]
  assign _T_801 = $signed(_T_799) & $signed(32'sh3); // @[Math.scala 406:56:@88585.4]
  assign _T_802 = $signed(_T_801); // @[Math.scala 406:56:@88586.4]
  assign _T_807 = x1236_number[31]; // @[FixedPoint.scala 50:25:@88592.4]
  assign _T_811 = _T_807 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@88594.4]
  assign _T_812 = x1236_number[31:2]; // @[FixedPoint.scala 18:52:@88595.4]
  assign x869_number = {_T_811,_T_812}; // @[Cat.scala 30:58:@88596.4]
  assign _GEN_2 = {{7'd0}, x869_number}; // @[Math.scala 450:32:@88601.4]
  assign _T_817 = _GEN_2 << 7; // @[Math.scala 450:32:@88601.4]
  assign _GEN_3 = {{6'd0}, x869_number}; // @[Math.scala 450:32:@88606.4]
  assign _T_821 = _GEN_3 << 6; // @[Math.scala 450:32:@88606.4]
  assign _T_860 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@88701.4 package.scala 96:25:@88702.4]
  assign _T_862 = io_rr ? _T_860 : 1'h0; // @[implicits.scala 55:10:@88703.4]
  assign _T_863 = _T_387 & _T_862; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 340:194:@88704.4]
  assign x1295_x867_D20 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@88680.4 package.scala 96:25:@88681.4]
  assign _T_864 = _T_863 & x1295_x867_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 340:283:@88705.4]
  assign x1296_b801_D52 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@88689.4 package.scala 96:25:@88690.4]
  assign _T_865 = _T_864 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 340:292:@88706.4]
  assign x1293_b802_D52 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@88662.4 package.scala 96:25:@88663.4]
  assign x1297_x850_rdcol_D30_number = RetimeWrapper_53_io_out; // @[package.scala 96:25:@88722.4 package.scala 96:25:@88723.4]
  assign _T_876 = $signed(x1297_x850_rdcol_D30_number); // @[Math.scala 465:37:@88728.4]
  assign x874 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@88736.4 package.scala 96:25:@88737.4]
  assign x875 = x1289_x864_D1 | x874; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 348:25:@88740.4]
  assign _T_908 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@88791.4 package.scala 96:25:@88792.4]
  assign _T_910 = io_rr ? _T_908 : 1'h0; // @[implicits.scala 55:10:@88793.4]
  assign _T_911 = _T_387 & _T_910; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:194:@88794.4]
  assign x1300_x876_D20 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@88779.4 package.scala 96:25:@88780.4]
  assign _T_912 = _T_911 & x1300_x876_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:283:@88795.4]
  assign _T_913 = _T_912 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:292:@88796.4]
  assign x1301_x844_rdcol_D30_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@88812.4 package.scala 96:25:@88813.4]
  assign _T_924 = $signed(x1301_x844_rdcol_D30_number); // @[Math.scala 465:37:@88818.4]
  assign x880 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@88826.4 package.scala 96:25:@88827.4]
  assign x881 = x1289_x864_D1 | x880; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 371:25:@88830.4]
  assign _T_956 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@88881.4 package.scala 96:25:@88882.4]
  assign _T_958 = io_rr ? _T_956 : 1'h0; // @[implicits.scala 55:10:@88883.4]
  assign _T_959 = _T_387 & _T_958; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:194:@88884.4]
  assign x1304_x882_D20 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@88869.4 package.scala 96:25:@88870.4]
  assign _T_960 = _T_959 & x1304_x882_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:283:@88885.4]
  assign _T_961 = _T_960 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:292:@88886.4]
  assign x1305_x838_rdcol_D30_number = RetimeWrapper_65_io_out; // @[package.scala 96:25:@88902.4 package.scala 96:25:@88903.4]
  assign _T_972 = $signed(x1305_x838_rdcol_D30_number); // @[Math.scala 465:37:@88908.4]
  assign x886 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@88916.4 package.scala 96:25:@88917.4]
  assign x887 = x1289_x864_D1 | x886; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 394:25:@88920.4]
  assign _T_1004 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@88971.4 package.scala 96:25:@88972.4]
  assign _T_1006 = io_rr ? _T_1004 : 1'h0; // @[implicits.scala 55:10:@88973.4]
  assign _T_1007 = _T_387 & _T_1006; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:194:@88974.4]
  assign x1307_x888_D20 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@88950.4 package.scala 96:25:@88951.4]
  assign _T_1008 = _T_1007 & x1307_x888_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:283:@88975.4]
  assign _T_1009 = _T_1008 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:292:@88976.4]
  assign x1309_x832_rdcol_D30_number = RetimeWrapper_71_io_out; // @[package.scala 96:25:@88992.4 package.scala 96:25:@88993.4]
  assign _T_1022 = $signed(x1309_x832_rdcol_D30_number); // @[Math.scala 465:37:@89000.4]
  assign x892 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@89008.4 package.scala 96:25:@89009.4]
  assign x893 = x1289_x864_D1 | x892; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 425:60:@89012.4]
  assign _T_1054 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@89063.4 package.scala 96:25:@89064.4]
  assign _T_1056 = io_rr ? _T_1054 : 1'h0; // @[implicits.scala 55:10:@89065.4]
  assign _T_1057 = _T_387 & _T_1056; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:194:@89066.4]
  assign x1312_x894_D20 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@89051.4 package.scala 96:25:@89052.4]
  assign _T_1058 = _T_1057 & x1312_x894_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:283:@89067.4]
  assign _T_1059 = _T_1058 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:292:@89068.4]
  assign x1313_x826_rdcol_D30_number = RetimeWrapper_77_io_out; // @[package.scala 96:25:@89084.4 package.scala 96:25:@89085.4]
  assign _T_1070 = $signed(x1313_x826_rdcol_D30_number); // @[Math.scala 465:37:@89090.4]
  assign x898 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@89098.4 package.scala 96:25:@89099.4]
  assign x899 = x1289_x864_D1 | x898; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 448:60:@89102.4]
  assign _T_1102 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@89153.4 package.scala 96:25:@89154.4]
  assign _T_1104 = io_rr ? _T_1102 : 1'h0; // @[implicits.scala 55:10:@89155.4]
  assign _T_1105 = _T_387 & _T_1104; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:194:@89156.4]
  assign x1315_x900_D20 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@89132.4 package.scala 96:25:@89133.4]
  assign _T_1106 = _T_1105 & x1315_x900_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:283:@89157.4]
  assign _T_1107 = _T_1106 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:292:@89158.4]
  assign x1317_x820_rdcol_D30_number = RetimeWrapper_83_io_out; // @[package.scala 96:25:@89174.4 package.scala 96:25:@89175.4]
  assign _T_1118 = $signed(x1317_x820_rdcol_D30_number); // @[Math.scala 465:37:@89180.4]
  assign x904 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@89188.4 package.scala 96:25:@89189.4]
  assign x905 = x1289_x864_D1 | x904; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 471:60:@89192.4]
  assign _T_1150 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@89243.4 package.scala 96:25:@89244.4]
  assign _T_1152 = io_rr ? _T_1150 : 1'h0; // @[implicits.scala 55:10:@89245.4]
  assign _T_1153 = _T_387 & _T_1152; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:194:@89246.4]
  assign x1319_x906_D20 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@89222.4 package.scala 96:25:@89223.4]
  assign _T_1154 = _T_1153 & x1319_x906_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:283:@89247.4]
  assign _T_1155 = _T_1154 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:292:@89248.4]
  assign x1321_b800_D30_number = RetimeWrapper_89_io_out; // @[package.scala 96:25:@89264.4 package.scala 96:25:@89265.4]
  assign _T_1166 = $signed(x1321_b800_D30_number); // @[Math.scala 465:37:@89270.4]
  assign x864 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@88536.4 package.scala 96:25:@88537.4]
  assign x910 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@89278.4 package.scala 96:25:@89279.4]
  assign x911 = x864 | x910; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 494:59:@89282.4]
  assign _T_1204 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@89351.4 package.scala 96:25:@89352.4]
  assign _T_1206 = io_rr ? _T_1204 : 1'h0; // @[implicits.scala 55:10:@89353.4]
  assign _T_1207 = _T_387 & _T_1206; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:194:@89354.4]
  assign x1326_x912_D21 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@89339.4 package.scala 96:25:@89340.4]
  assign _T_1208 = _T_1207 & x1326_x912_D21; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:283:@89355.4]
  assign _T_1209 = _T_1208 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:292:@89356.4]
  assign x916_rdcol_number = x916_rdcol_1_io_result; // @[Math.scala 154:22:@89375.4 Math.scala 155:14:@89376.4]
  assign _T_1224 = $signed(x916_rdcol_number); // @[Math.scala 465:37:@89381.4]
  assign x917 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@89389.4 package.scala 96:25:@89390.4]
  assign x918 = x1289_x864_D1 | x917; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 521:60:@89393.4]
  assign _T_1267 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@89459.4 package.scala 96:25:@89460.4]
  assign _T_1269 = io_rr ? _T_1267 : 1'h0; // @[implicits.scala 55:10:@89461.4]
  assign _T_1270 = _T_387 & _T_1269; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:194:@89462.4]
  assign x1328_x919_D20 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@89447.4 package.scala 96:25:@89448.4]
  assign _T_1271 = _T_1270 & x1328_x919_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:283:@89463.4]
  assign _T_1272 = _T_1271 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:292:@89464.4]
  assign x925_rdcol_number = x925_rdcol_1_io_result; // @[Math.scala 154:22:@89485.4 Math.scala 155:14:@89486.4]
  assign _T_1289 = $signed(x925_rdcol_number); // @[Math.scala 465:37:@89491.4]
  assign x926 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@89499.4 package.scala 96:25:@89500.4]
  assign x927 = x1289_x864_D1 | x926; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 554:60:@89503.4]
  assign _T_1332 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@89569.4 package.scala 96:25:@89570.4]
  assign _T_1334 = io_rr ? _T_1332 : 1'h0; // @[implicits.scala 55:10:@89571.4]
  assign _T_1335 = _T_387 & _T_1334; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 571:194:@89572.4]
  assign x1330_x928_D20 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@89557.4 package.scala 96:25:@89558.4]
  assign _T_1336 = _T_1335 & x1330_x928_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 571:283:@89573.4]
  assign _T_1337 = _T_1336 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 571:292:@89574.4]
  assign x934_rdrow_number = x934_rdrow_1_io_result; // @[Math.scala 195:22:@89593.4 Math.scala 196:14:@89594.4]
  assign _T_1354 = $signed(x934_rdrow_number); // @[Math.scala 406:49:@89600.4]
  assign _T_1356 = $signed(_T_1354) & $signed(32'sh3); // @[Math.scala 406:56:@89602.4]
  assign _T_1357 = $signed(_T_1356); // @[Math.scala 406:56:@89603.4]
  assign _T_1361 = $signed(RetimeWrapper_105_io_out); // @[package.scala 96:25:@89611.4]
  assign x1241_number = $unsigned(_T_1361); // @[implicits.scala 133:21:@89613.4]
  assign x936 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@89627.4 package.scala 96:25:@89628.4]
  assign x937 = x936 | x865; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 581:24:@89631.4]
  assign _T_1384 = $signed(x1241_number); // @[Math.scala 406:49:@89640.4]
  assign _T_1386 = $signed(_T_1384) & $signed(32'sh3); // @[Math.scala 406:56:@89642.4]
  assign _T_1387 = $signed(_T_1386); // @[Math.scala 406:56:@89643.4]
  assign _T_1392 = x1241_number[31]; // @[FixedPoint.scala 50:25:@89649.4]
  assign _T_1396 = _T_1392 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@89651.4]
  assign _T_1397 = x1241_number[31:2]; // @[FixedPoint.scala 18:52:@89652.4]
  assign x940_number = {_T_1396,_T_1397}; // @[Cat.scala 30:58:@89653.4]
  assign _GEN_4 = {{7'd0}, x940_number}; // @[Math.scala 450:32:@89658.4]
  assign _T_1402 = _GEN_4 << 7; // @[Math.scala 450:32:@89658.4]
  assign _GEN_5 = {{6'd0}, x940_number}; // @[Math.scala 450:32:@89663.4]
  assign _T_1406 = _GEN_5 << 6; // @[Math.scala 450:32:@89663.4]
  assign _T_1433 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@89722.4 package.scala 96:25:@89723.4]
  assign _T_1435 = io_rr ? _T_1433 : 1'h0; // @[implicits.scala 55:10:@89724.4]
  assign _T_1436 = _T_387 & _T_1435; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:194:@89725.4]
  assign x1333_x938_D20 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@89710.4 package.scala 96:25:@89711.4]
  assign _T_1437 = _T_1436 & x1333_x938_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:283:@89726.4]
  assign _T_1438 = _T_1437 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:292:@89727.4]
  assign x945 = x936 | x874; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 610:24:@89738.4]
  assign _T_1462 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@89771.4 package.scala 96:25:@89772.4]
  assign _T_1464 = io_rr ? _T_1462 : 1'h0; // @[implicits.scala 55:10:@89773.4]
  assign _T_1465 = _T_387 & _T_1464; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:194:@89774.4]
  assign x1334_x946_D20 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@89759.4 package.scala 96:25:@89760.4]
  assign _T_1466 = _T_1465 & x1334_x946_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:283:@89775.4]
  assign _T_1467 = _T_1466 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:292:@89776.4]
  assign x950 = x936 | x880; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 625:24:@89787.4]
  assign _T_1491 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@89820.4 package.scala 96:25:@89821.4]
  assign _T_1493 = io_rr ? _T_1491 : 1'h0; // @[implicits.scala 55:10:@89822.4]
  assign _T_1494 = _T_387 & _T_1493; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:194:@89823.4]
  assign x1335_x951_D20 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@89808.4 package.scala 96:25:@89809.4]
  assign _T_1495 = _T_1494 & x1335_x951_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:283:@89824.4]
  assign _T_1496 = _T_1495 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:292:@89825.4]
  assign x955 = x936 | x886; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 640:24:@89836.4]
  assign _T_1520 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@89869.4 package.scala 96:25:@89870.4]
  assign _T_1522 = io_rr ? _T_1520 : 1'h0; // @[implicits.scala 55:10:@89871.4]
  assign _T_1523 = _T_387 & _T_1522; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:194:@89872.4]
  assign x1336_x956_D20 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@89857.4 package.scala 96:25:@89858.4]
  assign _T_1524 = _T_1523 & x1336_x956_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:283:@89873.4]
  assign _T_1525 = _T_1524 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:292:@89874.4]
  assign x960 = x936 | x892; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 655:24:@89885.4]
  assign _T_1551 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@89920.4 package.scala 96:25:@89921.4]
  assign _T_1553 = io_rr ? _T_1551 : 1'h0; // @[implicits.scala 55:10:@89922.4]
  assign _T_1554 = _T_387 & _T_1553; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:194:@89923.4]
  assign x1337_x961_D20 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@89908.4 package.scala 96:25:@89909.4]
  assign _T_1555 = _T_1554 & x1337_x961_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:283:@89924.4]
  assign _T_1556 = _T_1555 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:292:@89925.4]
  assign x965 = x936 | x898; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 678:59:@89936.4]
  assign _T_1580 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@89969.4 package.scala 96:25:@89970.4]
  assign _T_1582 = io_rr ? _T_1580 : 1'h0; // @[implicits.scala 55:10:@89971.4]
  assign _T_1583 = _T_387 & _T_1582; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:194:@89972.4]
  assign x1338_x966_D20 = RetimeWrapper_119_io_out; // @[package.scala 96:25:@89957.4 package.scala 96:25:@89958.4]
  assign _T_1584 = _T_1583 & x1338_x966_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:283:@89973.4]
  assign _T_1585 = _T_1584 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:292:@89974.4]
  assign x970 = x936 | x904; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 693:59:@89985.4]
  assign _T_1609 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@90018.4 package.scala 96:25:@90019.4]
  assign _T_1611 = io_rr ? _T_1609 : 1'h0; // @[implicits.scala 55:10:@90020.4]
  assign _T_1612 = _T_387 & _T_1611; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:194:@90021.4]
  assign x1339_x971_D20 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@90006.4 package.scala 96:25:@90007.4]
  assign _T_1613 = _T_1612 & x1339_x971_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:283:@90022.4]
  assign _T_1614 = _T_1613 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:292:@90023.4]
  assign x1340_x910_D1 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@90039.4 package.scala 96:25:@90040.4]
  assign x975 = x936 | x1340_x910_D1; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 710:59:@90043.4]
  assign _T_1647 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@90094.4 package.scala 96:25:@90095.4]
  assign _T_1649 = io_rr ? _T_1647 : 1'h0; // @[implicits.scala 55:10:@90096.4]
  assign _T_1650 = _T_387 & _T_1649; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:194:@90097.4]
  assign x1343_x976_D20 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@90082.4 package.scala 96:25:@90083.4]
  assign _T_1651 = _T_1650 & x1343_x976_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:283:@90098.4]
  assign _T_1652 = _T_1651 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:292:@90099.4]
  assign x980 = x936 | x917; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 729:59:@90110.4]
  assign _T_1676 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@90143.4 package.scala 96:25:@90144.4]
  assign _T_1678 = io_rr ? _T_1676 : 1'h0; // @[implicits.scala 55:10:@90145.4]
  assign _T_1679 = _T_387 & _T_1678; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:194:@90146.4]
  assign x1344_x981_D20 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@90131.4 package.scala 96:25:@90132.4]
  assign _T_1680 = _T_1679 & x1344_x981_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:283:@90147.4]
  assign _T_1681 = _T_1680 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:292:@90148.4]
  assign x985 = x936 | x926; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 744:59:@90159.4]
  assign _T_1705 = RetimeWrapper_131_io_out; // @[package.scala 96:25:@90192.4 package.scala 96:25:@90193.4]
  assign _T_1707 = io_rr ? _T_1705 : 1'h0; // @[implicits.scala 55:10:@90194.4]
  assign _T_1708 = _T_387 & _T_1707; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:194:@90195.4]
  assign x1345_x986_D20 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@90180.4 package.scala 96:25:@90181.4]
  assign _T_1709 = _T_1708 & x1345_x986_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:283:@90196.4]
  assign _T_1710 = _T_1709 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:292:@90197.4]
  assign x990_rdrow_number = x990_rdrow_1_io_result; // @[Math.scala 195:22:@90216.4 Math.scala 196:14:@90217.4]
  assign _T_1727 = $signed(x990_rdrow_number); // @[Math.scala 406:49:@90223.4]
  assign _T_1729 = $signed(_T_1727) & $signed(32'sh3); // @[Math.scala 406:56:@90225.4]
  assign _T_1730 = $signed(_T_1729); // @[Math.scala 406:56:@90226.4]
  assign _T_1734 = $signed(RetimeWrapper_132_io_out); // @[package.scala 96:25:@90234.4]
  assign x1246_number = $unsigned(_T_1734); // @[implicits.scala 133:21:@90236.4]
  assign x992 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@90250.4 package.scala 96:25:@90251.4]
  assign x993 = x992 | x865; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 765:24:@90254.4]
  assign _T_1757 = $signed(x1246_number); // @[Math.scala 406:49:@90263.4]
  assign _T_1759 = $signed(_T_1757) & $signed(32'sh3); // @[Math.scala 406:56:@90265.4]
  assign _T_1760 = $signed(_T_1759); // @[Math.scala 406:56:@90266.4]
  assign _T_1765 = x1246_number[31]; // @[FixedPoint.scala 50:25:@90272.4]
  assign _T_1769 = _T_1765 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@90274.4]
  assign _T_1770 = x1246_number[31:2]; // @[FixedPoint.scala 18:52:@90275.4]
  assign x996_number = {_T_1769,_T_1770}; // @[Cat.scala 30:58:@90276.4]
  assign _GEN_6 = {{7'd0}, x996_number}; // @[Math.scala 450:32:@90281.4]
  assign _T_1775 = _GEN_6 << 7; // @[Math.scala 450:32:@90281.4]
  assign _GEN_7 = {{6'd0}, x996_number}; // @[Math.scala 450:32:@90286.4]
  assign _T_1779 = _GEN_7 << 6; // @[Math.scala 450:32:@90286.4]
  assign _T_1808 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@90347.4 package.scala 96:25:@90348.4]
  assign _T_1810 = io_rr ? _T_1808 : 1'h0; // @[implicits.scala 55:10:@90349.4]
  assign _T_1811 = _T_387 & _T_1810; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 798:194:@90350.4]
  assign x1347_x994_D20 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@90326.4 package.scala 96:25:@90327.4]
  assign _T_1812 = _T_1811 & x1347_x994_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 798:283:@90351.4]
  assign _T_1813 = _T_1812 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 798:292:@90352.4]
  assign x1001 = x992 | x874; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 802:60:@90363.4]
  assign _T_1837 = RetimeWrapper_139_io_out; // @[package.scala 96:25:@90396.4 package.scala 96:25:@90397.4]
  assign _T_1839 = io_rr ? _T_1837 : 1'h0; // @[implicits.scala 55:10:@90398.4]
  assign _T_1840 = _T_387 & _T_1839; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:199:@90399.4]
  assign x1349_x1002_D20 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@90384.4 package.scala 96:25:@90385.4]
  assign _T_1841 = _T_1840 & x1349_x1002_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:288:@90400.4]
  assign _T_1842 = _T_1841 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:297:@90401.4]
  assign x1006 = x992 | x880; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 817:60:@90412.4]
  assign _T_1866 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@90445.4 package.scala 96:25:@90446.4]
  assign _T_1868 = io_rr ? _T_1866 : 1'h0; // @[implicits.scala 55:10:@90447.4]
  assign _T_1869 = _T_387 & _T_1868; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:199:@90448.4]
  assign x1350_x1007_D20 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@90433.4 package.scala 96:25:@90434.4]
  assign _T_1870 = _T_1869 & x1350_x1007_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:288:@90449.4]
  assign _T_1871 = _T_1870 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:297:@90450.4]
  assign x1011 = x992 | x886; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 832:60:@90461.4]
  assign _T_1895 = RetimeWrapper_143_io_out; // @[package.scala 96:25:@90494.4 package.scala 96:25:@90495.4]
  assign _T_1897 = io_rr ? _T_1895 : 1'h0; // @[implicits.scala 55:10:@90496.4]
  assign _T_1898 = _T_387 & _T_1897; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:199:@90497.4]
  assign x1351_x1012_D20 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@90482.4 package.scala 96:25:@90483.4]
  assign _T_1899 = _T_1898 & x1351_x1012_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:288:@90498.4]
  assign _T_1900 = _T_1899 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:297:@90499.4]
  assign x1016 = x992 | x892; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 847:60:@90510.4]
  assign _T_1924 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@90543.4 package.scala 96:25:@90544.4]
  assign _T_1926 = io_rr ? _T_1924 : 1'h0; // @[implicits.scala 55:10:@90545.4]
  assign _T_1927 = _T_387 & _T_1926; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:199:@90546.4]
  assign x1352_x1017_D20 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@90531.4 package.scala 96:25:@90532.4]
  assign _T_1928 = _T_1927 & x1352_x1017_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:288:@90547.4]
  assign _T_1929 = _T_1928 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:297:@90548.4]
  assign x1021 = x992 | x898; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 862:60:@90559.4]
  assign _T_1953 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@90592.4 package.scala 96:25:@90593.4]
  assign _T_1955 = io_rr ? _T_1953 : 1'h0; // @[implicits.scala 55:10:@90594.4]
  assign _T_1956 = _T_387 & _T_1955; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:199:@90595.4]
  assign x1353_x1022_D20 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@90580.4 package.scala 96:25:@90581.4]
  assign _T_1957 = _T_1956 & x1353_x1022_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:288:@90596.4]
  assign _T_1958 = _T_1957 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:297:@90597.4]
  assign x1026 = x992 | x904; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 877:60:@90608.4]
  assign _T_1982 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@90641.4 package.scala 96:25:@90642.4]
  assign _T_1984 = io_rr ? _T_1982 : 1'h0; // @[implicits.scala 55:10:@90643.4]
  assign _T_1985 = _T_387 & _T_1984; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:199:@90644.4]
  assign x1354_x1027_D20 = RetimeWrapper_148_io_out; // @[package.scala 96:25:@90629.4 package.scala 96:25:@90630.4]
  assign _T_1986 = _T_1985 & x1354_x1027_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:288:@90645.4]
  assign _T_1987 = _T_1986 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:297:@90646.4]
  assign x1031 = x992 | x1340_x910_D1; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 892:60:@90657.4]
  assign _T_2017 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@90708.4 package.scala 96:25:@90709.4]
  assign _T_2019 = io_rr ? _T_2017 : 1'h0; // @[implicits.scala 55:10:@90710.4]
  assign _T_2020 = _T_387 & _T_2019; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:199:@90711.4]
  assign x1356_x1032_D20 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@90687.4 package.scala 96:25:@90688.4]
  assign _T_2021 = _T_2020 & x1356_x1032_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:288:@90712.4]
  assign _T_2022 = _T_2021 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:297:@90713.4]
  assign x1036 = x992 | x917; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 917:60:@90724.4]
  assign _T_2048 = RetimeWrapper_155_io_out; // @[package.scala 96:25:@90759.4 package.scala 96:25:@90760.4]
  assign _T_2050 = io_rr ? _T_2048 : 1'h0; // @[implicits.scala 55:10:@90761.4]
  assign _T_2051 = _T_387 & _T_2050; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:199:@90762.4]
  assign x1358_x1037_D20 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@90747.4 package.scala 96:25:@90748.4]
  assign _T_2052 = _T_2051 & x1358_x1037_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:288:@90763.4]
  assign _T_2053 = _T_2052 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:297:@90764.4]
  assign x1041 = x992 | x926; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 934:60:@90775.4]
  assign _T_2077 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@90808.4 package.scala 96:25:@90809.4]
  assign _T_2079 = io_rr ? _T_2077 : 1'h0; // @[implicits.scala 55:10:@90810.4]
  assign _T_2080 = _T_387 & _T_2079; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 945:199:@90811.4]
  assign x1359_x1042_D20 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@90796.4 package.scala 96:25:@90797.4]
  assign _T_2081 = _T_2080 & x1359_x1042_D20; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 945:288:@90812.4]
  assign _T_2082 = _T_2081 & x1296_b801_D52; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 945:297:@90813.4]
  assign x878_rd_0_number = x805_lb_0_io_rPort_1_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 359:29:@88782.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 363:341:@88803.4]
  assign _GEN_8 = {{1'd0}, x878_rd_0_number}; // @[Math.scala 450:32:@90825.4]
  assign x943_rd_0_number = x805_lb_0_io_rPort_12_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 602:29:@89713.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 606:411:@89734.4]
  assign _GEN_9 = {{1'd0}, x943_rd_0_number}; // @[Math.scala 450:32:@90837.4]
  assign x948_rd_0_number = x805_lb_0_io_rPort_5_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 617:29:@89762.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 621:411:@89783.4]
  assign _GEN_10 = {{2'd0}, x948_rd_0_number}; // @[Math.scala 450:32:@90849.4]
  assign x953_rd_0_number = x805_lb_0_io_rPort_8_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 632:29:@89811.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 636:411:@89832.4]
  assign _GEN_11 = {{1'd0}, x953_rd_0_number}; // @[Math.scala 450:32:@90861.4]
  assign x1004_rd_0_number = x805_lb_0_io_rPort_26_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 809:30:@90387.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 813:416:@90408.4]
  assign _GEN_12 = {{1'd0}, x1004_rd_0_number}; // @[Math.scala 450:32:@90873.4]
  assign x1058_sum_number = x1058_sum_1_io_result; // @[Math.scala 154:22:@90996.4 Math.scala 155:14:@90997.4]
  assign _T_2159 = x1058_sum_number[7:4]; // @[FixedPoint.scala 18:52:@91002.4]
  assign x884_rd_0_number = x805_lb_0_io_rPort_6_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 382:29:@88872.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 386:341:@88893.4]
  assign _GEN_13 = {{1'd0}, x884_rd_0_number}; // @[Math.scala 450:32:@91008.4]
  assign _GEN_14 = {{1'd0}, x948_rd_0_number}; // @[Math.scala 450:32:@91020.4]
  assign _GEN_15 = {{2'd0}, x953_rd_0_number}; // @[Math.scala 450:32:@91032.4]
  assign x958_rd_0_number = x805_lb_0_io_rPort_9_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 647:29:@89860.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 651:411:@89881.4]
  assign _GEN_16 = {{1'd0}, x958_rd_0_number}; // @[Math.scala 450:32:@91044.4]
  assign x1009_rd_0_number = x805_lb_0_io_rPort_27_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 824:30:@90436.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 828:416:@90457.4]
  assign _GEN_17 = {{1'd0}, x1009_rd_0_number}; // @[Math.scala 450:32:@91056.4]
  assign x1072_sum_number = x1072_sum_1_io_result; // @[Math.scala 154:22:@91179.4 Math.scala 155:14:@91180.4]
  assign _T_2235 = x1072_sum_number[7:4]; // @[FixedPoint.scala 18:52:@91185.4]
  assign x890_rd_0_number = x805_lb_0_io_rPort_10_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 405:29:@88962.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 409:341:@88983.4]
  assign _GEN_18 = {{1'd0}, x890_rd_0_number}; // @[Math.scala 450:32:@91191.4]
  assign _GEN_19 = {{2'd0}, x958_rd_0_number}; // @[Math.scala 450:32:@91205.4]
  assign x963_rd_0_number = x805_lb_0_io_rPort_20_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 670:29:@89911.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 674:411:@89932.4]
  assign _GEN_20 = {{1'd0}, x963_rd_0_number}; // @[Math.scala 450:32:@91217.4]
  assign x1014_rd_0_number = x805_lb_0_io_rPort_29_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 839:30:@90485.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 843:416:@90506.4]
  assign _GEN_21 = {{1'd0}, x1014_rd_0_number}; // @[Math.scala 450:32:@91229.4]
  assign x1085_sum_number = x1085_sum_1_io_result; // @[Math.scala 154:22:@91334.4 Math.scala 155:14:@91335.4]
  assign _T_2301 = x1085_sum_number[7:4]; // @[FixedPoint.scala 18:52:@91340.4]
  assign x896_rd_0_number = x805_lb_0_io_rPort_21_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 436:29:@89054.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 440:411:@89075.4]
  assign _GEN_22 = {{1'd0}, x896_rd_0_number}; // @[Math.scala 450:32:@91346.4]
  assign _GEN_23 = {{2'd0}, x963_rd_0_number}; // @[Math.scala 450:32:@91358.4]
  assign x968_rd_0_number = x805_lb_0_io_rPort_17_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 685:29:@89960.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 689:411:@89981.4]
  assign _GEN_24 = {{1'd0}, x968_rd_0_number}; // @[Math.scala 450:32:@91370.4]
  assign x1019_rd_0_number = x805_lb_0_io_rPort_24_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 854:30:@90534.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 858:416:@90555.4]
  assign _GEN_25 = {{1'd0}, x1019_rd_0_number}; // @[Math.scala 450:32:@91382.4]
  assign x1098_sum_number = x1098_sum_1_io_result; // @[Math.scala 154:22:@91487.4 Math.scala 155:14:@91488.4]
  assign _T_2365 = x1098_sum_number[7:4]; // @[FixedPoint.scala 18:52:@91493.4]
  assign x902_rd_0_number = x805_lb_0_io_rPort_3_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 459:29:@89144.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 463:411:@89165.4]
  assign _GEN_26 = {{1'd0}, x902_rd_0_number}; // @[Math.scala 450:32:@91499.4]
  assign _GEN_27 = {{2'd0}, x968_rd_0_number}; // @[Math.scala 450:32:@91511.4]
  assign x973_rd_0_number = x805_lb_0_io_rPort_2_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 700:29:@90009.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 704:411:@90030.4]
  assign _GEN_28 = {{1'd0}, x973_rd_0_number}; // @[Math.scala 450:32:@91523.4]
  assign x1024_rd_0_number = x805_lb_0_io_rPort_0_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 869:30:@90583.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 873:416:@90604.4]
  assign _GEN_29 = {{1'd0}, x1024_rd_0_number}; // @[Math.scala 450:32:@91535.4]
  assign x1111_sum_number = x1111_sum_1_io_result; // @[Math.scala 154:22:@91640.4 Math.scala 155:14:@91641.4]
  assign _T_2429 = x1111_sum_number[7:4]; // @[FixedPoint.scala 18:52:@91646.4]
  assign x908_rd_0_number = x805_lb_0_io_rPort_25_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 482:29:@89234.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 486:411:@89255.4]
  assign _GEN_30 = {{1'd0}, x908_rd_0_number}; // @[Math.scala 450:32:@91652.4]
  assign _GEN_31 = {{2'd0}, x973_rd_0_number}; // @[Math.scala 450:32:@91664.4]
  assign x978_rd_0_number = x805_lb_0_io_rPort_19_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 721:29:@90085.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 725:411:@90106.4]
  assign _GEN_32 = {{1'd0}, x978_rd_0_number}; // @[Math.scala 450:32:@91676.4]
  assign x1029_rd_0_number = x805_lb_0_io_rPort_11_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 884:30:@90632.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 888:416:@90653.4]
  assign _GEN_33 = {{1'd0}, x1029_rd_0_number}; // @[Math.scala 450:32:@91688.4]
  assign x1124_sum_number = x1124_sum_1_io_result; // @[Math.scala 154:22:@91795.4 Math.scala 155:14:@91796.4]
  assign _T_2495 = x1124_sum_number[7:4]; // @[FixedPoint.scala 18:52:@91801.4]
  assign x914_rd_0_number = x805_lb_0_io_rPort_22_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 509:29:@89342.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 513:411:@89363.4]
  assign _GEN_34 = {{1'd0}, x914_rd_0_number}; // @[Math.scala 450:32:@91807.4]
  assign _GEN_35 = {{2'd0}, x978_rd_0_number}; // @[Math.scala 450:32:@91819.4]
  assign x983_rd_0_number = x805_lb_0_io_rPort_14_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 736:29:@90134.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 740:411:@90155.4]
  assign _GEN_36 = {{1'd0}, x983_rd_0_number}; // @[Math.scala 450:32:@91831.4]
  assign x1034_rd_0_number = x805_lb_0_io_rPort_16_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 903:30:@90699.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 907:416:@90720.4]
  assign _GEN_37 = {{1'd0}, x1034_rd_0_number}; // @[Math.scala 450:32:@91843.4]
  assign x1137_sum_number = x1137_sum_1_io_result; // @[Math.scala 154:22:@91948.4 Math.scala 155:14:@91949.4]
  assign _T_2559 = x1137_sum_number[7:4]; // @[FixedPoint.scala 18:52:@91954.4]
  assign x923_rd_0_number = x805_lb_0_io_rPort_28_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 540:29:@89450.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 544:411:@89471.4]
  assign _GEN_38 = {{1'd0}, x923_rd_0_number}; // @[Math.scala 450:32:@91960.4]
  assign _GEN_39 = {{2'd0}, x983_rd_0_number}; // @[Math.scala 450:32:@91972.4]
  assign x988_rd_0_number = x805_lb_0_io_rPort_4_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 751:29:@90183.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 755:411:@90204.4]
  assign _GEN_40 = {{1'd0}, x988_rd_0_number}; // @[Math.scala 450:32:@91984.4]
  assign x1039_rd_0_number = x805_lb_0_io_rPort_7_output_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 926:30:@90750.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 930:416:@90771.4]
  assign _GEN_41 = {{1'd0}, x1039_rd_0_number}; // @[Math.scala 450:32:@91996.4]
  assign x1150_sum_number = x1150_sum_1_io_result; // @[Math.scala 154:22:@92101.4 Math.scala 155:14:@92102.4]
  assign _T_2623 = x1150_sum_number[7:4]; // @[FixedPoint.scala 18:52:@92107.4]
  assign _T_2642 = {4'h0,_T_2429,4'h0,_T_2495,4'h0,_T_2559,4'h0,_T_2623}; // @[Cat.scala 30:58:@92123.4]
  assign _T_2645 = {4'h0,_T_2159,4'h0,_T_2235,4'h0,_T_2301,4'h0,_T_2365}; // @[Cat.scala 30:58:@92126.4]
  assign _T_2658 = RetimeWrapper_215_io_out; // @[package.scala 96:25:@92162.4 package.scala 96:25:@92163.4]
  assign _T_2660 = io_rr ? _T_2658 : 1'h0; // @[implicits.scala 55:10:@92164.4]
  assign x1380_b801_D59 = RetimeWrapper_213_io_out; // @[package.scala 96:25:@92144.4 package.scala 96:25:@92145.4]
  assign _T_2661 = _T_2660 & x1380_b801_D59; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1225:117:@92165.4]
  assign x1381_b802_D59 = RetimeWrapper_214_io_out; // @[package.scala 96:25:@92153.4 package.scala 96:25:@92154.4]
  assign _T_2662 = _T_2661 & x1381_b802_D59; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1225:124:@92166.4]
  assign x1259_x814_D12_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@87728.4 package.scala 96:25:@87729.4]
  assign x1261_x1232_D26_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@87746.4 package.scala 96:25:@87747.4]
  assign x1263_x818_sum_D7_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@87764.4 package.scala 96:25:@87765.4]
  assign x1267_x824_sum_D6_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@87871.4 package.scala 96:25:@87872.4]
  assign x1268_x822_D11_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@87880.4 package.scala 96:25:@87881.4]
  assign x1269_x830_sum_D6_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@87960.4 package.scala 96:25:@87961.4]
  assign x1271_x828_D11_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@87978.4 package.scala 96:25:@87979.4]
  assign x1272_x834_D11_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@88060.4 package.scala 96:25:@88061.4]
  assign x1273_x836_sum_D6_number = RetimeWrapper_20_io_out; // @[package.scala 96:25:@88069.4 package.scala 96:25:@88070.4]
  assign x1275_x842_sum_D6_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@88158.4 package.scala 96:25:@88159.4]
  assign x1276_x840_D11_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@88167.4 package.scala 96:25:@88168.4]
  assign x1278_x846_D11_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@88256.4 package.scala 96:25:@88257.4]
  assign x1279_x848_sum_D6_number = RetimeWrapper_28_io_out; // @[package.scala 96:25:@88265.4 package.scala 96:25:@88266.4]
  assign x1281_x852_D11_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@88354.4 package.scala 96:25:@88355.4]
  assign x1283_x854_sum_D6_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@88372.4 package.scala 96:25:@88373.4]
  assign x1285_x858_D11_number = RetimeWrapper_36_io_out; // @[package.scala 96:25:@88461.4 package.scala 96:25:@88462.4]
  assign x1286_x860_sum_D6_number = RetimeWrapper_37_io_out; // @[package.scala 96:25:@88470.4 package.scala 96:25:@88471.4]
  assign x871_sum_number = x871_sum_1_io_result; // @[Math.scala 154:22:@88644.4 Math.scala 155:14:@88645.4]
  assign x1292_x1237_D21_number = RetimeWrapper_47_io_out; // @[package.scala 96:25:@88653.4 package.scala 96:25:@88654.4]
  assign x1294_x858_D35_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@88671.4 package.scala 96:25:@88672.4]
  assign x877_sum_number = x877_sum_1_io_result; // @[Math.scala 154:22:@88761.4 Math.scala 155:14:@88762.4]
  assign x1299_x852_D35_number = RetimeWrapper_56_io_out; // @[package.scala 96:25:@88770.4 package.scala 96:25:@88771.4]
  assign x883_sum_number = x883_sum_1_io_result; // @[Math.scala 154:22:@88851.4 Math.scala 155:14:@88852.4]
  assign x1303_x846_D35_number = RetimeWrapper_62_io_out; // @[package.scala 96:25:@88860.4 package.scala 96:25:@88861.4]
  assign x889_sum_number = x889_sum_1_io_result; // @[Math.scala 154:22:@88941.4 Math.scala 155:14:@88942.4]
  assign x1308_x840_D35_number = RetimeWrapper_69_io_out; // @[package.scala 96:25:@88959.4 package.scala 96:25:@88960.4]
  assign x895_sum_number = x895_sum_1_io_result; // @[Math.scala 154:22:@89033.4 Math.scala 155:14:@89034.4]
  assign x1311_x834_D35_number = RetimeWrapper_74_io_out; // @[package.scala 96:25:@89042.4 package.scala 96:25:@89043.4]
  assign x901_sum_number = x901_sum_1_io_result; // @[Math.scala 154:22:@89123.4 Math.scala 155:14:@89124.4]
  assign x1316_x828_D35_number = RetimeWrapper_81_io_out; // @[package.scala 96:25:@89141.4 package.scala 96:25:@89142.4]
  assign x907_sum_number = x907_sum_1_io_result; // @[Math.scala 154:22:@89213.4 Math.scala 155:14:@89214.4]
  assign x1320_x822_D35_number = RetimeWrapper_87_io_out; // @[package.scala 96:25:@89231.4 package.scala 96:25:@89232.4]
  assign x1324_x814_D36_number = RetimeWrapper_93_io_out; // @[package.scala 96:25:@89321.4 package.scala 96:25:@89322.4]
  assign x1325_x913_sum_D1_number = RetimeWrapper_94_io_out; // @[package.scala 96:25:@89330.4 package.scala 96:25:@89331.4]
  assign x922_sum_number = x922_sum_1_io_result; // @[Math.scala 154:22:@89429.4 Math.scala 155:14:@89430.4]
  assign x1327_x920_D5_number = RetimeWrapper_98_io_out; // @[package.scala 96:25:@89438.4 package.scala 96:25:@89439.4]
  assign x931_sum_number = x931_sum_1_io_result; // @[Math.scala 154:22:@89539.4 Math.scala 155:14:@89540.4]
  assign x1329_x929_D5_number = RetimeWrapper_102_io_out; // @[package.scala 96:25:@89548.4 package.scala 96:25:@89549.4]
  assign x942_sum_number = x942_sum_1_io_result; // @[Math.scala 154:22:@89692.4 Math.scala 155:14:@89693.4]
  assign x1332_x1242_D20_number = RetimeWrapper_108_io_out; // @[package.scala 96:25:@89701.4 package.scala 96:25:@89702.4]
  assign x947_sum_number = x947_sum_1_io_result; // @[Math.scala 154:22:@89750.4 Math.scala 155:14:@89751.4]
  assign x952_sum_number = x952_sum_1_io_result; // @[Math.scala 154:22:@89799.4 Math.scala 155:14:@89800.4]
  assign x957_sum_number = x957_sum_1_io_result; // @[Math.scala 154:22:@89848.4 Math.scala 155:14:@89849.4]
  assign x962_sum_number = x962_sum_1_io_result; // @[Math.scala 154:22:@89899.4 Math.scala 155:14:@89900.4]
  assign x967_sum_number = x967_sum_1_io_result; // @[Math.scala 154:22:@89948.4 Math.scala 155:14:@89949.4]
  assign x972_sum_number = x972_sum_1_io_result; // @[Math.scala 154:22:@89997.4 Math.scala 155:14:@89998.4]
  assign x1342_x977_sum_D1_number = RetimeWrapper_125_io_out; // @[package.scala 96:25:@90073.4 package.scala 96:25:@90074.4]
  assign x982_sum_number = x982_sum_1_io_result; // @[Math.scala 154:22:@90122.4 Math.scala 155:14:@90123.4]
  assign x987_sum_number = x987_sum_1_io_result; // @[Math.scala 154:22:@90171.4 Math.scala 155:14:@90172.4]
  assign x998_sum_number = x998_sum_1_io_result; // @[Math.scala 154:22:@90317.4 Math.scala 155:14:@90318.4]
  assign x1348_x1247_D20_number = RetimeWrapper_136_io_out; // @[package.scala 96:25:@90335.4 package.scala 96:25:@90336.4]
  assign x1003_sum_number = x1003_sum_1_io_result; // @[Math.scala 154:22:@90375.4 Math.scala 155:14:@90376.4]
  assign x1008_sum_number = x1008_sum_1_io_result; // @[Math.scala 154:22:@90424.4 Math.scala 155:14:@90425.4]
  assign x1013_sum_number = x1013_sum_1_io_result; // @[Math.scala 154:22:@90473.4 Math.scala 155:14:@90474.4]
  assign x1018_sum_number = x1018_sum_1_io_result; // @[Math.scala 154:22:@90522.4 Math.scala 155:14:@90523.4]
  assign x1023_sum_number = x1023_sum_1_io_result; // @[Math.scala 154:22:@90571.4 Math.scala 155:14:@90572.4]
  assign x1028_sum_number = x1028_sum_1_io_result; // @[Math.scala 154:22:@90620.4 Math.scala 155:14:@90621.4]
  assign x1357_x1033_sum_D1_number = RetimeWrapper_152_io_out; // @[package.scala 96:25:@90696.4 package.scala 96:25:@90697.4]
  assign x1038_sum_number = x1038_sum_1_io_result; // @[Math.scala 154:22:@90738.4 Math.scala 155:14:@90739.4]
  assign x1043_sum_number = x1043_sum_1_io_result; // @[Math.scala 154:22:@90787.4 Math.scala 155:14:@90788.4]
  assign _T_2090 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@90831.4 package.scala 96:25:@90832.4]
  assign _T_2096 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@90843.4 package.scala 96:25:@90844.4]
  assign _T_2102 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@90855.4 package.scala 96:25:@90856.4]
  assign _T_2108 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@90867.4 package.scala 96:25:@90868.4]
  assign _T_2114 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@90879.4 package.scala 96:25:@90880.4]
  assign _T_2166 = RetimeWrapper_167_io_out; // @[package.scala 96:25:@91014.4 package.scala 96:25:@91015.4]
  assign _T_2172 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@91026.4 package.scala 96:25:@91027.4]
  assign _T_2178 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@91038.4 package.scala 96:25:@91039.4]
  assign _T_2184 = RetimeWrapper_170_io_out; // @[package.scala 96:25:@91050.4 package.scala 96:25:@91051.4]
  assign _T_2190 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@91062.4 package.scala 96:25:@91063.4]
  assign _T_2242 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@91197.4 package.scala 96:25:@91198.4]
  assign _T_2250 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@91211.4 package.scala 96:25:@91212.4]
  assign _T_2256 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@91223.4 package.scala 96:25:@91224.4]
  assign _T_2262 = RetimeWrapper_179_io_out; // @[package.scala 96:25:@91235.4 package.scala 96:25:@91236.4]
  assign _T_2308 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@91352.4 package.scala 96:25:@91353.4]
  assign _T_2314 = RetimeWrapper_183_io_out; // @[package.scala 96:25:@91364.4 package.scala 96:25:@91365.4]
  assign _T_2320 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@91376.4 package.scala 96:25:@91377.4]
  assign _T_2326 = RetimeWrapper_185_io_out; // @[package.scala 96:25:@91388.4 package.scala 96:25:@91389.4]
  assign _T_2372 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@91505.4 package.scala 96:25:@91506.4]
  assign _T_2378 = RetimeWrapper_189_io_out; // @[package.scala 96:25:@91517.4 package.scala 96:25:@91518.4]
  assign _T_2384 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@91529.4 package.scala 96:25:@91530.4]
  assign _T_2390 = RetimeWrapper_191_io_out; // @[package.scala 96:25:@91541.4 package.scala 96:25:@91542.4]
  assign _T_2436 = RetimeWrapper_194_io_out; // @[package.scala 96:25:@91658.4 package.scala 96:25:@91659.4]
  assign _T_2442 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@91670.4 package.scala 96:25:@91671.4]
  assign _T_2448 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@91682.4 package.scala 96:25:@91683.4]
  assign _T_2454 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@91694.4 package.scala 96:25:@91695.4]
  assign _T_2502 = RetimeWrapper_200_io_out; // @[package.scala 96:25:@91813.4 package.scala 96:25:@91814.4]
  assign _T_2508 = RetimeWrapper_201_io_out; // @[package.scala 96:25:@91825.4 package.scala 96:25:@91826.4]
  assign _T_2514 = RetimeWrapper_202_io_out; // @[package.scala 96:25:@91837.4 package.scala 96:25:@91838.4]
  assign _T_2520 = RetimeWrapper_203_io_out; // @[package.scala 96:25:@91849.4 package.scala 96:25:@91850.4]
  assign _T_2566 = RetimeWrapper_206_io_out; // @[package.scala 96:25:@91966.4 package.scala 96:25:@91967.4]
  assign _T_2572 = RetimeWrapper_207_io_out; // @[package.scala 96:25:@91978.4 package.scala 96:25:@91979.4]
  assign _T_2578 = RetimeWrapper_208_io_out; // @[package.scala 96:25:@91990.4 package.scala 96:25:@91991.4]
  assign _T_2584 = RetimeWrapper_209_io_out; // @[package.scala 96:25:@92002.4 package.scala 96:25:@92003.4]
  assign io_in_x745_TVALID = _T_2662 & io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1225:22:@92168.4]
  assign io_in_x745_TDATA = {{192'd0}, RetimeWrapper_212_io_out}; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1226:24:@92169.4]
  assign io_in_x744_TREADY = _T_211 & _T_213; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 67:22:@87293.4 sm_x1156_inr_Foreach_SAMPLER_BOX.scala 69:22:@87301.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@87271.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@87283.4]
  assign RetimeWrapper_clock = clock; // @[:@87304.4]
  assign RetimeWrapper_reset = reset; // @[:@87305.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87307.4]
  assign RetimeWrapper_io_in = io_in_x744_TDATA[63:0]; // @[package.scala 94:16:@87306.4]
  assign x805_lb_0_clock = clock; // @[:@87314.4]
  assign x805_lb_0_reset = reset; // @[:@87315.4]
  assign x805_lb_0_io_rPort_29_banks_1 = x1308_x840_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90502.4]
  assign x805_lb_0_io_rPort_29_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90501.4]
  assign x805_lb_0_io_rPort_29_ofs_0 = x1013_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90503.4]
  assign x805_lb_0_io_rPort_29_en_0 = _T_1900 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90505.4]
  assign x805_lb_0_io_rPort_29_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90504.4]
  assign x805_lb_0_io_rPort_28_banks_1 = x1327_x920_D5_number[3:0]; // @[MemInterfaceType.scala 106:58:@89467.4]
  assign x805_lb_0_io_rPort_28_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@89466.4]
  assign x805_lb_0_io_rPort_28_ofs_0 = x922_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89468.4]
  assign x805_lb_0_io_rPort_28_en_0 = _T_1272 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89470.4]
  assign x805_lb_0_io_rPort_28_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89469.4]
  assign x805_lb_0_io_rPort_27_banks_1 = x1303_x846_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90453.4]
  assign x805_lb_0_io_rPort_27_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90452.4]
  assign x805_lb_0_io_rPort_27_ofs_0 = x1008_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90454.4]
  assign x805_lb_0_io_rPort_27_en_0 = _T_1871 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90456.4]
  assign x805_lb_0_io_rPort_27_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90455.4]
  assign x805_lb_0_io_rPort_26_banks_1 = x1299_x852_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90404.4]
  assign x805_lb_0_io_rPort_26_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90403.4]
  assign x805_lb_0_io_rPort_26_ofs_0 = x1003_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90405.4]
  assign x805_lb_0_io_rPort_26_en_0 = _T_1842 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90407.4]
  assign x805_lb_0_io_rPort_26_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90406.4]
  assign x805_lb_0_io_rPort_25_banks_1 = x1320_x822_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89251.4]
  assign x805_lb_0_io_rPort_25_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@89250.4]
  assign x805_lb_0_io_rPort_25_ofs_0 = x907_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89252.4]
  assign x805_lb_0_io_rPort_25_en_0 = _T_1155 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89254.4]
  assign x805_lb_0_io_rPort_25_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89253.4]
  assign x805_lb_0_io_rPort_24_banks_1 = x1311_x834_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90551.4]
  assign x805_lb_0_io_rPort_24_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90550.4]
  assign x805_lb_0_io_rPort_24_ofs_0 = x1018_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90552.4]
  assign x805_lb_0_io_rPort_24_en_0 = _T_1929 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90554.4]
  assign x805_lb_0_io_rPort_24_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90553.4]
  assign x805_lb_0_io_rPort_23_banks_1 = x1294_x858_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90355.4]
  assign x805_lb_0_io_rPort_23_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90354.4]
  assign x805_lb_0_io_rPort_23_ofs_0 = x998_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90356.4]
  assign x805_lb_0_io_rPort_23_en_0 = _T_1813 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90358.4]
  assign x805_lb_0_io_rPort_23_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90357.4]
  assign x805_lb_0_io_rPort_22_banks_1 = x1324_x814_D36_number[3:0]; // @[MemInterfaceType.scala 106:58:@89359.4]
  assign x805_lb_0_io_rPort_22_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@89358.4]
  assign x805_lb_0_io_rPort_22_ofs_0 = x1325_x913_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@89360.4]
  assign x805_lb_0_io_rPort_22_en_0 = _T_1209 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89362.4]
  assign x805_lb_0_io_rPort_22_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89361.4]
  assign x805_lb_0_io_rPort_21_banks_1 = x1311_x834_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89071.4]
  assign x805_lb_0_io_rPort_21_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@89070.4]
  assign x805_lb_0_io_rPort_21_ofs_0 = x895_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89072.4]
  assign x805_lb_0_io_rPort_21_en_0 = _T_1059 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89074.4]
  assign x805_lb_0_io_rPort_21_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89073.4]
  assign x805_lb_0_io_rPort_20_banks_1 = x1311_x834_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89928.4]
  assign x805_lb_0_io_rPort_20_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@89927.4]
  assign x805_lb_0_io_rPort_20_ofs_0 = x962_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89929.4]
  assign x805_lb_0_io_rPort_20_en_0 = _T_1556 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89931.4]
  assign x805_lb_0_io_rPort_20_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89930.4]
  assign x805_lb_0_io_rPort_19_banks_1 = x1324_x814_D36_number[3:0]; // @[MemInterfaceType.scala 106:58:@90102.4]
  assign x805_lb_0_io_rPort_19_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90101.4]
  assign x805_lb_0_io_rPort_19_ofs_0 = x1342_x977_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@90103.4]
  assign x805_lb_0_io_rPort_19_en_0 = _T_1652 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90105.4]
  assign x805_lb_0_io_rPort_19_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90104.4]
  assign x805_lb_0_io_rPort_18_banks_1 = x1294_x858_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@88709.4]
  assign x805_lb_0_io_rPort_18_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@88708.4]
  assign x805_lb_0_io_rPort_18_ofs_0 = x871_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@88710.4]
  assign x805_lb_0_io_rPort_18_en_0 = _T_865 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@88712.4]
  assign x805_lb_0_io_rPort_18_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@88711.4]
  assign x805_lb_0_io_rPort_17_banks_1 = x1316_x828_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89977.4]
  assign x805_lb_0_io_rPort_17_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@89976.4]
  assign x805_lb_0_io_rPort_17_ofs_0 = x967_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89978.4]
  assign x805_lb_0_io_rPort_17_en_0 = _T_1585 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89980.4]
  assign x805_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89979.4]
  assign x805_lb_0_io_rPort_16_banks_1 = x1324_x814_D36_number[3:0]; // @[MemInterfaceType.scala 106:58:@90716.4]
  assign x805_lb_0_io_rPort_16_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90715.4]
  assign x805_lb_0_io_rPort_16_ofs_0 = x1357_x1033_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@90717.4]
  assign x805_lb_0_io_rPort_16_en_0 = _T_2022 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90719.4]
  assign x805_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90718.4]
  assign x805_lb_0_io_rPort_15_banks_1 = x1329_x929_D5_number[3:0]; // @[MemInterfaceType.scala 106:58:@90816.4]
  assign x805_lb_0_io_rPort_15_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90815.4]
  assign x805_lb_0_io_rPort_15_ofs_0 = x1043_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90817.4]
  assign x805_lb_0_io_rPort_15_en_0 = _T_2082 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90819.4]
  assign x805_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90818.4]
  assign x805_lb_0_io_rPort_14_banks_1 = x1327_x920_D5_number[3:0]; // @[MemInterfaceType.scala 106:58:@90151.4]
  assign x805_lb_0_io_rPort_14_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90150.4]
  assign x805_lb_0_io_rPort_14_ofs_0 = x982_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90152.4]
  assign x805_lb_0_io_rPort_14_en_0 = _T_1681 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90154.4]
  assign x805_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90153.4]
  assign x805_lb_0_io_rPort_13_banks_1 = x1329_x929_D5_number[3:0]; // @[MemInterfaceType.scala 106:58:@89577.4]
  assign x805_lb_0_io_rPort_13_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@89576.4]
  assign x805_lb_0_io_rPort_13_ofs_0 = x931_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89578.4]
  assign x805_lb_0_io_rPort_13_en_0 = _T_1337 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89580.4]
  assign x805_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89579.4]
  assign x805_lb_0_io_rPort_12_banks_1 = x1294_x858_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89730.4]
  assign x805_lb_0_io_rPort_12_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@89729.4]
  assign x805_lb_0_io_rPort_12_ofs_0 = x942_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89731.4]
  assign x805_lb_0_io_rPort_12_en_0 = _T_1438 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89733.4]
  assign x805_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89732.4]
  assign x805_lb_0_io_rPort_11_banks_1 = x1320_x822_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90649.4]
  assign x805_lb_0_io_rPort_11_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90648.4]
  assign x805_lb_0_io_rPort_11_ofs_0 = x1028_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90650.4]
  assign x805_lb_0_io_rPort_11_en_0 = _T_1987 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90652.4]
  assign x805_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90651.4]
  assign x805_lb_0_io_rPort_10_banks_1 = x1308_x840_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@88979.4]
  assign x805_lb_0_io_rPort_10_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@88978.4]
  assign x805_lb_0_io_rPort_10_ofs_0 = x889_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@88980.4]
  assign x805_lb_0_io_rPort_10_en_0 = _T_1009 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@88982.4]
  assign x805_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@88981.4]
  assign x805_lb_0_io_rPort_9_banks_1 = x1308_x840_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89877.4]
  assign x805_lb_0_io_rPort_9_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@89876.4]
  assign x805_lb_0_io_rPort_9_ofs_0 = x957_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89878.4]
  assign x805_lb_0_io_rPort_9_en_0 = _T_1525 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89880.4]
  assign x805_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89879.4]
  assign x805_lb_0_io_rPort_8_banks_1 = x1303_x846_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89828.4]
  assign x805_lb_0_io_rPort_8_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@89827.4]
  assign x805_lb_0_io_rPort_8_ofs_0 = x952_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89829.4]
  assign x805_lb_0_io_rPort_8_en_0 = _T_1496 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89831.4]
  assign x805_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89830.4]
  assign x805_lb_0_io_rPort_7_banks_1 = x1327_x920_D5_number[3:0]; // @[MemInterfaceType.scala 106:58:@90767.4]
  assign x805_lb_0_io_rPort_7_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90766.4]
  assign x805_lb_0_io_rPort_7_ofs_0 = x1038_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90768.4]
  assign x805_lb_0_io_rPort_7_en_0 = _T_2053 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90770.4]
  assign x805_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90769.4]
  assign x805_lb_0_io_rPort_6_banks_1 = x1303_x846_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@88889.4]
  assign x805_lb_0_io_rPort_6_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@88888.4]
  assign x805_lb_0_io_rPort_6_ofs_0 = x883_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@88890.4]
  assign x805_lb_0_io_rPort_6_en_0 = _T_961 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@88892.4]
  assign x805_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@88891.4]
  assign x805_lb_0_io_rPort_5_banks_1 = x1299_x852_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89779.4]
  assign x805_lb_0_io_rPort_5_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@89778.4]
  assign x805_lb_0_io_rPort_5_ofs_0 = x947_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89780.4]
  assign x805_lb_0_io_rPort_5_en_0 = _T_1467 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89782.4]
  assign x805_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89781.4]
  assign x805_lb_0_io_rPort_4_banks_1 = x1329_x929_D5_number[3:0]; // @[MemInterfaceType.scala 106:58:@90200.4]
  assign x805_lb_0_io_rPort_4_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90199.4]
  assign x805_lb_0_io_rPort_4_ofs_0 = x987_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90201.4]
  assign x805_lb_0_io_rPort_4_en_0 = _T_1710 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90203.4]
  assign x805_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90202.4]
  assign x805_lb_0_io_rPort_3_banks_1 = x1316_x828_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@89161.4]
  assign x805_lb_0_io_rPort_3_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@89160.4]
  assign x805_lb_0_io_rPort_3_ofs_0 = x901_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@89162.4]
  assign x805_lb_0_io_rPort_3_en_0 = _T_1107 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@89164.4]
  assign x805_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@89163.4]
  assign x805_lb_0_io_rPort_2_banks_1 = x1320_x822_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90026.4]
  assign x805_lb_0_io_rPort_2_banks_0 = x1332_x1242_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90025.4]
  assign x805_lb_0_io_rPort_2_ofs_0 = x972_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90027.4]
  assign x805_lb_0_io_rPort_2_en_0 = _T_1614 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90029.4]
  assign x805_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90028.4]
  assign x805_lb_0_io_rPort_1_banks_1 = x1299_x852_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@88799.4]
  assign x805_lb_0_io_rPort_1_banks_0 = x1292_x1237_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@88798.4]
  assign x805_lb_0_io_rPort_1_ofs_0 = x877_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@88800.4]
  assign x805_lb_0_io_rPort_1_en_0 = _T_913 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@88802.4]
  assign x805_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@88801.4]
  assign x805_lb_0_io_rPort_0_banks_1 = x1316_x828_D35_number[3:0]; // @[MemInterfaceType.scala 106:58:@90600.4]
  assign x805_lb_0_io_rPort_0_banks_0 = x1348_x1247_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@90599.4]
  assign x805_lb_0_io_rPort_0_ofs_0 = x1023_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@90601.4]
  assign x805_lb_0_io_rPort_0_en_0 = _T_1958 & x1293_b802_D52; // @[MemInterfaceType.scala 110:79:@90603.4]
  assign x805_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@90602.4]
  assign x805_lb_0_io_wPort_7_banks_1 = x1281_x852_D11_number[3:0]; // @[MemInterfaceType.scala 88:58:@88393.4]
  assign x805_lb_0_io_wPort_7_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@88392.4]
  assign x805_lb_0_io_wPort_7_ofs_0 = x1283_x854_sum_D6_number[7:0]; // @[MemInterfaceType.scala 89:54:@88394.4]
  assign x805_lb_0_io_wPort_7_data_0 = RetimeWrapper_32_io_out; // @[MemInterfaceType.scala 90:56:@88395.4]
  assign x805_lb_0_io_wPort_7_en_0 = _T_691 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@88397.4]
  assign x805_lb_0_io_wPort_6_banks_1 = x1271_x828_D11_number[3:0]; // @[MemInterfaceType.scala 88:58:@87999.4]
  assign x805_lb_0_io_wPort_6_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@87998.4]
  assign x805_lb_0_io_wPort_6_ofs_0 = x1269_x830_sum_D6_number[7:0]; // @[MemInterfaceType.scala 89:54:@88000.4]
  assign x805_lb_0_io_wPort_6_data_0 = RetimeWrapper_16_io_out; // @[MemInterfaceType.scala 90:56:@88001.4]
  assign x805_lb_0_io_wPort_6_en_0 = _T_497 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@88003.4]
  assign x805_lb_0_io_wPort_5_banks_1 = x1276_x840_D11_number[3:0]; // @[MemInterfaceType.scala 88:58:@88197.4]
  assign x805_lb_0_io_wPort_5_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@88196.4]
  assign x805_lb_0_io_wPort_5_ofs_0 = x1275_x842_sum_D6_number[7:0]; // @[MemInterfaceType.scala 89:54:@88198.4]
  assign x805_lb_0_io_wPort_5_data_0 = RetimeWrapper_25_io_out; // @[MemInterfaceType.scala 90:56:@88199.4]
  assign x805_lb_0_io_wPort_5_en_0 = _T_595 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@88201.4]
  assign x805_lb_0_io_wPort_4_banks_1 = x1259_x814_D12_number[3:0]; // @[MemInterfaceType.scala 88:58:@87794.4]
  assign x805_lb_0_io_wPort_4_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@87793.4]
  assign x805_lb_0_io_wPort_4_ofs_0 = x1263_x818_sum_D7_number[7:0]; // @[MemInterfaceType.scala 89:54:@87795.4]
  assign x805_lb_0_io_wPort_4_data_0 = RetimeWrapper_6_io_out; // @[MemInterfaceType.scala 90:56:@87796.4]
  assign x805_lb_0_io_wPort_4_en_0 = _T_398 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@87798.4]
  assign x805_lb_0_io_wPort_3_banks_1 = x1272_x834_D11_number[3:0]; // @[MemInterfaceType.scala 88:58:@88099.4]
  assign x805_lb_0_io_wPort_3_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@88098.4]
  assign x805_lb_0_io_wPort_3_ofs_0 = x1273_x836_sum_D6_number[7:0]; // @[MemInterfaceType.scala 89:54:@88100.4]
  assign x805_lb_0_io_wPort_3_data_0 = RetimeWrapper_21_io_out; // @[MemInterfaceType.scala 90:56:@88101.4]
  assign x805_lb_0_io_wPort_3_en_0 = _T_547 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@88103.4]
  assign x805_lb_0_io_wPort_2_banks_1 = x1268_x822_D11_number[3:0]; // @[MemInterfaceType.scala 88:58:@87901.4]
  assign x805_lb_0_io_wPort_2_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@87900.4]
  assign x805_lb_0_io_wPort_2_ofs_0 = x1267_x824_sum_D6_number[7:0]; // @[MemInterfaceType.scala 89:54:@87902.4]
  assign x805_lb_0_io_wPort_2_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@87903.4]
  assign x805_lb_0_io_wPort_2_en_0 = _T_449 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@87905.4]
  assign x805_lb_0_io_wPort_1_banks_1 = x1278_x846_D11_number[3:0]; // @[MemInterfaceType.scala 88:58:@88295.4]
  assign x805_lb_0_io_wPort_1_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@88294.4]
  assign x805_lb_0_io_wPort_1_ofs_0 = x1279_x848_sum_D6_number[7:0]; // @[MemInterfaceType.scala 89:54:@88296.4]
  assign x805_lb_0_io_wPort_1_data_0 = RetimeWrapper_29_io_out; // @[MemInterfaceType.scala 90:56:@88297.4]
  assign x805_lb_0_io_wPort_1_en_0 = _T_643 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@88299.4]
  assign x805_lb_0_io_wPort_0_banks_1 = x1285_x858_D11_number[3:0]; // @[MemInterfaceType.scala 88:58:@88491.4]
  assign x805_lb_0_io_wPort_0_banks_0 = x1261_x1232_D26_number[2:0]; // @[MemInterfaceType.scala 88:58:@88490.4]
  assign x805_lb_0_io_wPort_0_ofs_0 = x1286_x860_sum_D6_number[7:0]; // @[MemInterfaceType.scala 89:54:@88492.4]
  assign x805_lb_0_io_wPort_0_data_0 = RetimeWrapper_35_io_out; // @[MemInterfaceType.scala 90:56:@88493.4]
  assign x805_lb_0_io_wPort_0_en_0 = _T_739 & x1260_b802_D28; // @[MemInterfaceType.scala 93:57:@88495.4]
  assign RetimeWrapper_1_clock = clock; // @[:@87632.4]
  assign RetimeWrapper_1_reset = reset; // @[:@87633.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87635.4]
  assign RetimeWrapper_1_io_in = _T_307 | _T_305; // @[package.scala 94:16:@87634.4]
  assign x814_1_clock = clock; // @[:@87654.4]
  assign x814_1_reset = reset; // @[:@87655.4]
  assign x814_1_io_a = __1_io_result; // @[Math.scala 367:17:@87656.4]
  assign x814_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@87658.4]
  assign x1235_sum_1_clock = clock; // @[:@87683.4]
  assign x1235_sum_1_reset = reset; // @[:@87684.4]
  assign x1235_sum_1_io_a = _T_347[31:0]; // @[Math.scala 151:17:@87685.4]
  assign x1235_sum_1_io_b = _T_351[31:0]; // @[Math.scala 152:17:@87686.4]
  assign x1235_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@87687.4]
  assign x817_div_1_clock = clock; // @[:@87695.4]
  assign x817_div_1_reset = reset; // @[:@87696.4]
  assign x817_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@87697.4]
  assign x817_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@87699.4]
  assign RetimeWrapper_2_clock = clock; // @[:@87705.4]
  assign RetimeWrapper_2_reset = reset; // @[:@87706.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87708.4]
  assign RetimeWrapper_2_io_in = x1235_sum_1_io_result; // @[package.scala 94:16:@87707.4]
  assign x818_sum_1_clock = clock; // @[:@87714.4]
  assign x818_sum_1_reset = reset; // @[:@87715.4]
  assign x818_sum_1_io_a = RetimeWrapper_2_io_out; // @[Math.scala 151:17:@87716.4]
  assign x818_sum_1_io_b = x817_div_1_io_result; // @[Math.scala 152:17:@87717.4]
  assign x818_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@87718.4]
  assign RetimeWrapper_3_clock = clock; // @[:@87724.4]
  assign RetimeWrapper_3_reset = reset; // @[:@87725.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87727.4]
  assign RetimeWrapper_3_io_in = x814_1_io_result; // @[package.scala 94:16:@87726.4]
  assign RetimeWrapper_4_clock = clock; // @[:@87733.4]
  assign RetimeWrapper_4_reset = reset; // @[:@87734.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87736.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@87735.4]
  assign RetimeWrapper_5_clock = clock; // @[:@87742.4]
  assign RetimeWrapper_5_reset = reset; // @[:@87743.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87745.4]
  assign RetimeWrapper_5_io_in = $unsigned(_T_325); // @[package.scala 94:16:@87744.4]
  assign RetimeWrapper_6_clock = clock; // @[:@87751.4]
  assign RetimeWrapper_6_reset = reset; // @[:@87752.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87754.4]
  assign RetimeWrapper_6_io_in = x1256_x803_D1_0_number[7:0]; // @[package.scala 94:16:@87753.4]
  assign RetimeWrapper_7_clock = clock; // @[:@87760.4]
  assign RetimeWrapper_7_reset = reset; // @[:@87761.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87763.4]
  assign RetimeWrapper_7_io_in = x818_sum_1_io_result; // @[package.scala 94:16:@87762.4]
  assign RetimeWrapper_8_clock = clock; // @[:@87769.4]
  assign RetimeWrapper_8_reset = reset; // @[:@87770.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87772.4]
  assign RetimeWrapper_8_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@87771.4]
  assign RetimeWrapper_9_clock = clock; // @[:@87780.4]
  assign RetimeWrapper_9_reset = reset; // @[:@87781.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87783.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@87782.4]
  assign x820_rdcol_1_clock = clock; // @[:@87803.4]
  assign x820_rdcol_1_reset = reset; // @[:@87804.4]
  assign x820_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@87805.4]
  assign x820_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@87806.4]
  assign x820_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@87807.4]
  assign x822_1_clock = clock; // @[:@87817.4]
  assign x822_1_reset = reset; // @[:@87818.4]
  assign x822_1_io_a = x820_rdcol_1_io_result; // @[Math.scala 367:17:@87819.4]
  assign x822_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@87821.4]
  assign x823_div_1_clock = clock; // @[:@87829.4]
  assign x823_div_1_reset = reset; // @[:@87830.4]
  assign x823_div_1_io_a = x820_rdcol_1_io_result; // @[Math.scala 328:17:@87831.4]
  assign x823_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@87833.4]
  assign RetimeWrapper_10_clock = clock; // @[:@87839.4]
  assign RetimeWrapper_10_reset = reset; // @[:@87840.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87842.4]
  assign RetimeWrapper_10_io_in = x1235_sum_1_io_result; // @[package.scala 94:16:@87841.4]
  assign x824_sum_1_clock = clock; // @[:@87848.4]
  assign x824_sum_1_reset = reset; // @[:@87849.4]
  assign x824_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@87850.4]
  assign x824_sum_1_io_b = x823_div_1_io_result; // @[Math.scala 152:17:@87851.4]
  assign x824_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@87852.4]
  assign RetimeWrapper_11_clock = clock; // @[:@87858.4]
  assign RetimeWrapper_11_reset = reset; // @[:@87859.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87861.4]
  assign RetimeWrapper_11_io_in = x1256_x803_D1_0_number[15:8]; // @[package.scala 94:16:@87860.4]
  assign RetimeWrapper_12_clock = clock; // @[:@87867.4]
  assign RetimeWrapper_12_reset = reset; // @[:@87868.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87870.4]
  assign RetimeWrapper_12_io_in = x824_sum_1_io_result; // @[package.scala 94:16:@87869.4]
  assign RetimeWrapper_13_clock = clock; // @[:@87876.4]
  assign RetimeWrapper_13_reset = reset; // @[:@87877.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87879.4]
  assign RetimeWrapper_13_io_in = x822_1_io_result; // @[package.scala 94:16:@87878.4]
  assign RetimeWrapper_14_clock = clock; // @[:@87887.4]
  assign RetimeWrapper_14_reset = reset; // @[:@87888.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87890.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@87889.4]
  assign x826_rdcol_1_clock = clock; // @[:@87910.4]
  assign x826_rdcol_1_reset = reset; // @[:@87911.4]
  assign x826_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@87912.4]
  assign x826_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@87913.4]
  assign x826_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@87914.4]
  assign x828_1_clock = clock; // @[:@87924.4]
  assign x828_1_reset = reset; // @[:@87925.4]
  assign x828_1_io_a = x826_rdcol_1_io_result; // @[Math.scala 367:17:@87926.4]
  assign x828_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@87928.4]
  assign x829_div_1_clock = clock; // @[:@87936.4]
  assign x829_div_1_reset = reset; // @[:@87937.4]
  assign x829_div_1_io_a = x826_rdcol_1_io_result; // @[Math.scala 328:17:@87938.4]
  assign x829_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@87940.4]
  assign x830_sum_1_clock = clock; // @[:@87946.4]
  assign x830_sum_1_reset = reset; // @[:@87947.4]
  assign x830_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@87948.4]
  assign x830_sum_1_io_b = x829_div_1_io_result; // @[Math.scala 152:17:@87949.4]
  assign x830_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@87950.4]
  assign RetimeWrapper_15_clock = clock; // @[:@87956.4]
  assign RetimeWrapper_15_reset = reset; // @[:@87957.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87959.4]
  assign RetimeWrapper_15_io_in = x830_sum_1_io_result; // @[package.scala 94:16:@87958.4]
  assign RetimeWrapper_16_clock = clock; // @[:@87965.4]
  assign RetimeWrapper_16_reset = reset; // @[:@87966.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87968.4]
  assign RetimeWrapper_16_io_in = x1256_x803_D1_0_number[23:16]; // @[package.scala 94:16:@87967.4]
  assign RetimeWrapper_17_clock = clock; // @[:@87974.4]
  assign RetimeWrapper_17_reset = reset; // @[:@87975.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87977.4]
  assign RetimeWrapper_17_io_in = x828_1_io_result; // @[package.scala 94:16:@87976.4]
  assign RetimeWrapper_18_clock = clock; // @[:@87985.4]
  assign RetimeWrapper_18_reset = reset; // @[:@87986.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@87988.4]
  assign RetimeWrapper_18_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@87987.4]
  assign x832_rdcol_1_clock = clock; // @[:@88008.4]
  assign x832_rdcol_1_reset = reset; // @[:@88009.4]
  assign x832_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@88010.4]
  assign x832_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@88011.4]
  assign x832_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88012.4]
  assign x834_1_clock = clock; // @[:@88024.4]
  assign x834_1_reset = reset; // @[:@88025.4]
  assign x834_1_io_a = x832_rdcol_1_io_result; // @[Math.scala 367:17:@88026.4]
  assign x834_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@88028.4]
  assign x835_div_1_clock = clock; // @[:@88036.4]
  assign x835_div_1_reset = reset; // @[:@88037.4]
  assign x835_div_1_io_a = x832_rdcol_1_io_result; // @[Math.scala 328:17:@88038.4]
  assign x835_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@88040.4]
  assign x836_sum_1_clock = clock; // @[:@88046.4]
  assign x836_sum_1_reset = reset; // @[:@88047.4]
  assign x836_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@88048.4]
  assign x836_sum_1_io_b = x835_div_1_io_result; // @[Math.scala 152:17:@88049.4]
  assign x836_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88050.4]
  assign RetimeWrapper_19_clock = clock; // @[:@88056.4]
  assign RetimeWrapper_19_reset = reset; // @[:@88057.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88059.4]
  assign RetimeWrapper_19_io_in = x834_1_io_result; // @[package.scala 94:16:@88058.4]
  assign RetimeWrapper_20_clock = clock; // @[:@88065.4]
  assign RetimeWrapper_20_reset = reset; // @[:@88066.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88068.4]
  assign RetimeWrapper_20_io_in = x836_sum_1_io_result; // @[package.scala 94:16:@88067.4]
  assign RetimeWrapper_21_clock = clock; // @[:@88074.4]
  assign RetimeWrapper_21_reset = reset; // @[:@88075.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88077.4]
  assign RetimeWrapper_21_io_in = x1256_x803_D1_0_number[31:24]; // @[package.scala 94:16:@88076.4]
  assign RetimeWrapper_22_clock = clock; // @[:@88085.4]
  assign RetimeWrapper_22_reset = reset; // @[:@88086.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88088.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88087.4]
  assign x838_rdcol_1_clock = clock; // @[:@88108.4]
  assign x838_rdcol_1_reset = reset; // @[:@88109.4]
  assign x838_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@88110.4]
  assign x838_rdcol_1_io_b = 32'h4; // @[Math.scala 152:17:@88111.4]
  assign x838_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88112.4]
  assign x840_1_clock = clock; // @[:@88122.4]
  assign x840_1_reset = reset; // @[:@88123.4]
  assign x840_1_io_a = x838_rdcol_1_io_result; // @[Math.scala 367:17:@88124.4]
  assign x840_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@88126.4]
  assign x841_div_1_clock = clock; // @[:@88134.4]
  assign x841_div_1_reset = reset; // @[:@88135.4]
  assign x841_div_1_io_a = x838_rdcol_1_io_result; // @[Math.scala 328:17:@88136.4]
  assign x841_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@88138.4]
  assign x842_sum_1_clock = clock; // @[:@88144.4]
  assign x842_sum_1_reset = reset; // @[:@88145.4]
  assign x842_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@88146.4]
  assign x842_sum_1_io_b = x841_div_1_io_result; // @[Math.scala 152:17:@88147.4]
  assign x842_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88148.4]
  assign RetimeWrapper_23_clock = clock; // @[:@88154.4]
  assign RetimeWrapper_23_reset = reset; // @[:@88155.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88157.4]
  assign RetimeWrapper_23_io_in = x842_sum_1_io_result; // @[package.scala 94:16:@88156.4]
  assign RetimeWrapper_24_clock = clock; // @[:@88163.4]
  assign RetimeWrapper_24_reset = reset; // @[:@88164.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88166.4]
  assign RetimeWrapper_24_io_in = x840_1_io_result; // @[package.scala 94:16:@88165.4]
  assign RetimeWrapper_25_clock = clock; // @[:@88172.4]
  assign RetimeWrapper_25_reset = reset; // @[:@88173.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88175.4]
  assign RetimeWrapper_25_io_in = x1256_x803_D1_0_number[39:32]; // @[package.scala 94:16:@88174.4]
  assign RetimeWrapper_26_clock = clock; // @[:@88183.4]
  assign RetimeWrapper_26_reset = reset; // @[:@88184.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88186.4]
  assign RetimeWrapper_26_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88185.4]
  assign x844_rdcol_1_clock = clock; // @[:@88206.4]
  assign x844_rdcol_1_reset = reset; // @[:@88207.4]
  assign x844_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@88208.4]
  assign x844_rdcol_1_io_b = 32'h5; // @[Math.scala 152:17:@88209.4]
  assign x844_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88210.4]
  assign x846_1_clock = clock; // @[:@88220.4]
  assign x846_1_reset = reset; // @[:@88221.4]
  assign x846_1_io_a = x844_rdcol_1_io_result; // @[Math.scala 367:17:@88222.4]
  assign x846_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@88224.4]
  assign x847_div_1_clock = clock; // @[:@88232.4]
  assign x847_div_1_reset = reset; // @[:@88233.4]
  assign x847_div_1_io_a = x844_rdcol_1_io_result; // @[Math.scala 328:17:@88234.4]
  assign x847_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@88236.4]
  assign x848_sum_1_clock = clock; // @[:@88242.4]
  assign x848_sum_1_reset = reset; // @[:@88243.4]
  assign x848_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@88244.4]
  assign x848_sum_1_io_b = x847_div_1_io_result; // @[Math.scala 152:17:@88245.4]
  assign x848_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88246.4]
  assign RetimeWrapper_27_clock = clock; // @[:@88252.4]
  assign RetimeWrapper_27_reset = reset; // @[:@88253.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88255.4]
  assign RetimeWrapper_27_io_in = x846_1_io_result; // @[package.scala 94:16:@88254.4]
  assign RetimeWrapper_28_clock = clock; // @[:@88261.4]
  assign RetimeWrapper_28_reset = reset; // @[:@88262.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88264.4]
  assign RetimeWrapper_28_io_in = x848_sum_1_io_result; // @[package.scala 94:16:@88263.4]
  assign RetimeWrapper_29_clock = clock; // @[:@88270.4]
  assign RetimeWrapper_29_reset = reset; // @[:@88271.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88273.4]
  assign RetimeWrapper_29_io_in = x1256_x803_D1_0_number[47:40]; // @[package.scala 94:16:@88272.4]
  assign RetimeWrapper_30_clock = clock; // @[:@88281.4]
  assign RetimeWrapper_30_reset = reset; // @[:@88282.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88284.4]
  assign RetimeWrapper_30_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88283.4]
  assign x850_rdcol_1_clock = clock; // @[:@88304.4]
  assign x850_rdcol_1_reset = reset; // @[:@88305.4]
  assign x850_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@88306.4]
  assign x850_rdcol_1_io_b = 32'h6; // @[Math.scala 152:17:@88307.4]
  assign x850_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88308.4]
  assign x852_1_clock = clock; // @[:@88318.4]
  assign x852_1_reset = reset; // @[:@88319.4]
  assign x852_1_io_a = x850_rdcol_1_io_result; // @[Math.scala 367:17:@88320.4]
  assign x852_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@88322.4]
  assign x853_div_1_clock = clock; // @[:@88330.4]
  assign x853_div_1_reset = reset; // @[:@88331.4]
  assign x853_div_1_io_a = x850_rdcol_1_io_result; // @[Math.scala 328:17:@88332.4]
  assign x853_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@88334.4]
  assign x854_sum_1_clock = clock; // @[:@88340.4]
  assign x854_sum_1_reset = reset; // @[:@88341.4]
  assign x854_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@88342.4]
  assign x854_sum_1_io_b = x853_div_1_io_result; // @[Math.scala 152:17:@88343.4]
  assign x854_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88344.4]
  assign RetimeWrapper_31_clock = clock; // @[:@88350.4]
  assign RetimeWrapper_31_reset = reset; // @[:@88351.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88353.4]
  assign RetimeWrapper_31_io_in = x852_1_io_result; // @[package.scala 94:16:@88352.4]
  assign RetimeWrapper_32_clock = clock; // @[:@88359.4]
  assign RetimeWrapper_32_reset = reset; // @[:@88360.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88362.4]
  assign RetimeWrapper_32_io_in = x1256_x803_D1_0_number[55:48]; // @[package.scala 94:16:@88361.4]
  assign RetimeWrapper_33_clock = clock; // @[:@88368.4]
  assign RetimeWrapper_33_reset = reset; // @[:@88369.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88371.4]
  assign RetimeWrapper_33_io_in = x854_sum_1_io_result; // @[package.scala 94:16:@88370.4]
  assign RetimeWrapper_34_clock = clock; // @[:@88379.4]
  assign RetimeWrapper_34_reset = reset; // @[:@88380.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88382.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88381.4]
  assign x856_rdcol_1_clock = clock; // @[:@88402.4]
  assign x856_rdcol_1_reset = reset; // @[:@88403.4]
  assign x856_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@88404.4]
  assign x856_rdcol_1_io_b = 32'h7; // @[Math.scala 152:17:@88405.4]
  assign x856_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88406.4]
  assign x858_1_clock = clock; // @[:@88416.4]
  assign x858_1_reset = reset; // @[:@88417.4]
  assign x858_1_io_a = x856_rdcol_1_io_result; // @[Math.scala 367:17:@88418.4]
  assign x858_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@88420.4]
  assign x859_div_1_clock = clock; // @[:@88428.4]
  assign x859_div_1_reset = reset; // @[:@88429.4]
  assign x859_div_1_io_a = x856_rdcol_1_io_result; // @[Math.scala 328:17:@88430.4]
  assign x859_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@88432.4]
  assign x860_sum_1_clock = clock; // @[:@88438.4]
  assign x860_sum_1_reset = reset; // @[:@88439.4]
  assign x860_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@88440.4]
  assign x860_sum_1_io_b = x859_div_1_io_result; // @[Math.scala 152:17:@88441.4]
  assign x860_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88442.4]
  assign RetimeWrapper_35_clock = clock; // @[:@88448.4]
  assign RetimeWrapper_35_reset = reset; // @[:@88449.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88451.4]
  assign RetimeWrapper_35_io_in = x1256_x803_D1_0_number[63:56]; // @[package.scala 94:16:@88450.4]
  assign RetimeWrapper_36_clock = clock; // @[:@88457.4]
  assign RetimeWrapper_36_reset = reset; // @[:@88458.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88460.4]
  assign RetimeWrapper_36_io_in = x858_1_io_result; // @[package.scala 94:16:@88459.4]
  assign RetimeWrapper_37_clock = clock; // @[:@88466.4]
  assign RetimeWrapper_37_reset = reset; // @[:@88467.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88469.4]
  assign RetimeWrapper_37_io_in = x860_sum_1_io_result; // @[package.scala 94:16:@88468.4]
  assign RetimeWrapper_38_clock = clock; // @[:@88477.4]
  assign RetimeWrapper_38_reset = reset; // @[:@88478.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88480.4]
  assign RetimeWrapper_38_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88479.4]
  assign RetimeWrapper_39_clock = clock; // @[:@88498.4]
  assign RetimeWrapper_39_reset = reset; // @[:@88499.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88501.4]
  assign RetimeWrapper_39_io_in = __io_result; // @[package.scala 94:16:@88500.4]
  assign RetimeWrapper_40_clock = clock; // @[:@88514.4]
  assign RetimeWrapper_40_reset = reset; // @[:@88515.4]
  assign RetimeWrapper_40_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@88518.4]
  assign RetimeWrapper_40_io_in = $unsigned(_T_754); // @[package.scala 94:16:@88517.4]
  assign RetimeWrapper_41_clock = clock; // @[:@88532.4]
  assign RetimeWrapper_41_reset = reset; // @[:@88533.4]
  assign RetimeWrapper_41_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@88535.4]
  assign RetimeWrapper_41_io_in = $signed(_T_751) < $signed(32'sh0); // @[package.scala 94:16:@88534.4]
  assign RetimeWrapper_42_clock = clock; // @[:@88541.4]
  assign RetimeWrapper_42_reset = reset; // @[:@88542.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88544.4]
  assign RetimeWrapper_42_io_in = x856_rdcol_1_io_result; // @[package.scala 94:16:@88543.4]
  assign RetimeWrapper_43_clock = clock; // @[:@88555.4]
  assign RetimeWrapper_43_reset = reset; // @[:@88556.4]
  assign RetimeWrapper_43_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@88558.4]
  assign RetimeWrapper_43_io_in = $signed(_T_778) < $signed(32'sh0); // @[package.scala 94:16:@88557.4]
  assign RetimeWrapper_44_clock = clock; // @[:@88564.4]
  assign RetimeWrapper_44_reset = reset; // @[:@88565.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88567.4]
  assign RetimeWrapper_44_io_in = RetimeWrapper_41_io_out; // @[package.scala 94:16:@88566.4]
  assign x1240_sum_1_clock = clock; // @[:@88611.4]
  assign x1240_sum_1_reset = reset; // @[:@88612.4]
  assign x1240_sum_1_io_a = _T_817[31:0]; // @[Math.scala 151:17:@88613.4]
  assign x1240_sum_1_io_b = _T_821[31:0]; // @[Math.scala 152:17:@88614.4]
  assign x1240_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88615.4]
  assign RetimeWrapper_45_clock = clock; // @[:@88621.4]
  assign RetimeWrapper_45_reset = reset; // @[:@88622.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88624.4]
  assign RetimeWrapper_45_io_in = x1240_sum_1_io_result; // @[package.scala 94:16:@88623.4]
  assign RetimeWrapper_46_clock = clock; // @[:@88630.4]
  assign RetimeWrapper_46_reset = reset; // @[:@88631.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88633.4]
  assign RetimeWrapper_46_io_in = x859_div_1_io_result; // @[package.scala 94:16:@88632.4]
  assign x871_sum_1_clock = clock; // @[:@88639.4]
  assign x871_sum_1_reset = reset; // @[:@88640.4]
  assign x871_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@88641.4]
  assign x871_sum_1_io_b = RetimeWrapper_46_io_out; // @[Math.scala 152:17:@88642.4]
  assign x871_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88643.4]
  assign RetimeWrapper_47_clock = clock; // @[:@88649.4]
  assign RetimeWrapper_47_reset = reset; // @[:@88650.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88652.4]
  assign RetimeWrapper_47_io_in = $unsigned(_T_802); // @[package.scala 94:16:@88651.4]
  assign RetimeWrapper_48_clock = clock; // @[:@88658.4]
  assign RetimeWrapper_48_reset = reset; // @[:@88659.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88661.4]
  assign RetimeWrapper_48_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@88660.4]
  assign RetimeWrapper_49_clock = clock; // @[:@88667.4]
  assign RetimeWrapper_49_reset = reset; // @[:@88668.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88670.4]
  assign RetimeWrapper_49_io_in = x858_1_io_result; // @[package.scala 94:16:@88669.4]
  assign RetimeWrapper_50_clock = clock; // @[:@88676.4]
  assign RetimeWrapper_50_reset = reset; // @[:@88677.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88679.4]
  assign RetimeWrapper_50_io_in = ~ x866; // @[package.scala 94:16:@88678.4]
  assign RetimeWrapper_51_clock = clock; // @[:@88685.4]
  assign RetimeWrapper_51_reset = reset; // @[:@88686.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88688.4]
  assign RetimeWrapper_51_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@88687.4]
  assign RetimeWrapper_52_clock = clock; // @[:@88697.4]
  assign RetimeWrapper_52_reset = reset; // @[:@88698.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88700.4]
  assign RetimeWrapper_52_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88699.4]
  assign RetimeWrapper_53_clock = clock; // @[:@88718.4]
  assign RetimeWrapper_53_reset = reset; // @[:@88719.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88721.4]
  assign RetimeWrapper_53_io_in = x850_rdcol_1_io_result; // @[package.scala 94:16:@88720.4]
  assign RetimeWrapper_54_clock = clock; // @[:@88732.4]
  assign RetimeWrapper_54_reset = reset; // @[:@88733.4]
  assign RetimeWrapper_54_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@88735.4]
  assign RetimeWrapper_54_io_in = $signed(_T_876) < $signed(32'sh0); // @[package.scala 94:16:@88734.4]
  assign RetimeWrapper_55_clock = clock; // @[:@88747.4]
  assign RetimeWrapper_55_reset = reset; // @[:@88748.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88750.4]
  assign RetimeWrapper_55_io_in = x853_div_1_io_result; // @[package.scala 94:16:@88749.4]
  assign x877_sum_1_clock = clock; // @[:@88756.4]
  assign x877_sum_1_reset = reset; // @[:@88757.4]
  assign x877_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@88758.4]
  assign x877_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@88759.4]
  assign x877_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88760.4]
  assign RetimeWrapper_56_clock = clock; // @[:@88766.4]
  assign RetimeWrapper_56_reset = reset; // @[:@88767.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88769.4]
  assign RetimeWrapper_56_io_in = x852_1_io_result; // @[package.scala 94:16:@88768.4]
  assign RetimeWrapper_57_clock = clock; // @[:@88775.4]
  assign RetimeWrapper_57_reset = reset; // @[:@88776.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88778.4]
  assign RetimeWrapper_57_io_in = ~ x875; // @[package.scala 94:16:@88777.4]
  assign RetimeWrapper_58_clock = clock; // @[:@88787.4]
  assign RetimeWrapper_58_reset = reset; // @[:@88788.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88790.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88789.4]
  assign RetimeWrapper_59_clock = clock; // @[:@88808.4]
  assign RetimeWrapper_59_reset = reset; // @[:@88809.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88811.4]
  assign RetimeWrapper_59_io_in = x844_rdcol_1_io_result; // @[package.scala 94:16:@88810.4]
  assign RetimeWrapper_60_clock = clock; // @[:@88822.4]
  assign RetimeWrapper_60_reset = reset; // @[:@88823.4]
  assign RetimeWrapper_60_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@88825.4]
  assign RetimeWrapper_60_io_in = $signed(_T_924) < $signed(32'sh0); // @[package.scala 94:16:@88824.4]
  assign RetimeWrapper_61_clock = clock; // @[:@88837.4]
  assign RetimeWrapper_61_reset = reset; // @[:@88838.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88840.4]
  assign RetimeWrapper_61_io_in = x847_div_1_io_result; // @[package.scala 94:16:@88839.4]
  assign x883_sum_1_clock = clock; // @[:@88846.4]
  assign x883_sum_1_reset = reset; // @[:@88847.4]
  assign x883_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@88848.4]
  assign x883_sum_1_io_b = RetimeWrapper_61_io_out; // @[Math.scala 152:17:@88849.4]
  assign x883_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88850.4]
  assign RetimeWrapper_62_clock = clock; // @[:@88856.4]
  assign RetimeWrapper_62_reset = reset; // @[:@88857.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88859.4]
  assign RetimeWrapper_62_io_in = x846_1_io_result; // @[package.scala 94:16:@88858.4]
  assign RetimeWrapper_63_clock = clock; // @[:@88865.4]
  assign RetimeWrapper_63_reset = reset; // @[:@88866.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88868.4]
  assign RetimeWrapper_63_io_in = ~ x881; // @[package.scala 94:16:@88867.4]
  assign RetimeWrapper_64_clock = clock; // @[:@88877.4]
  assign RetimeWrapper_64_reset = reset; // @[:@88878.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88880.4]
  assign RetimeWrapper_64_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88879.4]
  assign RetimeWrapper_65_clock = clock; // @[:@88898.4]
  assign RetimeWrapper_65_reset = reset; // @[:@88899.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88901.4]
  assign RetimeWrapper_65_io_in = x838_rdcol_1_io_result; // @[package.scala 94:16:@88900.4]
  assign RetimeWrapper_66_clock = clock; // @[:@88912.4]
  assign RetimeWrapper_66_reset = reset; // @[:@88913.4]
  assign RetimeWrapper_66_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@88915.4]
  assign RetimeWrapper_66_io_in = $signed(_T_972) < $signed(32'sh0); // @[package.scala 94:16:@88914.4]
  assign RetimeWrapper_67_clock = clock; // @[:@88927.4]
  assign RetimeWrapper_67_reset = reset; // @[:@88928.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88930.4]
  assign RetimeWrapper_67_io_in = x841_div_1_io_result; // @[package.scala 94:16:@88929.4]
  assign x889_sum_1_clock = clock; // @[:@88936.4]
  assign x889_sum_1_reset = reset; // @[:@88937.4]
  assign x889_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@88938.4]
  assign x889_sum_1_io_b = RetimeWrapper_67_io_out; // @[Math.scala 152:17:@88939.4]
  assign x889_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@88940.4]
  assign RetimeWrapper_68_clock = clock; // @[:@88946.4]
  assign RetimeWrapper_68_reset = reset; // @[:@88947.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88949.4]
  assign RetimeWrapper_68_io_in = ~ x887; // @[package.scala 94:16:@88948.4]
  assign RetimeWrapper_69_clock = clock; // @[:@88955.4]
  assign RetimeWrapper_69_reset = reset; // @[:@88956.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88958.4]
  assign RetimeWrapper_69_io_in = x840_1_io_result; // @[package.scala 94:16:@88957.4]
  assign RetimeWrapper_70_clock = clock; // @[:@88967.4]
  assign RetimeWrapper_70_reset = reset; // @[:@88968.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88970.4]
  assign RetimeWrapper_70_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@88969.4]
  assign RetimeWrapper_71_clock = clock; // @[:@88988.4]
  assign RetimeWrapper_71_reset = reset; // @[:@88989.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@88991.4]
  assign RetimeWrapper_71_io_in = x832_rdcol_1_io_result; // @[package.scala 94:16:@88990.4]
  assign RetimeWrapper_72_clock = clock; // @[:@89004.4]
  assign RetimeWrapper_72_reset = reset; // @[:@89005.4]
  assign RetimeWrapper_72_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89007.4]
  assign RetimeWrapper_72_io_in = $signed(_T_1022) < $signed(32'sh0); // @[package.scala 94:16:@89006.4]
  assign RetimeWrapper_73_clock = clock; // @[:@89019.4]
  assign RetimeWrapper_73_reset = reset; // @[:@89020.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89022.4]
  assign RetimeWrapper_73_io_in = x835_div_1_io_result; // @[package.scala 94:16:@89021.4]
  assign x895_sum_1_clock = clock; // @[:@89028.4]
  assign x895_sum_1_reset = reset; // @[:@89029.4]
  assign x895_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@89030.4]
  assign x895_sum_1_io_b = RetimeWrapper_73_io_out; // @[Math.scala 152:17:@89031.4]
  assign x895_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89032.4]
  assign RetimeWrapper_74_clock = clock; // @[:@89038.4]
  assign RetimeWrapper_74_reset = reset; // @[:@89039.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89041.4]
  assign RetimeWrapper_74_io_in = x834_1_io_result; // @[package.scala 94:16:@89040.4]
  assign RetimeWrapper_75_clock = clock; // @[:@89047.4]
  assign RetimeWrapper_75_reset = reset; // @[:@89048.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89050.4]
  assign RetimeWrapper_75_io_in = ~ x893; // @[package.scala 94:16:@89049.4]
  assign RetimeWrapper_76_clock = clock; // @[:@89059.4]
  assign RetimeWrapper_76_reset = reset; // @[:@89060.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89062.4]
  assign RetimeWrapper_76_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89061.4]
  assign RetimeWrapper_77_clock = clock; // @[:@89080.4]
  assign RetimeWrapper_77_reset = reset; // @[:@89081.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89083.4]
  assign RetimeWrapper_77_io_in = x826_rdcol_1_io_result; // @[package.scala 94:16:@89082.4]
  assign RetimeWrapper_78_clock = clock; // @[:@89094.4]
  assign RetimeWrapper_78_reset = reset; // @[:@89095.4]
  assign RetimeWrapper_78_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89097.4]
  assign RetimeWrapper_78_io_in = $signed(_T_1070) < $signed(32'sh0); // @[package.scala 94:16:@89096.4]
  assign RetimeWrapper_79_clock = clock; // @[:@89109.4]
  assign RetimeWrapper_79_reset = reset; // @[:@89110.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89112.4]
  assign RetimeWrapper_79_io_in = x829_div_1_io_result; // @[package.scala 94:16:@89111.4]
  assign x901_sum_1_clock = clock; // @[:@89118.4]
  assign x901_sum_1_reset = reset; // @[:@89119.4]
  assign x901_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@89120.4]
  assign x901_sum_1_io_b = RetimeWrapper_79_io_out; // @[Math.scala 152:17:@89121.4]
  assign x901_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89122.4]
  assign RetimeWrapper_80_clock = clock; // @[:@89128.4]
  assign RetimeWrapper_80_reset = reset; // @[:@89129.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89131.4]
  assign RetimeWrapper_80_io_in = ~ x899; // @[package.scala 94:16:@89130.4]
  assign RetimeWrapper_81_clock = clock; // @[:@89137.4]
  assign RetimeWrapper_81_reset = reset; // @[:@89138.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89140.4]
  assign RetimeWrapper_81_io_in = x828_1_io_result; // @[package.scala 94:16:@89139.4]
  assign RetimeWrapper_82_clock = clock; // @[:@89149.4]
  assign RetimeWrapper_82_reset = reset; // @[:@89150.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89152.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89151.4]
  assign RetimeWrapper_83_clock = clock; // @[:@89170.4]
  assign RetimeWrapper_83_reset = reset; // @[:@89171.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89173.4]
  assign RetimeWrapper_83_io_in = x820_rdcol_1_io_result; // @[package.scala 94:16:@89172.4]
  assign RetimeWrapper_84_clock = clock; // @[:@89184.4]
  assign RetimeWrapper_84_reset = reset; // @[:@89185.4]
  assign RetimeWrapper_84_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89187.4]
  assign RetimeWrapper_84_io_in = $signed(_T_1118) < $signed(32'sh0); // @[package.scala 94:16:@89186.4]
  assign RetimeWrapper_85_clock = clock; // @[:@89199.4]
  assign RetimeWrapper_85_reset = reset; // @[:@89200.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89202.4]
  assign RetimeWrapper_85_io_in = x823_div_1_io_result; // @[package.scala 94:16:@89201.4]
  assign x907_sum_1_clock = clock; // @[:@89208.4]
  assign x907_sum_1_reset = reset; // @[:@89209.4]
  assign x907_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@89210.4]
  assign x907_sum_1_io_b = RetimeWrapper_85_io_out; // @[Math.scala 152:17:@89211.4]
  assign x907_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89212.4]
  assign RetimeWrapper_86_clock = clock; // @[:@89218.4]
  assign RetimeWrapper_86_reset = reset; // @[:@89219.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89221.4]
  assign RetimeWrapper_86_io_in = ~ x905; // @[package.scala 94:16:@89220.4]
  assign RetimeWrapper_87_clock = clock; // @[:@89227.4]
  assign RetimeWrapper_87_reset = reset; // @[:@89228.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89230.4]
  assign RetimeWrapper_87_io_in = x822_1_io_result; // @[package.scala 94:16:@89229.4]
  assign RetimeWrapper_88_clock = clock; // @[:@89239.4]
  assign RetimeWrapper_88_reset = reset; // @[:@89240.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89242.4]
  assign RetimeWrapper_88_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89241.4]
  assign RetimeWrapper_89_clock = clock; // @[:@89260.4]
  assign RetimeWrapper_89_reset = reset; // @[:@89261.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89263.4]
  assign RetimeWrapper_89_io_in = __1_io_result; // @[package.scala 94:16:@89262.4]
  assign RetimeWrapper_90_clock = clock; // @[:@89274.4]
  assign RetimeWrapper_90_reset = reset; // @[:@89275.4]
  assign RetimeWrapper_90_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89277.4]
  assign RetimeWrapper_90_io_in = $signed(_T_1166) < $signed(32'sh0); // @[package.scala 94:16:@89276.4]
  assign RetimeWrapper_91_clock = clock; // @[:@89289.4]
  assign RetimeWrapper_91_reset = reset; // @[:@89290.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89292.4]
  assign RetimeWrapper_91_io_in = x1240_sum_1_io_result; // @[package.scala 94:16:@89291.4]
  assign RetimeWrapper_92_clock = clock; // @[:@89298.4]
  assign RetimeWrapper_92_reset = reset; // @[:@89299.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89301.4]
  assign RetimeWrapper_92_io_in = x817_div_1_io_result; // @[package.scala 94:16:@89300.4]
  assign x913_sum_1_clock = clock; // @[:@89307.4]
  assign x913_sum_1_reset = reset; // @[:@89308.4]
  assign x913_sum_1_io_a = RetimeWrapper_91_io_out; // @[Math.scala 151:17:@89309.4]
  assign x913_sum_1_io_b = RetimeWrapper_92_io_out; // @[Math.scala 152:17:@89310.4]
  assign x913_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89311.4]
  assign RetimeWrapper_93_clock = clock; // @[:@89317.4]
  assign RetimeWrapper_93_reset = reset; // @[:@89318.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89320.4]
  assign RetimeWrapper_93_io_in = x814_1_io_result; // @[package.scala 94:16:@89319.4]
  assign RetimeWrapper_94_clock = clock; // @[:@89326.4]
  assign RetimeWrapper_94_reset = reset; // @[:@89327.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89329.4]
  assign RetimeWrapper_94_io_in = x913_sum_1_io_result; // @[package.scala 94:16:@89328.4]
  assign RetimeWrapper_95_clock = clock; // @[:@89335.4]
  assign RetimeWrapper_95_reset = reset; // @[:@89336.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89338.4]
  assign RetimeWrapper_95_io_in = ~ x911; // @[package.scala 94:16:@89337.4]
  assign RetimeWrapper_96_clock = clock; // @[:@89347.4]
  assign RetimeWrapper_96_reset = reset; // @[:@89348.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89350.4]
  assign RetimeWrapper_96_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89349.4]
  assign x916_rdcol_1_clock = clock; // @[:@89370.4]
  assign x916_rdcol_1_reset = reset; // @[:@89371.4]
  assign x916_rdcol_1_io_a = RetimeWrapper_89_io_out; // @[Math.scala 151:17:@89372.4]
  assign x916_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@89373.4]
  assign x916_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89374.4]
  assign RetimeWrapper_97_clock = clock; // @[:@89385.4]
  assign RetimeWrapper_97_reset = reset; // @[:@89386.4]
  assign RetimeWrapper_97_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89388.4]
  assign RetimeWrapper_97_io_in = $signed(_T_1224) < $signed(32'sh0); // @[package.scala 94:16:@89387.4]
  assign x920_1_clock = clock; // @[:@89402.4]
  assign x920_1_reset = reset; // @[:@89403.4]
  assign x920_1_io_a = x916_rdcol_1_io_result; // @[Math.scala 367:17:@89404.4]
  assign x920_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@89406.4]
  assign x921_div_1_clock = clock; // @[:@89414.4]
  assign x921_div_1_reset = reset; // @[:@89415.4]
  assign x921_div_1_io_a = x916_rdcol_1_io_result; // @[Math.scala 328:17:@89416.4]
  assign x921_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@89418.4]
  assign x922_sum_1_clock = clock; // @[:@89424.4]
  assign x922_sum_1_reset = reset; // @[:@89425.4]
  assign x922_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@89426.4]
  assign x922_sum_1_io_b = x921_div_1_io_result; // @[Math.scala 152:17:@89427.4]
  assign x922_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89428.4]
  assign RetimeWrapper_98_clock = clock; // @[:@89434.4]
  assign RetimeWrapper_98_reset = reset; // @[:@89435.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89437.4]
  assign RetimeWrapper_98_io_in = x920_1_io_result; // @[package.scala 94:16:@89436.4]
  assign RetimeWrapper_99_clock = clock; // @[:@89443.4]
  assign RetimeWrapper_99_reset = reset; // @[:@89444.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89446.4]
  assign RetimeWrapper_99_io_in = ~ x918; // @[package.scala 94:16:@89445.4]
  assign RetimeWrapper_100_clock = clock; // @[:@89455.4]
  assign RetimeWrapper_100_reset = reset; // @[:@89456.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89458.4]
  assign RetimeWrapper_100_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89457.4]
  assign x925_rdcol_1_clock = clock; // @[:@89480.4]
  assign x925_rdcol_1_reset = reset; // @[:@89481.4]
  assign x925_rdcol_1_io_a = RetimeWrapper_89_io_out; // @[Math.scala 151:17:@89482.4]
  assign x925_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@89483.4]
  assign x925_rdcol_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89484.4]
  assign RetimeWrapper_101_clock = clock; // @[:@89495.4]
  assign RetimeWrapper_101_reset = reset; // @[:@89496.4]
  assign RetimeWrapper_101_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89498.4]
  assign RetimeWrapper_101_io_in = $signed(_T_1289) < $signed(32'sh0); // @[package.scala 94:16:@89497.4]
  assign x929_1_clock = clock; // @[:@89512.4]
  assign x929_1_reset = reset; // @[:@89513.4]
  assign x929_1_io_a = x925_rdcol_1_io_result; // @[Math.scala 367:17:@89514.4]
  assign x929_1_io_flow = io_in_x745_TREADY; // @[Math.scala 369:20:@89516.4]
  assign x930_div_1_clock = clock; // @[:@89524.4]
  assign x930_div_1_reset = reset; // @[:@89525.4]
  assign x930_div_1_io_a = x925_rdcol_1_io_result; // @[Math.scala 328:17:@89526.4]
  assign x930_div_1_io_flow = io_in_x745_TREADY; // @[Math.scala 330:20:@89528.4]
  assign x931_sum_1_clock = clock; // @[:@89534.4]
  assign x931_sum_1_reset = reset; // @[:@89535.4]
  assign x931_sum_1_io_a = RetimeWrapper_45_io_out; // @[Math.scala 151:17:@89536.4]
  assign x931_sum_1_io_b = x930_div_1_io_result; // @[Math.scala 152:17:@89537.4]
  assign x931_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89538.4]
  assign RetimeWrapper_102_clock = clock; // @[:@89544.4]
  assign RetimeWrapper_102_reset = reset; // @[:@89545.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89547.4]
  assign RetimeWrapper_102_io_in = x929_1_io_result; // @[package.scala 94:16:@89546.4]
  assign RetimeWrapper_103_clock = clock; // @[:@89553.4]
  assign RetimeWrapper_103_reset = reset; // @[:@89554.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89556.4]
  assign RetimeWrapper_103_io_in = ~ x927; // @[package.scala 94:16:@89555.4]
  assign RetimeWrapper_104_clock = clock; // @[:@89565.4]
  assign RetimeWrapper_104_reset = reset; // @[:@89566.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89568.4]
  assign RetimeWrapper_104_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89567.4]
  assign x934_rdrow_1_clock = clock; // @[:@89588.4]
  assign x934_rdrow_1_reset = reset; // @[:@89589.4]
  assign x934_rdrow_1_io_a = RetimeWrapper_39_io_out; // @[Math.scala 192:17:@89590.4]
  assign x934_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@89591.4]
  assign x934_rdrow_1_io_flow = io_in_x745_TREADY; // @[Math.scala 194:20:@89592.4]
  assign RetimeWrapper_105_clock = clock; // @[:@89605.4]
  assign RetimeWrapper_105_reset = reset; // @[:@89606.4]
  assign RetimeWrapper_105_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89609.4]
  assign RetimeWrapper_105_io_in = $unsigned(_T_1357); // @[package.scala 94:16:@89608.4]
  assign RetimeWrapper_106_clock = clock; // @[:@89623.4]
  assign RetimeWrapper_106_reset = reset; // @[:@89624.4]
  assign RetimeWrapper_106_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@89626.4]
  assign RetimeWrapper_106_io_in = $signed(_T_1354) < $signed(32'sh0); // @[package.scala 94:16:@89625.4]
  assign x1245_sum_1_clock = clock; // @[:@89668.4]
  assign x1245_sum_1_reset = reset; // @[:@89669.4]
  assign x1245_sum_1_io_a = _T_1402[31:0]; // @[Math.scala 151:17:@89670.4]
  assign x1245_sum_1_io_b = _T_1406[31:0]; // @[Math.scala 152:17:@89671.4]
  assign x1245_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89672.4]
  assign RetimeWrapper_107_clock = clock; // @[:@89678.4]
  assign RetimeWrapper_107_reset = reset; // @[:@89679.4]
  assign RetimeWrapper_107_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89681.4]
  assign RetimeWrapper_107_io_in = x1245_sum_1_io_result; // @[package.scala 94:16:@89680.4]
  assign x942_sum_1_clock = clock; // @[:@89687.4]
  assign x942_sum_1_reset = reset; // @[:@89688.4]
  assign x942_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@89689.4]
  assign x942_sum_1_io_b = RetimeWrapper_46_io_out; // @[Math.scala 152:17:@89690.4]
  assign x942_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89691.4]
  assign RetimeWrapper_108_clock = clock; // @[:@89697.4]
  assign RetimeWrapper_108_reset = reset; // @[:@89698.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89700.4]
  assign RetimeWrapper_108_io_in = $unsigned(_T_1387); // @[package.scala 94:16:@89699.4]
  assign RetimeWrapper_109_clock = clock; // @[:@89706.4]
  assign RetimeWrapper_109_reset = reset; // @[:@89707.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89709.4]
  assign RetimeWrapper_109_io_in = ~ x937; // @[package.scala 94:16:@89708.4]
  assign RetimeWrapper_110_clock = clock; // @[:@89718.4]
  assign RetimeWrapper_110_reset = reset; // @[:@89719.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89721.4]
  assign RetimeWrapper_110_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89720.4]
  assign x947_sum_1_clock = clock; // @[:@89745.4]
  assign x947_sum_1_reset = reset; // @[:@89746.4]
  assign x947_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@89747.4]
  assign x947_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@89748.4]
  assign x947_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89749.4]
  assign RetimeWrapper_111_clock = clock; // @[:@89755.4]
  assign RetimeWrapper_111_reset = reset; // @[:@89756.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89758.4]
  assign RetimeWrapper_111_io_in = ~ x945; // @[package.scala 94:16:@89757.4]
  assign RetimeWrapper_112_clock = clock; // @[:@89767.4]
  assign RetimeWrapper_112_reset = reset; // @[:@89768.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89770.4]
  assign RetimeWrapper_112_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89769.4]
  assign x952_sum_1_clock = clock; // @[:@89794.4]
  assign x952_sum_1_reset = reset; // @[:@89795.4]
  assign x952_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@89796.4]
  assign x952_sum_1_io_b = RetimeWrapper_61_io_out; // @[Math.scala 152:17:@89797.4]
  assign x952_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89798.4]
  assign RetimeWrapper_113_clock = clock; // @[:@89804.4]
  assign RetimeWrapper_113_reset = reset; // @[:@89805.4]
  assign RetimeWrapper_113_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89807.4]
  assign RetimeWrapper_113_io_in = ~ x950; // @[package.scala 94:16:@89806.4]
  assign RetimeWrapper_114_clock = clock; // @[:@89816.4]
  assign RetimeWrapper_114_reset = reset; // @[:@89817.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89819.4]
  assign RetimeWrapper_114_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89818.4]
  assign x957_sum_1_clock = clock; // @[:@89843.4]
  assign x957_sum_1_reset = reset; // @[:@89844.4]
  assign x957_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@89845.4]
  assign x957_sum_1_io_b = RetimeWrapper_67_io_out; // @[Math.scala 152:17:@89846.4]
  assign x957_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89847.4]
  assign RetimeWrapper_115_clock = clock; // @[:@89853.4]
  assign RetimeWrapper_115_reset = reset; // @[:@89854.4]
  assign RetimeWrapper_115_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89856.4]
  assign RetimeWrapper_115_io_in = ~ x955; // @[package.scala 94:16:@89855.4]
  assign RetimeWrapper_116_clock = clock; // @[:@89865.4]
  assign RetimeWrapper_116_reset = reset; // @[:@89866.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89868.4]
  assign RetimeWrapper_116_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89867.4]
  assign x962_sum_1_clock = clock; // @[:@89894.4]
  assign x962_sum_1_reset = reset; // @[:@89895.4]
  assign x962_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@89896.4]
  assign x962_sum_1_io_b = RetimeWrapper_73_io_out; // @[Math.scala 152:17:@89897.4]
  assign x962_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89898.4]
  assign RetimeWrapper_117_clock = clock; // @[:@89904.4]
  assign RetimeWrapper_117_reset = reset; // @[:@89905.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89907.4]
  assign RetimeWrapper_117_io_in = ~ x960; // @[package.scala 94:16:@89906.4]
  assign RetimeWrapper_118_clock = clock; // @[:@89916.4]
  assign RetimeWrapper_118_reset = reset; // @[:@89917.4]
  assign RetimeWrapper_118_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89919.4]
  assign RetimeWrapper_118_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89918.4]
  assign x967_sum_1_clock = clock; // @[:@89943.4]
  assign x967_sum_1_reset = reset; // @[:@89944.4]
  assign x967_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@89945.4]
  assign x967_sum_1_io_b = RetimeWrapper_79_io_out; // @[Math.scala 152:17:@89946.4]
  assign x967_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89947.4]
  assign RetimeWrapper_119_clock = clock; // @[:@89953.4]
  assign RetimeWrapper_119_reset = reset; // @[:@89954.4]
  assign RetimeWrapper_119_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89956.4]
  assign RetimeWrapper_119_io_in = ~ x965; // @[package.scala 94:16:@89955.4]
  assign RetimeWrapper_120_clock = clock; // @[:@89965.4]
  assign RetimeWrapper_120_reset = reset; // @[:@89966.4]
  assign RetimeWrapper_120_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@89968.4]
  assign RetimeWrapper_120_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@89967.4]
  assign x972_sum_1_clock = clock; // @[:@89992.4]
  assign x972_sum_1_reset = reset; // @[:@89993.4]
  assign x972_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@89994.4]
  assign x972_sum_1_io_b = RetimeWrapper_85_io_out; // @[Math.scala 152:17:@89995.4]
  assign x972_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@89996.4]
  assign RetimeWrapper_121_clock = clock; // @[:@90002.4]
  assign RetimeWrapper_121_reset = reset; // @[:@90003.4]
  assign RetimeWrapper_121_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90005.4]
  assign RetimeWrapper_121_io_in = ~ x970; // @[package.scala 94:16:@90004.4]
  assign RetimeWrapper_122_clock = clock; // @[:@90014.4]
  assign RetimeWrapper_122_reset = reset; // @[:@90015.4]
  assign RetimeWrapper_122_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90017.4]
  assign RetimeWrapper_122_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90016.4]
  assign RetimeWrapper_123_clock = clock; // @[:@90035.4]
  assign RetimeWrapper_123_reset = reset; // @[:@90036.4]
  assign RetimeWrapper_123_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90038.4]
  assign RetimeWrapper_123_io_in = RetimeWrapper_90_io_out; // @[package.scala 94:16:@90037.4]
  assign RetimeWrapper_124_clock = clock; // @[:@90050.4]
  assign RetimeWrapper_124_reset = reset; // @[:@90051.4]
  assign RetimeWrapper_124_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90053.4]
  assign RetimeWrapper_124_io_in = x1245_sum_1_io_result; // @[package.scala 94:16:@90052.4]
  assign x977_sum_1_clock = clock; // @[:@90059.4]
  assign x977_sum_1_reset = reset; // @[:@90060.4]
  assign x977_sum_1_io_a = RetimeWrapper_124_io_out; // @[Math.scala 151:17:@90061.4]
  assign x977_sum_1_io_b = RetimeWrapper_92_io_out; // @[Math.scala 152:17:@90062.4]
  assign x977_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90063.4]
  assign RetimeWrapper_125_clock = clock; // @[:@90069.4]
  assign RetimeWrapper_125_reset = reset; // @[:@90070.4]
  assign RetimeWrapper_125_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90072.4]
  assign RetimeWrapper_125_io_in = x977_sum_1_io_result; // @[package.scala 94:16:@90071.4]
  assign RetimeWrapper_126_clock = clock; // @[:@90078.4]
  assign RetimeWrapper_126_reset = reset; // @[:@90079.4]
  assign RetimeWrapper_126_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90081.4]
  assign RetimeWrapper_126_io_in = ~ x975; // @[package.scala 94:16:@90080.4]
  assign RetimeWrapper_127_clock = clock; // @[:@90090.4]
  assign RetimeWrapper_127_reset = reset; // @[:@90091.4]
  assign RetimeWrapper_127_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90093.4]
  assign RetimeWrapper_127_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90092.4]
  assign x982_sum_1_clock = clock; // @[:@90117.4]
  assign x982_sum_1_reset = reset; // @[:@90118.4]
  assign x982_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@90119.4]
  assign x982_sum_1_io_b = x921_div_1_io_result; // @[Math.scala 152:17:@90120.4]
  assign x982_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90121.4]
  assign RetimeWrapper_128_clock = clock; // @[:@90127.4]
  assign RetimeWrapper_128_reset = reset; // @[:@90128.4]
  assign RetimeWrapper_128_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90130.4]
  assign RetimeWrapper_128_io_in = ~ x980; // @[package.scala 94:16:@90129.4]
  assign RetimeWrapper_129_clock = clock; // @[:@90139.4]
  assign RetimeWrapper_129_reset = reset; // @[:@90140.4]
  assign RetimeWrapper_129_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90142.4]
  assign RetimeWrapper_129_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90141.4]
  assign x987_sum_1_clock = clock; // @[:@90166.4]
  assign x987_sum_1_reset = reset; // @[:@90167.4]
  assign x987_sum_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@90168.4]
  assign x987_sum_1_io_b = x930_div_1_io_result; // @[Math.scala 152:17:@90169.4]
  assign x987_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90170.4]
  assign RetimeWrapper_130_clock = clock; // @[:@90176.4]
  assign RetimeWrapper_130_reset = reset; // @[:@90177.4]
  assign RetimeWrapper_130_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90179.4]
  assign RetimeWrapper_130_io_in = ~ x985; // @[package.scala 94:16:@90178.4]
  assign RetimeWrapper_131_clock = clock; // @[:@90188.4]
  assign RetimeWrapper_131_reset = reset; // @[:@90189.4]
  assign RetimeWrapper_131_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90191.4]
  assign RetimeWrapper_131_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90190.4]
  assign x990_rdrow_1_clock = clock; // @[:@90211.4]
  assign x990_rdrow_1_reset = reset; // @[:@90212.4]
  assign x990_rdrow_1_io_a = RetimeWrapper_39_io_out; // @[Math.scala 192:17:@90213.4]
  assign x990_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@90214.4]
  assign x990_rdrow_1_io_flow = io_in_x745_TREADY; // @[Math.scala 194:20:@90215.4]
  assign RetimeWrapper_132_clock = clock; // @[:@90228.4]
  assign RetimeWrapper_132_reset = reset; // @[:@90229.4]
  assign RetimeWrapper_132_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@90232.4]
  assign RetimeWrapper_132_io_in = $unsigned(_T_1730); // @[package.scala 94:16:@90231.4]
  assign RetimeWrapper_133_clock = clock; // @[:@90246.4]
  assign RetimeWrapper_133_reset = reset; // @[:@90247.4]
  assign RetimeWrapper_133_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@90249.4]
  assign RetimeWrapper_133_io_in = $signed(_T_1727) < $signed(32'sh0); // @[package.scala 94:16:@90248.4]
  assign x1250_sum_1_clock = clock; // @[:@90291.4]
  assign x1250_sum_1_reset = reset; // @[:@90292.4]
  assign x1250_sum_1_io_a = _T_1775[31:0]; // @[Math.scala 151:17:@90293.4]
  assign x1250_sum_1_io_b = _T_1779[31:0]; // @[Math.scala 152:17:@90294.4]
  assign x1250_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90295.4]
  assign RetimeWrapper_134_clock = clock; // @[:@90301.4]
  assign RetimeWrapper_134_reset = reset; // @[:@90302.4]
  assign RetimeWrapper_134_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90304.4]
  assign RetimeWrapper_134_io_in = x1250_sum_1_io_result; // @[package.scala 94:16:@90303.4]
  assign x998_sum_1_clock = clock; // @[:@90312.4]
  assign x998_sum_1_reset = reset; // @[:@90313.4]
  assign x998_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90314.4]
  assign x998_sum_1_io_b = RetimeWrapper_46_io_out; // @[Math.scala 152:17:@90315.4]
  assign x998_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90316.4]
  assign RetimeWrapper_135_clock = clock; // @[:@90322.4]
  assign RetimeWrapper_135_reset = reset; // @[:@90323.4]
  assign RetimeWrapper_135_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90325.4]
  assign RetimeWrapper_135_io_in = ~ x993; // @[package.scala 94:16:@90324.4]
  assign RetimeWrapper_136_clock = clock; // @[:@90331.4]
  assign RetimeWrapper_136_reset = reset; // @[:@90332.4]
  assign RetimeWrapper_136_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90334.4]
  assign RetimeWrapper_136_io_in = $unsigned(_T_1760); // @[package.scala 94:16:@90333.4]
  assign RetimeWrapper_137_clock = clock; // @[:@90343.4]
  assign RetimeWrapper_137_reset = reset; // @[:@90344.4]
  assign RetimeWrapper_137_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90346.4]
  assign RetimeWrapper_137_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90345.4]
  assign x1003_sum_1_clock = clock; // @[:@90370.4]
  assign x1003_sum_1_reset = reset; // @[:@90371.4]
  assign x1003_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90372.4]
  assign x1003_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@90373.4]
  assign x1003_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90374.4]
  assign RetimeWrapper_138_clock = clock; // @[:@90380.4]
  assign RetimeWrapper_138_reset = reset; // @[:@90381.4]
  assign RetimeWrapper_138_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90383.4]
  assign RetimeWrapper_138_io_in = ~ x1001; // @[package.scala 94:16:@90382.4]
  assign RetimeWrapper_139_clock = clock; // @[:@90392.4]
  assign RetimeWrapper_139_reset = reset; // @[:@90393.4]
  assign RetimeWrapper_139_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90395.4]
  assign RetimeWrapper_139_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90394.4]
  assign x1008_sum_1_clock = clock; // @[:@90419.4]
  assign x1008_sum_1_reset = reset; // @[:@90420.4]
  assign x1008_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90421.4]
  assign x1008_sum_1_io_b = RetimeWrapper_61_io_out; // @[Math.scala 152:17:@90422.4]
  assign x1008_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90423.4]
  assign RetimeWrapper_140_clock = clock; // @[:@90429.4]
  assign RetimeWrapper_140_reset = reset; // @[:@90430.4]
  assign RetimeWrapper_140_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90432.4]
  assign RetimeWrapper_140_io_in = ~ x1006; // @[package.scala 94:16:@90431.4]
  assign RetimeWrapper_141_clock = clock; // @[:@90441.4]
  assign RetimeWrapper_141_reset = reset; // @[:@90442.4]
  assign RetimeWrapper_141_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90444.4]
  assign RetimeWrapper_141_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90443.4]
  assign x1013_sum_1_clock = clock; // @[:@90468.4]
  assign x1013_sum_1_reset = reset; // @[:@90469.4]
  assign x1013_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90470.4]
  assign x1013_sum_1_io_b = RetimeWrapper_67_io_out; // @[Math.scala 152:17:@90471.4]
  assign x1013_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90472.4]
  assign RetimeWrapper_142_clock = clock; // @[:@90478.4]
  assign RetimeWrapper_142_reset = reset; // @[:@90479.4]
  assign RetimeWrapper_142_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90481.4]
  assign RetimeWrapper_142_io_in = ~ x1011; // @[package.scala 94:16:@90480.4]
  assign RetimeWrapper_143_clock = clock; // @[:@90490.4]
  assign RetimeWrapper_143_reset = reset; // @[:@90491.4]
  assign RetimeWrapper_143_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90493.4]
  assign RetimeWrapper_143_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90492.4]
  assign x1018_sum_1_clock = clock; // @[:@90517.4]
  assign x1018_sum_1_reset = reset; // @[:@90518.4]
  assign x1018_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90519.4]
  assign x1018_sum_1_io_b = RetimeWrapper_73_io_out; // @[Math.scala 152:17:@90520.4]
  assign x1018_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90521.4]
  assign RetimeWrapper_144_clock = clock; // @[:@90527.4]
  assign RetimeWrapper_144_reset = reset; // @[:@90528.4]
  assign RetimeWrapper_144_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90530.4]
  assign RetimeWrapper_144_io_in = ~ x1016; // @[package.scala 94:16:@90529.4]
  assign RetimeWrapper_145_clock = clock; // @[:@90539.4]
  assign RetimeWrapper_145_reset = reset; // @[:@90540.4]
  assign RetimeWrapper_145_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90542.4]
  assign RetimeWrapper_145_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90541.4]
  assign x1023_sum_1_clock = clock; // @[:@90566.4]
  assign x1023_sum_1_reset = reset; // @[:@90567.4]
  assign x1023_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90568.4]
  assign x1023_sum_1_io_b = RetimeWrapper_79_io_out; // @[Math.scala 152:17:@90569.4]
  assign x1023_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90570.4]
  assign RetimeWrapper_146_clock = clock; // @[:@90576.4]
  assign RetimeWrapper_146_reset = reset; // @[:@90577.4]
  assign RetimeWrapper_146_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90579.4]
  assign RetimeWrapper_146_io_in = ~ x1021; // @[package.scala 94:16:@90578.4]
  assign RetimeWrapper_147_clock = clock; // @[:@90588.4]
  assign RetimeWrapper_147_reset = reset; // @[:@90589.4]
  assign RetimeWrapper_147_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90591.4]
  assign RetimeWrapper_147_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90590.4]
  assign x1028_sum_1_clock = clock; // @[:@90615.4]
  assign x1028_sum_1_reset = reset; // @[:@90616.4]
  assign x1028_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90617.4]
  assign x1028_sum_1_io_b = RetimeWrapper_85_io_out; // @[Math.scala 152:17:@90618.4]
  assign x1028_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90619.4]
  assign RetimeWrapper_148_clock = clock; // @[:@90625.4]
  assign RetimeWrapper_148_reset = reset; // @[:@90626.4]
  assign RetimeWrapper_148_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90628.4]
  assign RetimeWrapper_148_io_in = ~ x1026; // @[package.scala 94:16:@90627.4]
  assign RetimeWrapper_149_clock = clock; // @[:@90637.4]
  assign RetimeWrapper_149_reset = reset; // @[:@90638.4]
  assign RetimeWrapper_149_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90640.4]
  assign RetimeWrapper_149_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90639.4]
  assign RetimeWrapper_150_clock = clock; // @[:@90664.4]
  assign RetimeWrapper_150_reset = reset; // @[:@90665.4]
  assign RetimeWrapper_150_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90667.4]
  assign RetimeWrapper_150_io_in = x1250_sum_1_io_result; // @[package.scala 94:16:@90666.4]
  assign x1033_sum_1_clock = clock; // @[:@90673.4]
  assign x1033_sum_1_reset = reset; // @[:@90674.4]
  assign x1033_sum_1_io_a = RetimeWrapper_150_io_out; // @[Math.scala 151:17:@90675.4]
  assign x1033_sum_1_io_b = RetimeWrapper_92_io_out; // @[Math.scala 152:17:@90676.4]
  assign x1033_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90677.4]
  assign RetimeWrapper_151_clock = clock; // @[:@90683.4]
  assign RetimeWrapper_151_reset = reset; // @[:@90684.4]
  assign RetimeWrapper_151_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90686.4]
  assign RetimeWrapper_151_io_in = ~ x1031; // @[package.scala 94:16:@90685.4]
  assign RetimeWrapper_152_clock = clock; // @[:@90692.4]
  assign RetimeWrapper_152_reset = reset; // @[:@90693.4]
  assign RetimeWrapper_152_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90695.4]
  assign RetimeWrapper_152_io_in = x1033_sum_1_io_result; // @[package.scala 94:16:@90694.4]
  assign RetimeWrapper_153_clock = clock; // @[:@90704.4]
  assign RetimeWrapper_153_reset = reset; // @[:@90705.4]
  assign RetimeWrapper_153_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90707.4]
  assign RetimeWrapper_153_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90706.4]
  assign x1038_sum_1_clock = clock; // @[:@90733.4]
  assign x1038_sum_1_reset = reset; // @[:@90734.4]
  assign x1038_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90735.4]
  assign x1038_sum_1_io_b = x921_div_1_io_result; // @[Math.scala 152:17:@90736.4]
  assign x1038_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90737.4]
  assign RetimeWrapper_154_clock = clock; // @[:@90743.4]
  assign RetimeWrapper_154_reset = reset; // @[:@90744.4]
  assign RetimeWrapper_154_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90746.4]
  assign RetimeWrapper_154_io_in = ~ x1036; // @[package.scala 94:16:@90745.4]
  assign RetimeWrapper_155_clock = clock; // @[:@90755.4]
  assign RetimeWrapper_155_reset = reset; // @[:@90756.4]
  assign RetimeWrapper_155_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90758.4]
  assign RetimeWrapper_155_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90757.4]
  assign x1043_sum_1_clock = clock; // @[:@90782.4]
  assign x1043_sum_1_reset = reset; // @[:@90783.4]
  assign x1043_sum_1_io_a = RetimeWrapper_134_io_out; // @[Math.scala 151:17:@90784.4]
  assign x1043_sum_1_io_b = x930_div_1_io_result; // @[Math.scala 152:17:@90785.4]
  assign x1043_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90786.4]
  assign RetimeWrapper_156_clock = clock; // @[:@90792.4]
  assign RetimeWrapper_156_reset = reset; // @[:@90793.4]
  assign RetimeWrapper_156_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90795.4]
  assign RetimeWrapper_156_io_in = ~ x1041; // @[package.scala 94:16:@90794.4]
  assign RetimeWrapper_157_clock = clock; // @[:@90804.4]
  assign RetimeWrapper_157_reset = reset; // @[:@90805.4]
  assign RetimeWrapper_157_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90807.4]
  assign RetimeWrapper_157_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@90806.4]
  assign RetimeWrapper_158_clock = clock; // @[:@90827.4]
  assign RetimeWrapper_158_reset = reset; // @[:@90828.4]
  assign RetimeWrapper_158_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@90830.4]
  assign RetimeWrapper_158_io_in = _GEN_8 << 1; // @[package.scala 94:16:@90829.4]
  assign RetimeWrapper_159_clock = clock; // @[:@90839.4]
  assign RetimeWrapper_159_reset = reset; // @[:@90840.4]
  assign RetimeWrapper_159_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@90842.4]
  assign RetimeWrapper_159_io_in = _GEN_9 << 1; // @[package.scala 94:16:@90841.4]
  assign RetimeWrapper_160_clock = clock; // @[:@90851.4]
  assign RetimeWrapper_160_reset = reset; // @[:@90852.4]
  assign RetimeWrapper_160_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@90854.4]
  assign RetimeWrapper_160_io_in = _GEN_10 << 2; // @[package.scala 94:16:@90853.4]
  assign RetimeWrapper_161_clock = clock; // @[:@90863.4]
  assign RetimeWrapper_161_reset = reset; // @[:@90864.4]
  assign RetimeWrapper_161_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@90866.4]
  assign RetimeWrapper_161_io_in = _GEN_11 << 1; // @[package.scala 94:16:@90865.4]
  assign RetimeWrapper_162_clock = clock; // @[:@90875.4]
  assign RetimeWrapper_162_reset = reset; // @[:@90876.4]
  assign RetimeWrapper_162_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@90878.4]
  assign RetimeWrapper_162_io_in = _GEN_12 << 1; // @[package.scala 94:16:@90877.4]
  assign RetimeWrapper_163_clock = clock; // @[:@90885.4]
  assign RetimeWrapper_163_reset = reset; // @[:@90886.4]
  assign RetimeWrapper_163_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90888.4]
  assign RetimeWrapper_163_io_in = x805_lb_0_io_rPort_18_output_0; // @[package.scala 94:16:@90887.4]
  assign x1051_x15_1_io_a = RetimeWrapper_163_io_out; // @[Math.scala 151:17:@90896.4]
  assign x1051_x15_1_io_b = _T_2090[7:0]; // @[Math.scala 152:17:@90897.4]
  assign RetimeWrapper_164_clock = clock; // @[:@90904.4]
  assign RetimeWrapper_164_reset = reset; // @[:@90905.4]
  assign RetimeWrapper_164_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90907.4]
  assign RetimeWrapper_164_io_in = x805_lb_0_io_rPort_6_output_0; // @[package.scala 94:16:@90906.4]
  assign x1052_x16_1_io_a = RetimeWrapper_164_io_out; // @[Math.scala 151:17:@90915.4]
  assign x1052_x16_1_io_b = _T_2096[7:0]; // @[Math.scala 152:17:@90916.4]
  assign x1053_x15_1_io_a = _T_2102[7:0]; // @[Math.scala 151:17:@90925.4]
  assign x1053_x15_1_io_b = _T_2108[7:0]; // @[Math.scala 152:17:@90926.4]
  assign RetimeWrapper_165_clock = clock; // @[:@90933.4]
  assign RetimeWrapper_165_reset = reset; // @[:@90934.4]
  assign RetimeWrapper_165_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90936.4]
  assign RetimeWrapper_165_io_in = x805_lb_0_io_rPort_23_output_0; // @[package.scala 94:16:@90935.4]
  assign x1054_x16_1_io_a = RetimeWrapper_165_io_out; // @[Math.scala 151:17:@90944.4]
  assign x1054_x16_1_io_b = _T_2114[7:0]; // @[Math.scala 152:17:@90945.4]
  assign x1055_x15_1_io_a = x1051_x15_1_io_result; // @[Math.scala 151:17:@90954.4]
  assign x1055_x15_1_io_b = x1052_x16_1_io_result; // @[Math.scala 152:17:@90955.4]
  assign x1056_x16_1_io_a = x1053_x15_1_io_result; // @[Math.scala 151:17:@90964.4]
  assign x1056_x16_1_io_b = x1054_x16_1_io_result; // @[Math.scala 152:17:@90965.4]
  assign x1057_x15_1_io_a = x1055_x15_1_io_result; // @[Math.scala 151:17:@90974.4]
  assign x1057_x15_1_io_b = x1056_x16_1_io_result; // @[Math.scala 152:17:@90975.4]
  assign RetimeWrapper_166_clock = clock; // @[:@90982.4]
  assign RetimeWrapper_166_reset = reset; // @[:@90983.4]
  assign RetimeWrapper_166_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@90985.4]
  assign RetimeWrapper_166_io_in = x805_lb_0_io_rPort_27_output_0; // @[package.scala 94:16:@90984.4]
  assign x1058_sum_1_clock = clock; // @[:@90991.4]
  assign x1058_sum_1_reset = reset; // @[:@90992.4]
  assign x1058_sum_1_io_a = x1057_x15_1_io_result; // @[Math.scala 151:17:@90993.4]
  assign x1058_sum_1_io_b = RetimeWrapper_166_io_out; // @[Math.scala 152:17:@90994.4]
  assign x1058_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@90995.4]
  assign RetimeWrapper_167_clock = clock; // @[:@91010.4]
  assign RetimeWrapper_167_reset = reset; // @[:@91011.4]
  assign RetimeWrapper_167_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91013.4]
  assign RetimeWrapper_167_io_in = _GEN_13 << 1; // @[package.scala 94:16:@91012.4]
  assign RetimeWrapper_168_clock = clock; // @[:@91022.4]
  assign RetimeWrapper_168_reset = reset; // @[:@91023.4]
  assign RetimeWrapper_168_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91025.4]
  assign RetimeWrapper_168_io_in = _GEN_14 << 1; // @[package.scala 94:16:@91024.4]
  assign RetimeWrapper_169_clock = clock; // @[:@91034.4]
  assign RetimeWrapper_169_reset = reset; // @[:@91035.4]
  assign RetimeWrapper_169_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91037.4]
  assign RetimeWrapper_169_io_in = _GEN_15 << 2; // @[package.scala 94:16:@91036.4]
  assign RetimeWrapper_170_clock = clock; // @[:@91046.4]
  assign RetimeWrapper_170_reset = reset; // @[:@91047.4]
  assign RetimeWrapper_170_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91049.4]
  assign RetimeWrapper_170_io_in = _GEN_16 << 1; // @[package.scala 94:16:@91048.4]
  assign RetimeWrapper_171_clock = clock; // @[:@91058.4]
  assign RetimeWrapper_171_reset = reset; // @[:@91059.4]
  assign RetimeWrapper_171_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91061.4]
  assign RetimeWrapper_171_io_in = _GEN_17 << 1; // @[package.scala 94:16:@91060.4]
  assign RetimeWrapper_172_clock = clock; // @[:@91068.4]
  assign RetimeWrapper_172_reset = reset; // @[:@91069.4]
  assign RetimeWrapper_172_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91071.4]
  assign RetimeWrapper_172_io_in = x805_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@91070.4]
  assign x1065_x15_1_io_a = RetimeWrapper_172_io_out; // @[Math.scala 151:17:@91079.4]
  assign x1065_x15_1_io_b = _T_2166[7:0]; // @[Math.scala 152:17:@91080.4]
  assign RetimeWrapper_173_clock = clock; // @[:@91087.4]
  assign RetimeWrapper_173_reset = reset; // @[:@91088.4]
  assign RetimeWrapper_173_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91090.4]
  assign RetimeWrapper_173_io_in = x805_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@91089.4]
  assign x1066_x16_1_io_a = RetimeWrapper_173_io_out; // @[Math.scala 151:17:@91098.4]
  assign x1066_x16_1_io_b = _T_2172[7:0]; // @[Math.scala 152:17:@91099.4]
  assign x1067_x15_1_io_a = _T_2178[7:0]; // @[Math.scala 151:17:@91108.4]
  assign x1067_x15_1_io_b = _T_2184[7:0]; // @[Math.scala 152:17:@91109.4]
  assign RetimeWrapper_174_clock = clock; // @[:@91116.4]
  assign RetimeWrapper_174_reset = reset; // @[:@91117.4]
  assign RetimeWrapper_174_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91119.4]
  assign RetimeWrapper_174_io_in = x805_lb_0_io_rPort_26_output_0; // @[package.scala 94:16:@91118.4]
  assign x1068_x16_1_io_a = RetimeWrapper_174_io_out; // @[Math.scala 151:17:@91127.4]
  assign x1068_x16_1_io_b = _T_2190[7:0]; // @[Math.scala 152:17:@91128.4]
  assign x1069_x15_1_io_a = x1065_x15_1_io_result; // @[Math.scala 151:17:@91137.4]
  assign x1069_x15_1_io_b = x1066_x16_1_io_result; // @[Math.scala 152:17:@91138.4]
  assign x1070_x16_1_io_a = x1067_x15_1_io_result; // @[Math.scala 151:17:@91147.4]
  assign x1070_x16_1_io_b = x1068_x16_1_io_result; // @[Math.scala 152:17:@91148.4]
  assign x1071_x15_1_io_a = x1069_x15_1_io_result; // @[Math.scala 151:17:@91157.4]
  assign x1071_x15_1_io_b = x1070_x16_1_io_result; // @[Math.scala 152:17:@91158.4]
  assign RetimeWrapper_175_clock = clock; // @[:@91165.4]
  assign RetimeWrapper_175_reset = reset; // @[:@91166.4]
  assign RetimeWrapper_175_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91168.4]
  assign RetimeWrapper_175_io_in = x805_lb_0_io_rPort_29_output_0; // @[package.scala 94:16:@91167.4]
  assign x1072_sum_1_clock = clock; // @[:@91174.4]
  assign x1072_sum_1_reset = reset; // @[:@91175.4]
  assign x1072_sum_1_io_a = x1071_x15_1_io_result; // @[Math.scala 151:17:@91176.4]
  assign x1072_sum_1_io_b = RetimeWrapper_175_io_out; // @[Math.scala 152:17:@91177.4]
  assign x1072_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@91178.4]
  assign RetimeWrapper_176_clock = clock; // @[:@91193.4]
  assign RetimeWrapper_176_reset = reset; // @[:@91194.4]
  assign RetimeWrapper_176_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91196.4]
  assign RetimeWrapper_176_io_in = _GEN_18 << 1; // @[package.scala 94:16:@91195.4]
  assign RetimeWrapper_177_clock = clock; // @[:@91207.4]
  assign RetimeWrapper_177_reset = reset; // @[:@91208.4]
  assign RetimeWrapper_177_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91210.4]
  assign RetimeWrapper_177_io_in = _GEN_19 << 2; // @[package.scala 94:16:@91209.4]
  assign RetimeWrapper_178_clock = clock; // @[:@91219.4]
  assign RetimeWrapper_178_reset = reset; // @[:@91220.4]
  assign RetimeWrapper_178_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91222.4]
  assign RetimeWrapper_178_io_in = _GEN_20 << 1; // @[package.scala 94:16:@91221.4]
  assign RetimeWrapper_179_clock = clock; // @[:@91231.4]
  assign RetimeWrapper_179_reset = reset; // @[:@91232.4]
  assign RetimeWrapper_179_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91234.4]
  assign RetimeWrapper_179_io_in = _GEN_21 << 1; // @[package.scala 94:16:@91233.4]
  assign x1078_x15_1_io_a = RetimeWrapper_164_io_out; // @[Math.scala 151:17:@91243.4]
  assign x1078_x15_1_io_b = _T_2242[7:0]; // @[Math.scala 152:17:@91244.4]
  assign RetimeWrapper_180_clock = clock; // @[:@91251.4]
  assign RetimeWrapper_180_reset = reset; // @[:@91252.4]
  assign RetimeWrapper_180_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91254.4]
  assign RetimeWrapper_180_io_in = x805_lb_0_io_rPort_21_output_0; // @[package.scala 94:16:@91253.4]
  assign x1079_x16_1_io_a = RetimeWrapper_180_io_out; // @[Math.scala 151:17:@91262.4]
  assign x1079_x16_1_io_b = _T_2108[7:0]; // @[Math.scala 152:17:@91263.4]
  assign x1080_x15_1_io_a = _T_2250[7:0]; // @[Math.scala 151:17:@91272.4]
  assign x1080_x15_1_io_b = _T_2256[7:0]; // @[Math.scala 152:17:@91273.4]
  assign x1081_x16_1_io_a = RetimeWrapper_166_io_out; // @[Math.scala 151:17:@91282.4]
  assign x1081_x16_1_io_b = _T_2262[7:0]; // @[Math.scala 152:17:@91283.4]
  assign x1082_x15_1_io_a = x1078_x15_1_io_result; // @[Math.scala 151:17:@91292.4]
  assign x1082_x15_1_io_b = x1079_x16_1_io_result; // @[Math.scala 152:17:@91293.4]
  assign x1083_x16_1_io_a = x1080_x15_1_io_result; // @[Math.scala 151:17:@91302.4]
  assign x1083_x16_1_io_b = x1081_x16_1_io_result; // @[Math.scala 152:17:@91303.4]
  assign x1084_x15_1_io_a = x1082_x15_1_io_result; // @[Math.scala 151:17:@91312.4]
  assign x1084_x15_1_io_b = x1083_x16_1_io_result; // @[Math.scala 152:17:@91313.4]
  assign RetimeWrapper_181_clock = clock; // @[:@91320.4]
  assign RetimeWrapper_181_reset = reset; // @[:@91321.4]
  assign RetimeWrapper_181_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91323.4]
  assign RetimeWrapper_181_io_in = x805_lb_0_io_rPort_24_output_0; // @[package.scala 94:16:@91322.4]
  assign x1085_sum_1_clock = clock; // @[:@91329.4]
  assign x1085_sum_1_reset = reset; // @[:@91330.4]
  assign x1085_sum_1_io_a = x1084_x15_1_io_result; // @[Math.scala 151:17:@91331.4]
  assign x1085_sum_1_io_b = RetimeWrapper_181_io_out; // @[Math.scala 152:17:@91332.4]
  assign x1085_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@91333.4]
  assign RetimeWrapper_182_clock = clock; // @[:@91348.4]
  assign RetimeWrapper_182_reset = reset; // @[:@91349.4]
  assign RetimeWrapper_182_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91351.4]
  assign RetimeWrapper_182_io_in = _GEN_22 << 1; // @[package.scala 94:16:@91350.4]
  assign RetimeWrapper_183_clock = clock; // @[:@91360.4]
  assign RetimeWrapper_183_reset = reset; // @[:@91361.4]
  assign RetimeWrapper_183_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91363.4]
  assign RetimeWrapper_183_io_in = _GEN_23 << 2; // @[package.scala 94:16:@91362.4]
  assign RetimeWrapper_184_clock = clock; // @[:@91372.4]
  assign RetimeWrapper_184_reset = reset; // @[:@91373.4]
  assign RetimeWrapper_184_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91375.4]
  assign RetimeWrapper_184_io_in = _GEN_24 << 1; // @[package.scala 94:16:@91374.4]
  assign RetimeWrapper_185_clock = clock; // @[:@91384.4]
  assign RetimeWrapper_185_reset = reset; // @[:@91385.4]
  assign RetimeWrapper_185_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91387.4]
  assign RetimeWrapper_185_io_in = _GEN_25 << 1; // @[package.scala 94:16:@91386.4]
  assign x1091_x15_1_io_a = RetimeWrapper_173_io_out; // @[Math.scala 151:17:@91396.4]
  assign x1091_x15_1_io_b = _T_2308[7:0]; // @[Math.scala 152:17:@91397.4]
  assign RetimeWrapper_186_clock = clock; // @[:@91404.4]
  assign RetimeWrapper_186_reset = reset; // @[:@91405.4]
  assign RetimeWrapper_186_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91407.4]
  assign RetimeWrapper_186_io_in = x805_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@91406.4]
  assign x1092_x16_1_io_a = RetimeWrapper_186_io_out; // @[Math.scala 151:17:@91415.4]
  assign x1092_x16_1_io_b = _T_2184[7:0]; // @[Math.scala 152:17:@91416.4]
  assign x1093_x15_1_io_a = _T_2314[7:0]; // @[Math.scala 151:17:@91425.4]
  assign x1093_x15_1_io_b = _T_2320[7:0]; // @[Math.scala 152:17:@91426.4]
  assign x1094_x16_1_io_a = RetimeWrapper_175_io_out; // @[Math.scala 151:17:@91435.4]
  assign x1094_x16_1_io_b = _T_2326[7:0]; // @[Math.scala 152:17:@91436.4]
  assign x1095_x15_1_io_a = x1091_x15_1_io_result; // @[Math.scala 151:17:@91445.4]
  assign x1095_x15_1_io_b = x1092_x16_1_io_result; // @[Math.scala 152:17:@91446.4]
  assign x1096_x16_1_io_a = x1093_x15_1_io_result; // @[Math.scala 151:17:@91455.4]
  assign x1096_x16_1_io_b = x1094_x16_1_io_result; // @[Math.scala 152:17:@91456.4]
  assign x1097_x15_1_io_a = x1095_x15_1_io_result; // @[Math.scala 151:17:@91465.4]
  assign x1097_x15_1_io_b = x1096_x16_1_io_result; // @[Math.scala 152:17:@91466.4]
  assign RetimeWrapper_187_clock = clock; // @[:@91473.4]
  assign RetimeWrapper_187_reset = reset; // @[:@91474.4]
  assign RetimeWrapper_187_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91476.4]
  assign RetimeWrapper_187_io_in = x805_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@91475.4]
  assign x1098_sum_1_clock = clock; // @[:@91482.4]
  assign x1098_sum_1_reset = reset; // @[:@91483.4]
  assign x1098_sum_1_io_a = x1097_x15_1_io_result; // @[Math.scala 151:17:@91484.4]
  assign x1098_sum_1_io_b = RetimeWrapper_187_io_out; // @[Math.scala 152:17:@91485.4]
  assign x1098_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@91486.4]
  assign RetimeWrapper_188_clock = clock; // @[:@91501.4]
  assign RetimeWrapper_188_reset = reset; // @[:@91502.4]
  assign RetimeWrapper_188_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91504.4]
  assign RetimeWrapper_188_io_in = _GEN_26 << 1; // @[package.scala 94:16:@91503.4]
  assign RetimeWrapper_189_clock = clock; // @[:@91513.4]
  assign RetimeWrapper_189_reset = reset; // @[:@91514.4]
  assign RetimeWrapper_189_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91516.4]
  assign RetimeWrapper_189_io_in = _GEN_27 << 2; // @[package.scala 94:16:@91515.4]
  assign RetimeWrapper_190_clock = clock; // @[:@91525.4]
  assign RetimeWrapper_190_reset = reset; // @[:@91526.4]
  assign RetimeWrapper_190_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91528.4]
  assign RetimeWrapper_190_io_in = _GEN_28 << 1; // @[package.scala 94:16:@91527.4]
  assign RetimeWrapper_191_clock = clock; // @[:@91537.4]
  assign RetimeWrapper_191_reset = reset; // @[:@91538.4]
  assign RetimeWrapper_191_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91540.4]
  assign RetimeWrapper_191_io_in = _GEN_29 << 1; // @[package.scala 94:16:@91539.4]
  assign x1104_x15_1_io_a = RetimeWrapper_180_io_out; // @[Math.scala 151:17:@91549.4]
  assign x1104_x15_1_io_b = _T_2372[7:0]; // @[Math.scala 152:17:@91550.4]
  assign RetimeWrapper_192_clock = clock; // @[:@91557.4]
  assign RetimeWrapper_192_reset = reset; // @[:@91558.4]
  assign RetimeWrapper_192_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91560.4]
  assign RetimeWrapper_192_io_in = x805_lb_0_io_rPort_25_output_0; // @[package.scala 94:16:@91559.4]
  assign x1105_x16_1_io_a = RetimeWrapper_192_io_out; // @[Math.scala 151:17:@91568.4]
  assign x1105_x16_1_io_b = _T_2256[7:0]; // @[Math.scala 152:17:@91569.4]
  assign x1106_x15_1_io_a = _T_2378[7:0]; // @[Math.scala 151:17:@91578.4]
  assign x1106_x15_1_io_b = _T_2384[7:0]; // @[Math.scala 152:17:@91579.4]
  assign x1107_x16_1_io_a = RetimeWrapper_181_io_out; // @[Math.scala 151:17:@91588.4]
  assign x1107_x16_1_io_b = _T_2390[7:0]; // @[Math.scala 152:17:@91589.4]
  assign x1108_x15_1_io_a = x1104_x15_1_io_result; // @[Math.scala 151:17:@91598.4]
  assign x1108_x15_1_io_b = x1105_x16_1_io_result; // @[Math.scala 152:17:@91599.4]
  assign x1109_x16_1_io_a = x1106_x15_1_io_result; // @[Math.scala 151:17:@91608.4]
  assign x1109_x16_1_io_b = x1107_x16_1_io_result; // @[Math.scala 152:17:@91609.4]
  assign x1110_x15_1_io_a = x1108_x15_1_io_result; // @[Math.scala 151:17:@91618.4]
  assign x1110_x15_1_io_b = x1109_x16_1_io_result; // @[Math.scala 152:17:@91619.4]
  assign RetimeWrapper_193_clock = clock; // @[:@91626.4]
  assign RetimeWrapper_193_reset = reset; // @[:@91627.4]
  assign RetimeWrapper_193_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91629.4]
  assign RetimeWrapper_193_io_in = x805_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@91628.4]
  assign x1111_sum_1_clock = clock; // @[:@91635.4]
  assign x1111_sum_1_reset = reset; // @[:@91636.4]
  assign x1111_sum_1_io_a = x1110_x15_1_io_result; // @[Math.scala 151:17:@91637.4]
  assign x1111_sum_1_io_b = RetimeWrapper_193_io_out; // @[Math.scala 152:17:@91638.4]
  assign x1111_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@91639.4]
  assign RetimeWrapper_194_clock = clock; // @[:@91654.4]
  assign RetimeWrapper_194_reset = reset; // @[:@91655.4]
  assign RetimeWrapper_194_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91657.4]
  assign RetimeWrapper_194_io_in = _GEN_30 << 1; // @[package.scala 94:16:@91656.4]
  assign RetimeWrapper_195_clock = clock; // @[:@91666.4]
  assign RetimeWrapper_195_reset = reset; // @[:@91667.4]
  assign RetimeWrapper_195_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91669.4]
  assign RetimeWrapper_195_io_in = _GEN_31 << 2; // @[package.scala 94:16:@91668.4]
  assign RetimeWrapper_196_clock = clock; // @[:@91678.4]
  assign RetimeWrapper_196_reset = reset; // @[:@91679.4]
  assign RetimeWrapper_196_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91681.4]
  assign RetimeWrapper_196_io_in = _GEN_32 << 1; // @[package.scala 94:16:@91680.4]
  assign RetimeWrapper_197_clock = clock; // @[:@91690.4]
  assign RetimeWrapper_197_reset = reset; // @[:@91691.4]
  assign RetimeWrapper_197_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91693.4]
  assign RetimeWrapper_197_io_in = _GEN_33 << 1; // @[package.scala 94:16:@91692.4]
  assign x1117_x15_1_io_a = RetimeWrapper_186_io_out; // @[Math.scala 151:17:@91702.4]
  assign x1117_x15_1_io_b = _T_2436[7:0]; // @[Math.scala 152:17:@91703.4]
  assign RetimeWrapper_198_clock = clock; // @[:@91710.4]
  assign RetimeWrapper_198_reset = reset; // @[:@91711.4]
  assign RetimeWrapper_198_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91713.4]
  assign RetimeWrapper_198_io_in = x805_lb_0_io_rPort_22_output_0; // @[package.scala 94:16:@91712.4]
  assign x1118_x16_1_io_a = RetimeWrapper_198_io_out; // @[Math.scala 151:17:@91723.4]
  assign x1118_x16_1_io_b = _T_2320[7:0]; // @[Math.scala 152:17:@91724.4]
  assign x1119_x15_1_io_a = _T_2442[7:0]; // @[Math.scala 151:17:@91733.4]
  assign x1119_x15_1_io_b = _T_2448[7:0]; // @[Math.scala 152:17:@91734.4]
  assign x1120_x16_1_io_a = RetimeWrapper_187_io_out; // @[Math.scala 151:17:@91743.4]
  assign x1120_x16_1_io_b = _T_2454[7:0]; // @[Math.scala 152:17:@91744.4]
  assign x1121_x15_1_io_a = x1117_x15_1_io_result; // @[Math.scala 151:17:@91753.4]
  assign x1121_x15_1_io_b = x1118_x16_1_io_result; // @[Math.scala 152:17:@91754.4]
  assign x1122_x16_1_io_a = x1119_x15_1_io_result; // @[Math.scala 151:17:@91763.4]
  assign x1122_x16_1_io_b = x1120_x16_1_io_result; // @[Math.scala 152:17:@91764.4]
  assign x1123_x15_1_io_a = x1121_x15_1_io_result; // @[Math.scala 151:17:@91773.4]
  assign x1123_x15_1_io_b = x1122_x16_1_io_result; // @[Math.scala 152:17:@91774.4]
  assign RetimeWrapper_199_clock = clock; // @[:@91781.4]
  assign RetimeWrapper_199_reset = reset; // @[:@91782.4]
  assign RetimeWrapper_199_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91784.4]
  assign RetimeWrapper_199_io_in = x805_lb_0_io_rPort_16_output_0; // @[package.scala 94:16:@91783.4]
  assign x1124_sum_1_clock = clock; // @[:@91790.4]
  assign x1124_sum_1_reset = reset; // @[:@91791.4]
  assign x1124_sum_1_io_a = x1123_x15_1_io_result; // @[Math.scala 151:17:@91792.4]
  assign x1124_sum_1_io_b = RetimeWrapper_199_io_out; // @[Math.scala 152:17:@91793.4]
  assign x1124_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@91794.4]
  assign RetimeWrapper_200_clock = clock; // @[:@91809.4]
  assign RetimeWrapper_200_reset = reset; // @[:@91810.4]
  assign RetimeWrapper_200_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91812.4]
  assign RetimeWrapper_200_io_in = _GEN_34 << 1; // @[package.scala 94:16:@91811.4]
  assign RetimeWrapper_201_clock = clock; // @[:@91821.4]
  assign RetimeWrapper_201_reset = reset; // @[:@91822.4]
  assign RetimeWrapper_201_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91824.4]
  assign RetimeWrapper_201_io_in = _GEN_35 << 2; // @[package.scala 94:16:@91823.4]
  assign RetimeWrapper_202_clock = clock; // @[:@91833.4]
  assign RetimeWrapper_202_reset = reset; // @[:@91834.4]
  assign RetimeWrapper_202_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91836.4]
  assign RetimeWrapper_202_io_in = _GEN_36 << 1; // @[package.scala 94:16:@91835.4]
  assign RetimeWrapper_203_clock = clock; // @[:@91845.4]
  assign RetimeWrapper_203_reset = reset; // @[:@91846.4]
  assign RetimeWrapper_203_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91848.4]
  assign RetimeWrapper_203_io_in = _GEN_37 << 1; // @[package.scala 94:16:@91847.4]
  assign x1130_x15_1_io_a = RetimeWrapper_192_io_out; // @[Math.scala 151:17:@91857.4]
  assign x1130_x15_1_io_b = _T_2502[7:0]; // @[Math.scala 152:17:@91858.4]
  assign RetimeWrapper_204_clock = clock; // @[:@91865.4]
  assign RetimeWrapper_204_reset = reset; // @[:@91866.4]
  assign RetimeWrapper_204_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91868.4]
  assign RetimeWrapper_204_io_in = x805_lb_0_io_rPort_28_output_0; // @[package.scala 94:16:@91867.4]
  assign x1131_x16_1_io_a = RetimeWrapper_204_io_out; // @[Math.scala 151:17:@91876.4]
  assign x1131_x16_1_io_b = _T_2384[7:0]; // @[Math.scala 152:17:@91877.4]
  assign x1132_x15_1_io_a = _T_2508[7:0]; // @[Math.scala 151:17:@91886.4]
  assign x1132_x15_1_io_b = _T_2514[7:0]; // @[Math.scala 152:17:@91887.4]
  assign x1133_x16_1_io_a = RetimeWrapper_193_io_out; // @[Math.scala 151:17:@91896.4]
  assign x1133_x16_1_io_b = _T_2520[7:0]; // @[Math.scala 152:17:@91897.4]
  assign x1134_x15_1_io_a = x1130_x15_1_io_result; // @[Math.scala 151:17:@91906.4]
  assign x1134_x15_1_io_b = x1131_x16_1_io_result; // @[Math.scala 152:17:@91907.4]
  assign x1135_x16_1_io_a = x1132_x15_1_io_result; // @[Math.scala 151:17:@91916.4]
  assign x1135_x16_1_io_b = x1133_x16_1_io_result; // @[Math.scala 152:17:@91917.4]
  assign x1136_x15_1_io_a = x1134_x15_1_io_result; // @[Math.scala 151:17:@91926.4]
  assign x1136_x15_1_io_b = x1135_x16_1_io_result; // @[Math.scala 152:17:@91927.4]
  assign RetimeWrapper_205_clock = clock; // @[:@91934.4]
  assign RetimeWrapper_205_reset = reset; // @[:@91935.4]
  assign RetimeWrapper_205_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@91937.4]
  assign RetimeWrapper_205_io_in = x805_lb_0_io_rPort_7_output_0; // @[package.scala 94:16:@91936.4]
  assign x1137_sum_1_clock = clock; // @[:@91943.4]
  assign x1137_sum_1_reset = reset; // @[:@91944.4]
  assign x1137_sum_1_io_a = x1136_x15_1_io_result; // @[Math.scala 151:17:@91945.4]
  assign x1137_sum_1_io_b = RetimeWrapper_205_io_out; // @[Math.scala 152:17:@91946.4]
  assign x1137_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@91947.4]
  assign RetimeWrapper_206_clock = clock; // @[:@91962.4]
  assign RetimeWrapper_206_reset = reset; // @[:@91963.4]
  assign RetimeWrapper_206_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91965.4]
  assign RetimeWrapper_206_io_in = _GEN_38 << 1; // @[package.scala 94:16:@91964.4]
  assign RetimeWrapper_207_clock = clock; // @[:@91974.4]
  assign RetimeWrapper_207_reset = reset; // @[:@91975.4]
  assign RetimeWrapper_207_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91977.4]
  assign RetimeWrapper_207_io_in = _GEN_39 << 2; // @[package.scala 94:16:@91976.4]
  assign RetimeWrapper_208_clock = clock; // @[:@91986.4]
  assign RetimeWrapper_208_reset = reset; // @[:@91987.4]
  assign RetimeWrapper_208_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@91989.4]
  assign RetimeWrapper_208_io_in = _GEN_40 << 1; // @[package.scala 94:16:@91988.4]
  assign RetimeWrapper_209_clock = clock; // @[:@91998.4]
  assign RetimeWrapper_209_reset = reset; // @[:@91999.4]
  assign RetimeWrapper_209_io_flow = io_in_x745_TREADY; // @[package.scala 95:18:@92001.4]
  assign RetimeWrapper_209_io_in = _GEN_41 << 1; // @[package.scala 94:16:@92000.4]
  assign x1143_x15_1_io_a = RetimeWrapper_198_io_out; // @[Math.scala 151:17:@92010.4]
  assign x1143_x15_1_io_b = _T_2566[7:0]; // @[Math.scala 152:17:@92011.4]
  assign RetimeWrapper_210_clock = clock; // @[:@92018.4]
  assign RetimeWrapper_210_reset = reset; // @[:@92019.4]
  assign RetimeWrapper_210_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@92021.4]
  assign RetimeWrapper_210_io_in = x805_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@92020.4]
  assign x1144_x16_1_io_a = RetimeWrapper_210_io_out; // @[Math.scala 151:17:@92029.4]
  assign x1144_x16_1_io_b = _T_2448[7:0]; // @[Math.scala 152:17:@92030.4]
  assign x1145_x15_1_io_a = _T_2572[7:0]; // @[Math.scala 151:17:@92039.4]
  assign x1145_x15_1_io_b = _T_2578[7:0]; // @[Math.scala 152:17:@92040.4]
  assign x1146_x16_1_io_a = RetimeWrapper_199_io_out; // @[Math.scala 151:17:@92049.4]
  assign x1146_x16_1_io_b = _T_2584[7:0]; // @[Math.scala 152:17:@92050.4]
  assign x1147_x15_1_io_a = x1143_x15_1_io_result; // @[Math.scala 151:17:@92059.4]
  assign x1147_x15_1_io_b = x1144_x16_1_io_result; // @[Math.scala 152:17:@92060.4]
  assign x1148_x16_1_io_a = x1145_x15_1_io_result; // @[Math.scala 151:17:@92069.4]
  assign x1148_x16_1_io_b = x1146_x16_1_io_result; // @[Math.scala 152:17:@92070.4]
  assign x1149_x15_1_io_a = x1147_x15_1_io_result; // @[Math.scala 151:17:@92079.4]
  assign x1149_x15_1_io_b = x1148_x16_1_io_result; // @[Math.scala 152:17:@92080.4]
  assign RetimeWrapper_211_clock = clock; // @[:@92087.4]
  assign RetimeWrapper_211_reset = reset; // @[:@92088.4]
  assign RetimeWrapper_211_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@92090.4]
  assign RetimeWrapper_211_io_in = x805_lb_0_io_rPort_15_output_0; // @[package.scala 94:16:@92089.4]
  assign x1150_sum_1_clock = clock; // @[:@92096.4]
  assign x1150_sum_1_reset = reset; // @[:@92097.4]
  assign x1150_sum_1_io_a = x1149_x15_1_io_result; // @[Math.scala 151:17:@92098.4]
  assign x1150_sum_1_io_b = RetimeWrapper_211_io_out; // @[Math.scala 152:17:@92099.4]
  assign x1150_sum_1_io_flow = io_in_x745_TREADY; // @[Math.scala 153:20:@92100.4]
  assign RetimeWrapper_212_clock = clock; // @[:@92131.4]
  assign RetimeWrapper_212_reset = reset; // @[:@92132.4]
  assign RetimeWrapper_212_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@92134.4]
  assign RetimeWrapper_212_io_in = {_T_2645,_T_2642}; // @[package.scala 94:16:@92133.4]
  assign RetimeWrapper_213_clock = clock; // @[:@92140.4]
  assign RetimeWrapper_213_reset = reset; // @[:@92141.4]
  assign RetimeWrapper_213_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@92143.4]
  assign RetimeWrapper_213_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@92142.4]
  assign RetimeWrapper_214_clock = clock; // @[:@92149.4]
  assign RetimeWrapper_214_reset = reset; // @[:@92150.4]
  assign RetimeWrapper_214_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@92152.4]
  assign RetimeWrapper_214_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@92151.4]
  assign RetimeWrapper_215_clock = clock; // @[:@92158.4]
  assign RetimeWrapper_215_reset = reset; // @[:@92159.4]
  assign RetimeWrapper_215_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@92161.4]
  assign RetimeWrapper_215_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@92160.4]
endmodule
module x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1( // @[:@92179.2]
  input          clock, // @[:@92180.4]
  input          reset, // @[:@92181.4]
  output         io_in_x745_TVALID, // @[:@92182.4]
  input          io_in_x745_TREADY, // @[:@92182.4]
  output [255:0] io_in_x745_TDATA, // @[:@92182.4]
  input          io_in_x744_TVALID, // @[:@92182.4]
  output         io_in_x744_TREADY, // @[:@92182.4]
  input  [255:0] io_in_x744_TDATA, // @[:@92182.4]
  input  [7:0]   io_in_x744_TID, // @[:@92182.4]
  input  [7:0]   io_in_x744_TDEST, // @[:@92182.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@92182.4]
  input          io_sigsIn_smChildAcks_0, // @[:@92182.4]
  output         io_sigsOut_smDoneIn_0, // @[:@92182.4]
  input          io_rr // @[:@92182.4]
);
  wire  x798_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire  x798_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire  x798_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire  x798_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire [12:0] x798_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire [12:0] x798_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire  x798_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire  x798_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire  x798_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@92216.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@92304.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@92304.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@92304.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@92304.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@92304.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@92346.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@92346.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@92346.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@92346.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@92346.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@92354.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@92354.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@92354.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@92354.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@92354.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TVALID; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TREADY; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire [255:0] x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TDATA; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TREADY; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire [255:0] x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TDATA; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire [7:0] x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TID; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire [7:0] x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TDEST; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire [31:0] x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire [31:0] x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
  wire  _T_240; // @[package.scala 96:25:@92309.4 package.scala 96:25:@92310.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x1157_outr_UnitPipe.scala 69:67:@92315.4]
  wire  _T_253; // @[package.scala 96:25:@92351.4 package.scala 96:25:@92352.4]
  wire  _T_259; // @[package.scala 96:25:@92359.4 package.scala 96:25:@92360.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@92362.4]
  wire  x1156_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@92363.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@92371.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@92372.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@92384.4]
  x752_ctrchain x798_ctrchain ( // @[SpatialBlocks.scala 37:22:@92216.4]
    .clock(x798_ctrchain_clock),
    .reset(x798_ctrchain_reset),
    .io_input_reset(x798_ctrchain_io_input_reset),
    .io_input_enable(x798_ctrchain_io_input_enable),
    .io_output_counts_1(x798_ctrchain_io_output_counts_1),
    .io_output_counts_0(x798_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x798_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x798_ctrchain_io_output_oobs_1),
    .io_output_done(x798_ctrchain_io_output_done)
  );
  x1156_inr_Foreach_SAMPLER_BOX_sm x1156_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 32:18:@92276.4]
    .clock(x1156_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x1156_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x1156_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x1156_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x1156_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x1156_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x1156_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x1156_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x1156_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@92304.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@92346.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@92354.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1 x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1238:24:@92388.4]
    .clock(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x745_TVALID(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TVALID),
    .io_in_x745_TREADY(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TREADY),
    .io_in_x745_TDATA(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TDATA),
    .io_in_x744_TREADY(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TREADY),
    .io_in_x744_TDATA(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TDATA),
    .io_in_x744_TID(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TID),
    .io_in_x744_TDEST(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TDEST),
    .io_sigsIn_backpressure(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@92309.4 package.scala 96:25:@92310.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x744_TVALID | x1156_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x1157_outr_UnitPipe.scala 69:67:@92315.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@92351.4 package.scala 96:25:@92352.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@92359.4 package.scala 96:25:@92360.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@92362.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@92363.4]
  assign _T_264 = x1156_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@92371.4]
  assign _T_265 = ~ x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@92372.4]
  assign _T_272 = x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@92384.4]
  assign io_in_x745_TVALID = x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TVALID; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 48:23:@92447.4]
  assign io_in_x745_TDATA = x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TDATA; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 48:23:@92445.4]
  assign io_in_x744_TREADY = x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TREADY; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 49:23:@92455.4]
  assign io_sigsOut_smDoneIn_0 = x1156_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@92369.4]
  assign x798_ctrchain_clock = clock; // @[:@92217.4]
  assign x798_ctrchain_reset = reset; // @[:@92218.4]
  assign x798_ctrchain_io_input_reset = x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@92387.4]
  assign x798_ctrchain_io_input_enable = _T_272 & x1156_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@92339.4 SpatialBlocks.scala 159:42:@92386.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@92277.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@92278.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sm_io_enable = x1156_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x1156_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@92366.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x1157_outr_UnitPipe.scala 67:51:@92312.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@92368.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x745_TREADY | x1156_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@92340.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x1157_outr_UnitPipe.scala 71:49:@92318.4]
  assign RetimeWrapper_clock = clock; // @[:@92305.4]
  assign RetimeWrapper_reset = reset; // @[:@92306.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@92308.4]
  assign RetimeWrapper_io_in = x798_ctrchain_io_output_done; // @[package.scala 94:16:@92307.4]
  assign RetimeWrapper_1_clock = clock; // @[:@92347.4]
  assign RetimeWrapper_1_reset = reset; // @[:@92348.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@92350.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@92349.4]
  assign RetimeWrapper_2_clock = clock; // @[:@92355.4]
  assign RetimeWrapper_2_reset = reset; // @[:@92356.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@92358.4]
  assign RetimeWrapper_2_io_in = x1156_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@92357.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@92389.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@92390.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x745_TREADY = io_in_x745_TREADY; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 48:23:@92446.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TDATA = io_in_x744_TDATA; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 49:23:@92454.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TID = io_in_x744_TID; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 49:23:@92450.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x744_TDEST = io_in_x744_TDEST; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 49:23:@92449.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x745_TREADY | x1156_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1243:22:@92473.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1243:22:@92471.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x1156_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1243:22:@92469.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x798_ctrchain_io_output_counts_1[12]}},x798_ctrchain_io_output_counts_1}; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1243:22:@92464.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x798_ctrchain_io_output_counts_0[12]}},x798_ctrchain_io_output_counts_0}; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1243:22:@92463.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x798_ctrchain_io_output_oobs_0; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1243:22:@92461.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x798_ctrchain_io_output_oobs_1; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1243:22:@92462.4]
  assign x1156_inr_Foreach_SAMPLER_BOX_kernelx1156_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x1156_inr_Foreach_SAMPLER_BOX.scala 1242:18:@92457.4]
endmodule
module x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1( // @[:@92487.2]
  input          clock, // @[:@92488.4]
  input          reset, // @[:@92489.4]
  output         io_in_x745_TVALID, // @[:@92490.4]
  input          io_in_x745_TREADY, // @[:@92490.4]
  output [255:0] io_in_x745_TDATA, // @[:@92490.4]
  input          io_in_x744_TVALID, // @[:@92490.4]
  output         io_in_x744_TREADY, // @[:@92490.4]
  input  [255:0] io_in_x744_TDATA, // @[:@92490.4]
  input  [7:0]   io_in_x744_TID, // @[:@92490.4]
  input  [7:0]   io_in_x744_TDEST, // @[:@92490.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@92490.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@92490.4]
  input          io_sigsIn_smChildAcks_0, // @[:@92490.4]
  input          io_sigsIn_smChildAcks_1, // @[:@92490.4]
  output         io_sigsOut_smDoneIn_0, // @[:@92490.4]
  output         io_sigsOut_smDoneIn_1, // @[:@92490.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@92490.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@92490.4]
  input          io_rr // @[:@92490.4]
);
  wire  x747_fifoinraw_0_clock; // @[m_x747_fifoinraw_0.scala 27:17:@92504.4]
  wire  x747_fifoinraw_0_reset; // @[m_x747_fifoinraw_0.scala 27:17:@92504.4]
  wire  x748_fifoinpacked_0_clock; // @[m_x748_fifoinpacked_0.scala 27:17:@92528.4]
  wire  x748_fifoinpacked_0_reset; // @[m_x748_fifoinpacked_0.scala 27:17:@92528.4]
  wire  x748_fifoinpacked_0_io_wPort_0_en_0; // @[m_x748_fifoinpacked_0.scala 27:17:@92528.4]
  wire  x748_fifoinpacked_0_io_full; // @[m_x748_fifoinpacked_0.scala 27:17:@92528.4]
  wire  x748_fifoinpacked_0_io_active_0_in; // @[m_x748_fifoinpacked_0.scala 27:17:@92528.4]
  wire  x748_fifoinpacked_0_io_active_0_out; // @[m_x748_fifoinpacked_0.scala 27:17:@92528.4]
  wire  x749_fifooutraw_0_clock; // @[m_x749_fifooutraw_0.scala 27:17:@92552.4]
  wire  x749_fifooutraw_0_reset; // @[m_x749_fifooutraw_0.scala 27:17:@92552.4]
  wire  x752_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire  x752_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire  x752_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire  x752_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire [12:0] x752_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire [12:0] x752_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire  x752_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire  x752_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire  x752_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@92576.4]
  wire  x794_inr_Foreach_sm_clock; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_reset; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_enable; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_done; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_doneLatch; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_ctrDone; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_datapathEn; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_ctrInc; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_ctrRst; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_parentAck; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_backpressure; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  x794_inr_Foreach_sm_io_break; // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@92664.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@92664.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@92664.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@92664.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@92664.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@92710.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@92710.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@92710.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@92710.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@92710.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@92718.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@92718.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@92718.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@92718.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@92718.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_clock; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_reset; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_wPort_0_en_0; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_full; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_active_0_in; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_active_0_out; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire [31:0] x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire [31:0] x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_rr; // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
  wire  x1157_outr_UnitPipe_sm_clock; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_reset; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_enable; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_done; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_rst; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_ctrDone; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_ctrInc; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_parentAck; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  x1157_outr_UnitPipe_sm_io_childAck_0; // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@92942.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@92942.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@92942.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@92942.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@92942.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@92950.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@92950.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@92950.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@92950.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@92950.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_clock; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_reset; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TVALID; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TREADY; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire [255:0] x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TDATA; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TVALID; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TREADY; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire [255:0] x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TDATA; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire [7:0] x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TID; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire [7:0] x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TDEST; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_rr; // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
  wire  _T_254; // @[package.scala 96:25:@92669.4 package.scala 96:25:@92670.4]
  wire  _T_260; // @[implicits.scala 47:10:@92673.4]
  wire  _T_261; // @[sm_x1158_outr_UnitPipe.scala 70:41:@92674.4]
  wire  _T_262; // @[sm_x1158_outr_UnitPipe.scala 70:78:@92675.4]
  wire  _T_263; // @[sm_x1158_outr_UnitPipe.scala 70:76:@92676.4]
  wire  _T_275; // @[package.scala 96:25:@92715.4 package.scala 96:25:@92716.4]
  wire  _T_281; // @[package.scala 96:25:@92723.4 package.scala 96:25:@92724.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@92726.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@92735.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@92736.4]
  wire  _T_354; // @[package.scala 100:49:@92913.4]
  reg  _T_357; // @[package.scala 48:56:@92914.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@92947.4 package.scala 96:25:@92948.4]
  wire  _T_377; // @[package.scala 96:25:@92955.4 package.scala 96:25:@92956.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@92958.4]
  x747_fifoinraw_0 x747_fifoinraw_0 ( // @[m_x747_fifoinraw_0.scala 27:17:@92504.4]
    .clock(x747_fifoinraw_0_clock),
    .reset(x747_fifoinraw_0_reset)
  );
  x748_fifoinpacked_0 x748_fifoinpacked_0 ( // @[m_x748_fifoinpacked_0.scala 27:17:@92528.4]
    .clock(x748_fifoinpacked_0_clock),
    .reset(x748_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x748_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x748_fifoinpacked_0_io_full),
    .io_active_0_in(x748_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x748_fifoinpacked_0_io_active_0_out)
  );
  x747_fifoinraw_0 x749_fifooutraw_0 ( // @[m_x749_fifooutraw_0.scala 27:17:@92552.4]
    .clock(x749_fifooutraw_0_clock),
    .reset(x749_fifooutraw_0_reset)
  );
  x752_ctrchain x752_ctrchain ( // @[SpatialBlocks.scala 37:22:@92576.4]
    .clock(x752_ctrchain_clock),
    .reset(x752_ctrchain_reset),
    .io_input_reset(x752_ctrchain_io_input_reset),
    .io_input_enable(x752_ctrchain_io_input_enable),
    .io_output_counts_1(x752_ctrchain_io_output_counts_1),
    .io_output_counts_0(x752_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x752_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x752_ctrchain_io_output_oobs_1),
    .io_output_done(x752_ctrchain_io_output_done)
  );
  x794_inr_Foreach_sm x794_inr_Foreach_sm ( // @[sm_x794_inr_Foreach.scala 32:18:@92636.4]
    .clock(x794_inr_Foreach_sm_clock),
    .reset(x794_inr_Foreach_sm_reset),
    .io_enable(x794_inr_Foreach_sm_io_enable),
    .io_done(x794_inr_Foreach_sm_io_done),
    .io_doneLatch(x794_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x794_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x794_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x794_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x794_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x794_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x794_inr_Foreach_sm_io_backpressure),
    .io_break(x794_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@92664.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@92710.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@92718.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x794_inr_Foreach_kernelx794_inr_Foreach_concrete1 x794_inr_Foreach_kernelx794_inr_Foreach_concrete1 ( // @[sm_x794_inr_Foreach.scala 178:24:@92753.4]
    .clock(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_clock),
    .reset(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_reset),
    .io_in_x748_fifoinpacked_0_wPort_0_en_0(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_wPort_0_en_0),
    .io_in_x748_fifoinpacked_0_full(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_full),
    .io_in_x748_fifoinpacked_0_active_0_in(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_active_0_in),
    .io_in_x748_fifoinpacked_0_active_0_out(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x1157_outr_UnitPipe_sm ( // @[sm_x1157_outr_UnitPipe.scala 32:18:@92885.4]
    .clock(x1157_outr_UnitPipe_sm_clock),
    .reset(x1157_outr_UnitPipe_sm_reset),
    .io_enable(x1157_outr_UnitPipe_sm_io_enable),
    .io_done(x1157_outr_UnitPipe_sm_io_done),
    .io_rst(x1157_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x1157_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x1157_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x1157_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x1157_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x1157_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x1157_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@92942.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@92950.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1 x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1 ( // @[sm_x1157_outr_UnitPipe.scala 76:24:@92980.4]
    .clock(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_clock),
    .reset(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_reset),
    .io_in_x745_TVALID(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TVALID),
    .io_in_x745_TREADY(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TREADY),
    .io_in_x745_TDATA(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TDATA),
    .io_in_x744_TVALID(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TVALID),
    .io_in_x744_TREADY(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TREADY),
    .io_in_x744_TDATA(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TDATA),
    .io_in_x744_TID(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TID),
    .io_in_x744_TDEST(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TDEST),
    .io_sigsIn_smEnableOuts_0(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@92669.4 package.scala 96:25:@92670.4]
  assign _T_260 = x748_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@92673.4]
  assign _T_261 = ~ _T_260; // @[sm_x1158_outr_UnitPipe.scala 70:41:@92674.4]
  assign _T_262 = ~ x748_fifoinpacked_0_io_active_0_out; // @[sm_x1158_outr_UnitPipe.scala 70:78:@92675.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x1158_outr_UnitPipe.scala 70:76:@92676.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@92715.4 package.scala 96:25:@92716.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@92723.4 package.scala 96:25:@92724.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@92726.4]
  assign _T_286 = x794_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@92735.4]
  assign _T_287 = ~ x794_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@92736.4]
  assign _T_354 = x1157_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@92913.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@92947.4 package.scala 96:25:@92948.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@92955.4 package.scala 96:25:@92956.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@92958.4]
  assign io_in_x745_TVALID = x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TVALID; // @[sm_x1157_outr_UnitPipe.scala 48:23:@93037.4]
  assign io_in_x745_TDATA = x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TDATA; // @[sm_x1157_outr_UnitPipe.scala 48:23:@93035.4]
  assign io_in_x744_TREADY = x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TREADY; // @[sm_x1157_outr_UnitPipe.scala 49:23:@93045.4]
  assign io_sigsOut_smDoneIn_0 = x794_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@92733.4]
  assign io_sigsOut_smDoneIn_1 = x1157_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@92965.4]
  assign io_sigsOut_smCtrCopyDone_0 = x794_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@92752.4]
  assign io_sigsOut_smCtrCopyDone_1 = x1157_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@92979.4]
  assign x747_fifoinraw_0_clock = clock; // @[:@92505.4]
  assign x747_fifoinraw_0_reset = reset; // @[:@92506.4]
  assign x748_fifoinpacked_0_clock = clock; // @[:@92529.4]
  assign x748_fifoinpacked_0_reset = reset; // @[:@92530.4]
  assign x748_fifoinpacked_0_io_wPort_0_en_0 = x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@92813.4]
  assign x748_fifoinpacked_0_io_active_0_in = x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@92812.4]
  assign x749_fifooutraw_0_clock = clock; // @[:@92553.4]
  assign x749_fifooutraw_0_reset = reset; // @[:@92554.4]
  assign x752_ctrchain_clock = clock; // @[:@92577.4]
  assign x752_ctrchain_reset = reset; // @[:@92578.4]
  assign x752_ctrchain_io_input_reset = x794_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@92751.4]
  assign x752_ctrchain_io_input_enable = x794_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@92703.4 SpatialBlocks.scala 159:42:@92750.4]
  assign x794_inr_Foreach_sm_clock = clock; // @[:@92637.4]
  assign x794_inr_Foreach_sm_reset = reset; // @[:@92638.4]
  assign x794_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@92730.4]
  assign x794_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x1158_outr_UnitPipe.scala 69:38:@92672.4]
  assign x794_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@92732.4]
  assign x794_inr_Foreach_sm_io_backpressure = _T_263 | x794_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@92704.4]
  assign x794_inr_Foreach_sm_io_break = 1'h0; // @[sm_x1158_outr_UnitPipe.scala 73:36:@92682.4]
  assign RetimeWrapper_clock = clock; // @[:@92665.4]
  assign RetimeWrapper_reset = reset; // @[:@92666.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@92668.4]
  assign RetimeWrapper_io_in = x752_ctrchain_io_output_done; // @[package.scala 94:16:@92667.4]
  assign RetimeWrapper_1_clock = clock; // @[:@92711.4]
  assign RetimeWrapper_1_reset = reset; // @[:@92712.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@92714.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@92713.4]
  assign RetimeWrapper_2_clock = clock; // @[:@92719.4]
  assign RetimeWrapper_2_reset = reset; // @[:@92720.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@92722.4]
  assign RetimeWrapper_2_io_in = x794_inr_Foreach_sm_io_done; // @[package.scala 94:16:@92721.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_clock = clock; // @[:@92754.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_reset = reset; // @[:@92755.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_full = x748_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@92807.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_in_x748_fifoinpacked_0_active_0_out = x748_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@92806.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x794_inr_Foreach_sm_io_doneLatch; // @[sm_x794_inr_Foreach.scala 183:22:@92836.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x794_inr_Foreach.scala 183:22:@92834.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_break = x794_inr_Foreach_sm_io_break; // @[sm_x794_inr_Foreach.scala 183:22:@92832.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x752_ctrchain_io_output_counts_1[12]}},x752_ctrchain_io_output_counts_1}; // @[sm_x794_inr_Foreach.scala 183:22:@92827.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x752_ctrchain_io_output_counts_0[12]}},x752_ctrchain_io_output_counts_0}; // @[sm_x794_inr_Foreach.scala 183:22:@92826.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x752_ctrchain_io_output_oobs_0; // @[sm_x794_inr_Foreach.scala 183:22:@92824.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x752_ctrchain_io_output_oobs_1; // @[sm_x794_inr_Foreach.scala 183:22:@92825.4]
  assign x794_inr_Foreach_kernelx794_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x794_inr_Foreach.scala 182:18:@92820.4]
  assign x1157_outr_UnitPipe_sm_clock = clock; // @[:@92886.4]
  assign x1157_outr_UnitPipe_sm_reset = reset; // @[:@92887.4]
  assign x1157_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@92962.4]
  assign x1157_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@92937.4]
  assign x1157_outr_UnitPipe_sm_io_ctrDone = x1157_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x1158_outr_UnitPipe.scala 78:41:@92917.4]
  assign x1157_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@92964.4]
  assign x1157_outr_UnitPipe_sm_io_doneIn_0 = x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@92934.4]
  assign RetimeWrapper_3_clock = clock; // @[:@92943.4]
  assign RetimeWrapper_3_reset = reset; // @[:@92944.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@92946.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@92945.4]
  assign RetimeWrapper_4_clock = clock; // @[:@92951.4]
  assign RetimeWrapper_4_reset = reset; // @[:@92952.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@92954.4]
  assign RetimeWrapper_4_io_in = x1157_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@92953.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_clock = clock; // @[:@92981.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_reset = reset; // @[:@92982.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x745_TREADY = io_in_x745_TREADY; // @[sm_x1157_outr_UnitPipe.scala 48:23:@93036.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TVALID = io_in_x744_TVALID; // @[sm_x1157_outr_UnitPipe.scala 49:23:@93046.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TDATA = io_in_x744_TDATA; // @[sm_x1157_outr_UnitPipe.scala 49:23:@93044.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TID = io_in_x744_TID; // @[sm_x1157_outr_UnitPipe.scala 49:23:@93040.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_in_x744_TDEST = io_in_x744_TDEST; // @[sm_x1157_outr_UnitPipe.scala 49:23:@93039.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x1157_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x1157_outr_UnitPipe.scala 81:22:@93055.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x1157_outr_UnitPipe_sm_io_childAck_0; // @[sm_x1157_outr_UnitPipe.scala 81:22:@93053.4]
  assign x1157_outr_UnitPipe_kernelx1157_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x1157_outr_UnitPipe.scala 80:18:@93047.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x1180_outr_UnitPipe_sm( // @[:@93544.2]
  input   clock, // @[:@93545.4]
  input   reset, // @[:@93546.4]
  input   io_enable, // @[:@93547.4]
  output  io_done, // @[:@93547.4]
  input   io_parentAck, // @[:@93547.4]
  input   io_doneIn_0, // @[:@93547.4]
  input   io_doneIn_1, // @[:@93547.4]
  input   io_doneIn_2, // @[:@93547.4]
  output  io_enableOut_0, // @[:@93547.4]
  output  io_enableOut_1, // @[:@93547.4]
  output  io_enableOut_2, // @[:@93547.4]
  output  io_childAck_0, // @[:@93547.4]
  output  io_childAck_1, // @[:@93547.4]
  output  io_childAck_2, // @[:@93547.4]
  input   io_ctrCopyDone_0, // @[:@93547.4]
  input   io_ctrCopyDone_1, // @[:@93547.4]
  input   io_ctrCopyDone_2 // @[:@93547.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@93550.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@93550.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@93550.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@93550.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@93550.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@93550.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@93553.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@93553.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@93553.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@93553.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@93553.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@93553.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@93556.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@93556.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@93556.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@93556.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@93556.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@93556.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@93559.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@93559.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@93559.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@93559.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@93559.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@93559.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@93562.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@93562.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@93562.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@93562.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@93562.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@93562.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@93565.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@93565.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@93565.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@93565.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@93565.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@93565.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@93606.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@93606.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@93606.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@93606.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@93606.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@93606.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@93609.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@93609.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@93609.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@93609.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@93609.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@93609.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@93612.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@93612.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@93612.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@93612.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@93612.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@93612.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@93663.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@93663.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@93663.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@93663.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@93663.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@93677.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@93677.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@93677.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@93677.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@93677.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@93695.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@93695.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@93695.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@93695.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@93695.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@93732.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@93732.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@93732.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@93732.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@93732.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@93746.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@93746.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@93746.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@93746.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@93746.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@93764.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@93764.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@93764.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@93764.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@93764.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@93801.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@93801.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@93801.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@93801.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@93801.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@93815.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@93815.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@93815.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@93815.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@93815.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@93833.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@93833.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@93833.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@93833.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@93833.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@93890.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@93890.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@93890.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@93890.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@93890.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@93907.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@93907.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@93907.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@93907.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@93907.4]
  wire  _T_77; // @[Controllers.scala 80:47:@93568.4]
  wire  allDone; // @[Controllers.scala 80:47:@93569.4]
  wire  _T_151; // @[Controllers.scala 165:35:@93647.4]
  wire  _T_153; // @[Controllers.scala 165:60:@93648.4]
  wire  _T_154; // @[Controllers.scala 165:58:@93649.4]
  wire  _T_156; // @[Controllers.scala 165:76:@93650.4]
  wire  _T_157; // @[Controllers.scala 165:74:@93651.4]
  wire  _T_161; // @[Controllers.scala 165:109:@93654.4]
  wire  _T_164; // @[Controllers.scala 165:141:@93656.4]
  wire  _T_172; // @[package.scala 96:25:@93668.4 package.scala 96:25:@93669.4]
  wire  _T_176; // @[Controllers.scala 167:54:@93671.4]
  wire  _T_177; // @[Controllers.scala 167:52:@93672.4]
  wire  _T_184; // @[package.scala 96:25:@93682.4 package.scala 96:25:@93683.4]
  wire  _T_202; // @[package.scala 96:25:@93700.4 package.scala 96:25:@93701.4]
  wire  _T_206; // @[Controllers.scala 169:67:@93703.4]
  wire  _T_207; // @[Controllers.scala 169:86:@93704.4]
  wire  _T_219; // @[Controllers.scala 165:35:@93716.4]
  wire  _T_221; // @[Controllers.scala 165:60:@93717.4]
  wire  _T_222; // @[Controllers.scala 165:58:@93718.4]
  wire  _T_224; // @[Controllers.scala 165:76:@93719.4]
  wire  _T_225; // @[Controllers.scala 165:74:@93720.4]
  wire  _T_229; // @[Controllers.scala 165:109:@93723.4]
  wire  _T_232; // @[Controllers.scala 165:141:@93725.4]
  wire  _T_240; // @[package.scala 96:25:@93737.4 package.scala 96:25:@93738.4]
  wire  _T_244; // @[Controllers.scala 167:54:@93740.4]
  wire  _T_245; // @[Controllers.scala 167:52:@93741.4]
  wire  _T_252; // @[package.scala 96:25:@93751.4 package.scala 96:25:@93752.4]
  wire  _T_270; // @[package.scala 96:25:@93769.4 package.scala 96:25:@93770.4]
  wire  _T_274; // @[Controllers.scala 169:67:@93772.4]
  wire  _T_275; // @[Controllers.scala 169:86:@93773.4]
  wire  _T_287; // @[Controllers.scala 165:35:@93785.4]
  wire  _T_289; // @[Controllers.scala 165:60:@93786.4]
  wire  _T_290; // @[Controllers.scala 165:58:@93787.4]
  wire  _T_292; // @[Controllers.scala 165:76:@93788.4]
  wire  _T_293; // @[Controllers.scala 165:74:@93789.4]
  wire  _T_297; // @[Controllers.scala 165:109:@93792.4]
  wire  _T_300; // @[Controllers.scala 165:141:@93794.4]
  wire  _T_308; // @[package.scala 96:25:@93806.4 package.scala 96:25:@93807.4]
  wire  _T_312; // @[Controllers.scala 167:54:@93809.4]
  wire  _T_313; // @[Controllers.scala 167:52:@93810.4]
  wire  _T_320; // @[package.scala 96:25:@93820.4 package.scala 96:25:@93821.4]
  wire  _T_338; // @[package.scala 96:25:@93838.4 package.scala 96:25:@93839.4]
  wire  _T_342; // @[Controllers.scala 169:67:@93841.4]
  wire  _T_343; // @[Controllers.scala 169:86:@93842.4]
  wire  _T_358; // @[Controllers.scala 213:68:@93860.4]
  wire  _T_360; // @[Controllers.scala 213:90:@93862.4]
  wire  _T_362; // @[Controllers.scala 213:132:@93864.4]
  wire  _T_366; // @[Controllers.scala 213:68:@93869.4]
  wire  _T_368; // @[Controllers.scala 213:90:@93871.4]
  wire  _T_374; // @[Controllers.scala 213:68:@93877.4]
  wire  _T_376; // @[Controllers.scala 213:90:@93879.4]
  wire  _T_383; // @[package.scala 100:49:@93885.4]
  reg  _T_386; // @[package.scala 48:56:@93886.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@93888.4]
  reg  _T_400; // @[package.scala 48:56:@93904.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@93550.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@93553.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@93556.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@93559.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@93562.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@93565.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@93606.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@93609.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@93612.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@93663.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@93677.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@93695.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@93732.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@93746.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@93764.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@93801.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@93815.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@93833.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@93890.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@93907.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@93568.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@93569.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@93647.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@93648.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@93649.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@93650.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@93651.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@93654.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@93656.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@93668.4 package.scala 96:25:@93669.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@93671.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@93672.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@93682.4 package.scala 96:25:@93683.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@93700.4 package.scala 96:25:@93701.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@93703.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@93704.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@93716.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@93717.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@93718.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@93719.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@93720.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@93723.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@93725.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@93737.4 package.scala 96:25:@93738.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@93740.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@93741.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@93751.4 package.scala 96:25:@93752.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@93769.4 package.scala 96:25:@93770.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@93772.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@93773.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@93785.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@93786.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@93787.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@93788.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@93789.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@93792.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@93794.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@93806.4 package.scala 96:25:@93807.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@93809.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@93810.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@93820.4 package.scala 96:25:@93821.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@93838.4 package.scala 96:25:@93839.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@93841.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@93842.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@93860.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@93862.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@93864.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@93869.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@93871.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@93877.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@93879.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@93885.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@93888.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@93914.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@93868.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@93876.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@93884.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@93855.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@93857.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@93859.4]
  assign active_0_clock = clock; // @[:@93551.4]
  assign active_0_reset = reset; // @[:@93552.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@93658.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@93662.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@93572.4]
  assign active_1_clock = clock; // @[:@93554.4]
  assign active_1_reset = reset; // @[:@93555.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@93727.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@93731.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@93573.4]
  assign active_2_clock = clock; // @[:@93557.4]
  assign active_2_reset = reset; // @[:@93558.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@93796.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@93800.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@93574.4]
  assign done_0_clock = clock; // @[:@93560.4]
  assign done_0_reset = reset; // @[:@93561.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@93708.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@93586.4 Controllers.scala 170:32:@93715.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@93575.4]
  assign done_1_clock = clock; // @[:@93563.4]
  assign done_1_reset = reset; // @[:@93564.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@93777.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@93595.4 Controllers.scala 170:32:@93784.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@93576.4]
  assign done_2_clock = clock; // @[:@93566.4]
  assign done_2_reset = reset; // @[:@93567.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@93846.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@93604.4 Controllers.scala 170:32:@93853.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@93577.4]
  assign iterDone_0_clock = clock; // @[:@93607.4]
  assign iterDone_0_reset = reset; // @[:@93608.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@93676.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@93626.4 Controllers.scala 168:36:@93692.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@93615.4]
  assign iterDone_1_clock = clock; // @[:@93610.4]
  assign iterDone_1_reset = reset; // @[:@93611.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@93745.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@93635.4 Controllers.scala 168:36:@93761.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@93616.4]
  assign iterDone_2_clock = clock; // @[:@93613.4]
  assign iterDone_2_reset = reset; // @[:@93614.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@93814.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@93644.4 Controllers.scala 168:36:@93830.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@93617.4]
  assign RetimeWrapper_clock = clock; // @[:@93664.4]
  assign RetimeWrapper_reset = reset; // @[:@93665.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@93667.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@93666.4]
  assign RetimeWrapper_1_clock = clock; // @[:@93678.4]
  assign RetimeWrapper_1_reset = reset; // @[:@93679.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@93681.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@93680.4]
  assign RetimeWrapper_2_clock = clock; // @[:@93696.4]
  assign RetimeWrapper_2_reset = reset; // @[:@93697.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@93699.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@93698.4]
  assign RetimeWrapper_3_clock = clock; // @[:@93733.4]
  assign RetimeWrapper_3_reset = reset; // @[:@93734.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@93736.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@93735.4]
  assign RetimeWrapper_4_clock = clock; // @[:@93747.4]
  assign RetimeWrapper_4_reset = reset; // @[:@93748.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@93750.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@93749.4]
  assign RetimeWrapper_5_clock = clock; // @[:@93765.4]
  assign RetimeWrapper_5_reset = reset; // @[:@93766.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@93768.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@93767.4]
  assign RetimeWrapper_6_clock = clock; // @[:@93802.4]
  assign RetimeWrapper_6_reset = reset; // @[:@93803.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@93805.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@93804.4]
  assign RetimeWrapper_7_clock = clock; // @[:@93816.4]
  assign RetimeWrapper_7_reset = reset; // @[:@93817.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@93819.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@93818.4]
  assign RetimeWrapper_8_clock = clock; // @[:@93834.4]
  assign RetimeWrapper_8_reset = reset; // @[:@93835.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@93837.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@93836.4]
  assign RetimeWrapper_9_clock = clock; // @[:@93891.4]
  assign RetimeWrapper_9_reset = reset; // @[:@93892.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@93894.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@93893.4]
  assign RetimeWrapper_10_clock = clock; // @[:@93908.4]
  assign RetimeWrapper_10_reset = reset; // @[:@93909.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@93911.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@93910.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x1166_inr_UnitPipe_sm( // @[:@94087.2]
  input   clock, // @[:@94088.4]
  input   reset, // @[:@94089.4]
  input   io_enable, // @[:@94090.4]
  output  io_done, // @[:@94090.4]
  output  io_doneLatch, // @[:@94090.4]
  input   io_ctrDone, // @[:@94090.4]
  output  io_datapathEn, // @[:@94090.4]
  output  io_ctrInc, // @[:@94090.4]
  input   io_parentAck, // @[:@94090.4]
  input   io_backpressure // @[:@94090.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@94092.4]
  wire  active_reset; // @[Controllers.scala 261:22:@94092.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@94092.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@94092.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@94092.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@94092.4]
  wire  done_clock; // @[Controllers.scala 262:20:@94095.4]
  wire  done_reset; // @[Controllers.scala 262:20:@94095.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@94095.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@94095.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@94095.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@94095.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@94149.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@94149.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@94149.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@94149.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@94149.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@94157.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@94157.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@94157.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@94157.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@94157.4]
  wire  _T_80; // @[Controllers.scala 264:48:@94100.4]
  wire  _T_81; // @[Controllers.scala 264:46:@94101.4]
  wire  _T_82; // @[Controllers.scala 264:62:@94102.4]
  wire  _T_83; // @[Controllers.scala 264:60:@94103.4]
  wire  _T_100; // @[package.scala 100:49:@94120.4]
  reg  _T_103; // @[package.scala 48:56:@94121.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@94129.4]
  wire  _T_116; // @[Controllers.scala 283:41:@94137.4]
  wire  _T_117; // @[Controllers.scala 283:59:@94138.4]
  wire  _T_119; // @[Controllers.scala 284:37:@94141.4]
  reg  _T_125; // @[package.scala 48:56:@94145.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@94167.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@94170.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@94172.4]
  wire  _T_152; // @[Controllers.scala 292:61:@94173.4]
  wire  _T_153; // @[Controllers.scala 292:24:@94174.4]
  SRFF active ( // @[Controllers.scala 261:22:@94092.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@94095.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@94149.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@94157.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@94100.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@94101.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@94102.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@94103.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@94120.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@94129.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@94137.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@94138.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@94141.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@94172.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@94173.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@94174.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@94148.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@94176.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@94140.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@94143.4]
  assign active_clock = clock; // @[:@94093.4]
  assign active_reset = reset; // @[:@94094.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@94105.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@94109.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@94110.4]
  assign done_clock = clock; // @[:@94096.4]
  assign done_reset = reset; // @[:@94097.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@94125.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@94118.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@94119.4]
  assign RetimeWrapper_clock = clock; // @[:@94150.4]
  assign RetimeWrapper_reset = reset; // @[:@94151.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@94153.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@94152.4]
  assign RetimeWrapper_1_clock = clock; // @[:@94158.4]
  assign RetimeWrapper_1_reset = reset; // @[:@94159.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@94161.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@94160.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1( // @[:@94251.2]
  output        io_in_x1159_valid, // @[:@94254.4]
  output [63:0] io_in_x1159_bits_addr, // @[:@94254.4]
  output [31:0] io_in_x1159_bits_size, // @[:@94254.4]
  input  [63:0] io_in_x742_outdram_number, // @[:@94254.4]
  input         io_sigsIn_backpressure, // @[:@94254.4]
  input         io_sigsIn_datapathEn, // @[:@94254.4]
  input         io_rr // @[:@94254.4]
);
  wire [96:0] x1163_tuple; // @[Cat.scala 30:58:@94268.4]
  wire  _T_135; // @[implicits.scala 55:10:@94271.4]
  assign x1163_tuple = {33'h1fa400,io_in_x742_outdram_number}; // @[Cat.scala 30:58:@94268.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@94271.4]
  assign io_in_x1159_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x1166_inr_UnitPipe.scala 65:19:@94274.4]
  assign io_in_x1159_bits_addr = x1163_tuple[63:0]; // @[sm_x1166_inr_UnitPipe.scala 66:23:@94276.4]
  assign io_in_x1159_bits_size = x1163_tuple[95:64]; // @[sm_x1166_inr_UnitPipe.scala 67:23:@94278.4]
endmodule
module FF_13( // @[:@94280.2]
  input         clock, // @[:@94281.4]
  input         reset, // @[:@94282.4]
  output [22:0] io_rPort_0_output_0, // @[:@94283.4]
  input  [22:0] io_wPort_0_data_0, // @[:@94283.4]
  input         io_wPort_0_reset, // @[:@94283.4]
  input         io_wPort_0_en_0 // @[:@94283.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 311:19:@94298.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 315:32:@94300.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 315:12:@94301.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@94300.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 315:12:@94301.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@94303.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@94318.2]
  input         clock, // @[:@94319.4]
  input         reset, // @[:@94320.4]
  input         io_input_reset, // @[:@94321.4]
  input         io_input_enable, // @[:@94321.4]
  output [22:0] io_output_count_0, // @[:@94321.4]
  output        io_output_oobs_0, // @[:@94321.4]
  output        io_output_done // @[:@94321.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@94334.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@94334.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@94334.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@94334.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@94334.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@94334.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@94350.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@94350.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@94350.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@94350.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@94350.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@94350.4]
  wire  _T_36; // @[Counter.scala 264:45:@94353.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@94378.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@94379.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@94380.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@94381.4]
  wire  _T_57; // @[Counter.scala 293:18:@94383.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@94391.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@94394.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@94395.4]
  wire  _T_75; // @[Counter.scala 322:102:@94399.4]
  wire  _T_77; // @[Counter.scala 322:130:@94400.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@94334.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@94350.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@94353.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@94378.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@94379.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@94380.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@94381.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@94383.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@94391.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@94394.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@94395.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@94399.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@94400.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@94398.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@94402.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@94404.4]
  assign bases_0_clock = clock; // @[:@94335.4]
  assign bases_0_reset = reset; // @[:@94336.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@94397.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@94376.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@94377.4]
  assign SRFF_clock = clock; // @[:@94351.4]
  assign SRFF_reset = reset; // @[:@94352.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@94355.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@94357.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@94358.4]
endmodule
module x1168_ctrchain( // @[:@94409.2]
  input         clock, // @[:@94410.4]
  input         reset, // @[:@94411.4]
  input         io_input_reset, // @[:@94412.4]
  input         io_input_enable, // @[:@94412.4]
  output [22:0] io_output_counts_0, // @[:@94412.4]
  output        io_output_oobs_0, // @[:@94412.4]
  output        io_output_done // @[:@94412.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@94414.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@94414.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@94414.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@94414.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@94414.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@94414.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@94414.4]
  reg  wasDone; // @[Counter.scala 542:24:@94423.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@94429.4]
  wire  _T_47; // @[Counter.scala 546:80:@94430.4]
  reg  doneLatch; // @[Counter.scala 550:26:@94435.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@94436.4]
  wire  _T_55; // @[Counter.scala 551:19:@94437.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@94414.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@94429.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@94430.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@94436.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@94437.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@94439.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@94441.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@94432.4]
  assign ctrs_0_clock = clock; // @[:@94415.4]
  assign ctrs_0_reset = reset; // @[:@94416.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@94420.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@94421.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x1175_inr_Foreach_sm( // @[:@94629.2]
  input   clock, // @[:@94630.4]
  input   reset, // @[:@94631.4]
  input   io_enable, // @[:@94632.4]
  output  io_done, // @[:@94632.4]
  output  io_doneLatch, // @[:@94632.4]
  input   io_ctrDone, // @[:@94632.4]
  output  io_datapathEn, // @[:@94632.4]
  output  io_ctrInc, // @[:@94632.4]
  output  io_ctrRst, // @[:@94632.4]
  input   io_parentAck, // @[:@94632.4]
  input   io_backpressure, // @[:@94632.4]
  input   io_break // @[:@94632.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@94634.4]
  wire  active_reset; // @[Controllers.scala 261:22:@94634.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@94634.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@94634.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@94634.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@94634.4]
  wire  done_clock; // @[Controllers.scala 262:20:@94637.4]
  wire  done_reset; // @[Controllers.scala 262:20:@94637.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@94637.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@94637.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@94637.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@94637.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@94671.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@94671.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@94671.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@94671.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@94671.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@94693.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@94693.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@94693.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@94693.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@94693.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@94705.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@94705.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@94705.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@94705.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@94705.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@94713.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@94713.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@94713.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@94713.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@94713.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@94729.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@94729.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@94729.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@94729.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@94729.4]
  wire  _T_80; // @[Controllers.scala 264:48:@94642.4]
  wire  _T_81; // @[Controllers.scala 264:46:@94643.4]
  wire  _T_82; // @[Controllers.scala 264:62:@94644.4]
  wire  _T_83; // @[Controllers.scala 264:60:@94645.4]
  wire  _T_100; // @[package.scala 100:49:@94662.4]
  reg  _T_103; // @[package.scala 48:56:@94663.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@94676.4 package.scala 96:25:@94677.4]
  wire  _T_110; // @[package.scala 100:49:@94678.4]
  reg  _T_113; // @[package.scala 48:56:@94679.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@94681.4]
  wire  _T_118; // @[Controllers.scala 283:41:@94686.4]
  wire  _T_119; // @[Controllers.scala 283:59:@94687.4]
  wire  _T_121; // @[Controllers.scala 284:37:@94690.4]
  wire  _T_124; // @[package.scala 96:25:@94698.4 package.scala 96:25:@94699.4]
  wire  _T_126; // @[package.scala 100:49:@94700.4]
  reg  _T_129; // @[package.scala 48:56:@94701.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@94723.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@94725.4]
  reg  _T_153; // @[package.scala 48:56:@94726.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@94734.4 package.scala 96:25:@94735.4]
  wire  _T_158; // @[Controllers.scala 292:61:@94736.4]
  wire  _T_159; // @[Controllers.scala 292:24:@94737.4]
  SRFF active ( // @[Controllers.scala 261:22:@94634.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@94637.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@94671.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@94693.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@94705.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@94713.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@94729.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@94642.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@94643.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@94644.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@94645.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@94662.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@94676.4 package.scala 96:25:@94677.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@94678.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@94681.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@94686.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@94687.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@94690.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@94698.4 package.scala 96:25:@94699.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@94700.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@94725.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@94734.4 package.scala 96:25:@94735.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@94736.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@94737.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@94704.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@94739.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@94689.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@94692.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@94684.4]
  assign active_clock = clock; // @[:@94635.4]
  assign active_reset = reset; // @[:@94636.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@94647.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@94651.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@94652.4]
  assign done_clock = clock; // @[:@94638.4]
  assign done_reset = reset; // @[:@94639.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@94667.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@94660.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@94661.4]
  assign RetimeWrapper_clock = clock; // @[:@94672.4]
  assign RetimeWrapper_reset = reset; // @[:@94673.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@94675.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@94674.4]
  assign RetimeWrapper_1_clock = clock; // @[:@94694.4]
  assign RetimeWrapper_1_reset = reset; // @[:@94695.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@94697.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@94696.4]
  assign RetimeWrapper_2_clock = clock; // @[:@94706.4]
  assign RetimeWrapper_2_reset = reset; // @[:@94707.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@94709.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@94708.4]
  assign RetimeWrapper_3_clock = clock; // @[:@94714.4]
  assign RetimeWrapper_3_reset = reset; // @[:@94715.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@94717.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@94716.4]
  assign RetimeWrapper_4_clock = clock; // @[:@94730.4]
  assign RetimeWrapper_4_reset = reset; // @[:@94731.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@94733.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@94732.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1( // @[:@94951.2]
  input         clock, // @[:@94952.4]
  input         reset, // @[:@94953.4]
  output [20:0] io_in_x746_outbuf_0_rPort_0_ofs_0, // @[:@94954.4]
  output        io_in_x746_outbuf_0_rPort_0_en_0, // @[:@94954.4]
  output        io_in_x746_outbuf_0_rPort_0_backpressure, // @[:@94954.4]
  input  [7:0]  io_in_x746_outbuf_0_rPort_0_output_0, // @[:@94954.4]
  output        io_in_x1160_valid, // @[:@94954.4]
  output [7:0]  io_in_x1160_bits_wdata_0, // @[:@94954.4]
  output        io_in_x1160_bits_wstrb, // @[:@94954.4]
  input         io_sigsIn_backpressure, // @[:@94954.4]
  input         io_sigsIn_datapathEn, // @[:@94954.4]
  input         io_sigsIn_break, // @[:@94954.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@94954.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@94954.4]
  input         io_rr // @[:@94954.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@94981.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@94981.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@95010.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@95010.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@95010.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@95010.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@95010.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@95019.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@95019.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@95019.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@95019.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@95019.4]
  wire  b1170; // @[sm_x1175_inr_Foreach.scala 62:19:@94989.4]
  wire  _T_274; // @[sm_x1175_inr_Foreach.scala 67:134:@94993.4]
  wire  _T_278; // @[implicits.scala 55:10:@94996.4]
  wire  _T_279; // @[sm_x1175_inr_Foreach.scala 67:151:@94997.4]
  wire [8:0] x1173_tuple; // @[Cat.scala 30:58:@95007.4]
  wire  _T_290; // @[package.scala 96:25:@95024.4 package.scala 96:25:@95025.4]
  wire  _T_292; // @[implicits.scala 55:10:@95026.4]
  wire  x1382_b1170_D2; // @[package.scala 96:25:@95015.4 package.scala 96:25:@95016.4]
  wire  _T_293; // @[sm_x1175_inr_Foreach.scala 74:113:@95027.4]
  wire [31:0] b1169_number; // @[Math.scala 712:22:@94986.4 Math.scala 713:14:@94987.4]
  _ _ ( // @[Math.scala 709:24:@94981.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@95010.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@95019.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b1170 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x1175_inr_Foreach.scala 62:19:@94989.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x1175_inr_Foreach.scala 67:134:@94993.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@94996.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x1175_inr_Foreach.scala 67:151:@94997.4]
  assign x1173_tuple = {1'h1,io_in_x746_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@95007.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@95024.4 package.scala 96:25:@95025.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@95026.4]
  assign x1382_b1170_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@95015.4 package.scala 96:25:@95016.4]
  assign _T_293 = _T_292 & x1382_b1170_D2; // @[sm_x1175_inr_Foreach.scala 74:113:@95027.4]
  assign b1169_number = __io_result; // @[Math.scala 712:22:@94986.4 Math.scala 713:14:@94987.4]
  assign io_in_x746_outbuf_0_rPort_0_ofs_0 = b1169_number[20:0]; // @[MemInterfaceType.scala 107:54:@95000.4]
  assign io_in_x746_outbuf_0_rPort_0_en_0 = _T_279 & b1170; // @[MemInterfaceType.scala 110:79:@95002.4]
  assign io_in_x746_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@95001.4]
  assign io_in_x1160_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x1175_inr_Foreach.scala 74:19:@95029.4]
  assign io_in_x1160_bits_wdata_0 = x1173_tuple[7:0]; // @[sm_x1175_inr_Foreach.scala 75:27:@95031.4]
  assign io_in_x1160_bits_wstrb = x1173_tuple[8]; // @[sm_x1175_inr_Foreach.scala 76:24:@95033.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@94984.4]
  assign RetimeWrapper_clock = clock; // @[:@95011.4]
  assign RetimeWrapper_reset = reset; // @[:@95012.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@95014.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@95013.4]
  assign RetimeWrapper_1_clock = clock; // @[:@95020.4]
  assign RetimeWrapper_1_reset = reset; // @[:@95021.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@95023.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@95022.4]
endmodule
module x1179_inr_UnitPipe_sm( // @[:@95189.2]
  input   clock, // @[:@95190.4]
  input   reset, // @[:@95191.4]
  input   io_enable, // @[:@95192.4]
  output  io_done, // @[:@95192.4]
  output  io_doneLatch, // @[:@95192.4]
  input   io_ctrDone, // @[:@95192.4]
  output  io_datapathEn, // @[:@95192.4]
  output  io_ctrInc, // @[:@95192.4]
  input   io_parentAck // @[:@95192.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@95194.4]
  wire  active_reset; // @[Controllers.scala 261:22:@95194.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@95194.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@95194.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@95194.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@95194.4]
  wire  done_clock; // @[Controllers.scala 262:20:@95197.4]
  wire  done_reset; // @[Controllers.scala 262:20:@95197.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@95197.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@95197.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@95197.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@95197.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@95231.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@95231.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@95231.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@95231.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@95231.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@95253.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@95253.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@95253.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@95253.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@95253.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@95265.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@95265.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@95265.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@95265.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@95265.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@95273.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@95273.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@95273.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@95273.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@95273.4]
  wire  _T_80; // @[Controllers.scala 264:48:@95202.4]
  wire  _T_81; // @[Controllers.scala 264:46:@95203.4]
  wire  _T_82; // @[Controllers.scala 264:62:@95204.4]
  wire  _T_100; // @[package.scala 100:49:@95222.4]
  reg  _T_103; // @[package.scala 48:56:@95223.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@95246.4]
  wire  _T_124; // @[package.scala 96:25:@95258.4 package.scala 96:25:@95259.4]
  wire  _T_126; // @[package.scala 100:49:@95260.4]
  reg  _T_129; // @[package.scala 48:56:@95261.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@95283.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@95285.4]
  reg  _T_153; // @[package.scala 48:56:@95286.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@95288.4]
  wire  _T_156; // @[Controllers.scala 292:61:@95289.4]
  wire  _T_157; // @[Controllers.scala 292:24:@95290.4]
  SRFF active ( // @[Controllers.scala 261:22:@95194.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@95197.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@95231.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@95253.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@95265.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@95273.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@95202.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@95203.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@95204.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@95222.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@95246.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@95258.4 package.scala 96:25:@95259.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@95260.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@95285.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@95288.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@95289.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@95290.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@95264.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@95292.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@95249.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@95252.4]
  assign active_clock = clock; // @[:@95195.4]
  assign active_reset = reset; // @[:@95196.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@95207.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@95211.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@95212.4]
  assign done_clock = clock; // @[:@95198.4]
  assign done_reset = reset; // @[:@95199.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@95227.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@95220.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@95221.4]
  assign RetimeWrapper_clock = clock; // @[:@95232.4]
  assign RetimeWrapper_reset = reset; // @[:@95233.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@95235.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@95234.4]
  assign RetimeWrapper_1_clock = clock; // @[:@95254.4]
  assign RetimeWrapper_1_reset = reset; // @[:@95255.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@95257.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@95256.4]
  assign RetimeWrapper_2_clock = clock; // @[:@95266.4]
  assign RetimeWrapper_2_reset = reset; // @[:@95267.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@95269.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@95268.4]
  assign RetimeWrapper_3_clock = clock; // @[:@95274.4]
  assign RetimeWrapper_3_reset = reset; // @[:@95275.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@95277.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@95276.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1( // @[:@95367.2]
  output  io_in_x1161_ready, // @[:@95370.4]
  input   io_sigsIn_datapathEn // @[:@95370.4]
);
  assign io_in_x1161_ready = io_sigsIn_datapathEn; // @[sm_x1179_inr_UnitPipe.scala 57:19:@95382.4]
endmodule
module x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1( // @[:@95385.2]
  input         clock, // @[:@95386.4]
  input         reset, // @[:@95387.4]
  output [20:0] io_in_x746_outbuf_0_rPort_0_ofs_0, // @[:@95388.4]
  output        io_in_x746_outbuf_0_rPort_0_en_0, // @[:@95388.4]
  output        io_in_x746_outbuf_0_rPort_0_backpressure, // @[:@95388.4]
  input  [7:0]  io_in_x746_outbuf_0_rPort_0_output_0, // @[:@95388.4]
  input         io_in_x1159_ready, // @[:@95388.4]
  output        io_in_x1159_valid, // @[:@95388.4]
  output [63:0] io_in_x1159_bits_addr, // @[:@95388.4]
  output [31:0] io_in_x1159_bits_size, // @[:@95388.4]
  input  [63:0] io_in_x742_outdram_number, // @[:@95388.4]
  input         io_in_x1160_ready, // @[:@95388.4]
  output        io_in_x1160_valid, // @[:@95388.4]
  output [7:0]  io_in_x1160_bits_wdata_0, // @[:@95388.4]
  output        io_in_x1160_bits_wstrb, // @[:@95388.4]
  output        io_in_x1161_ready, // @[:@95388.4]
  input         io_in_x1161_valid, // @[:@95388.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@95388.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@95388.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@95388.4]
  input         io_sigsIn_smChildAcks_0, // @[:@95388.4]
  input         io_sigsIn_smChildAcks_1, // @[:@95388.4]
  input         io_sigsIn_smChildAcks_2, // @[:@95388.4]
  output        io_sigsOut_smDoneIn_0, // @[:@95388.4]
  output        io_sigsOut_smDoneIn_1, // @[:@95388.4]
  output        io_sigsOut_smDoneIn_2, // @[:@95388.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@95388.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@95388.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@95388.4]
  input         io_rr // @[:@95388.4]
);
  wire  x1166_inr_UnitPipe_sm_clock; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_reset; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_enable; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_done; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_doneLatch; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_ctrDone; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_datapathEn; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_ctrInc; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_parentAck; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  x1166_inr_UnitPipe_sm_io_backpressure; // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@95512.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@95512.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@95512.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@95512.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@95512.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@95520.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@95520.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@95520.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@95520.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@95520.4]
  wire  x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_valid; // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
  wire [63:0] x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_bits_addr; // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
  wire [31:0] x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_bits_size; // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
  wire [63:0] x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x742_outdram_number; // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
  wire  x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
  wire  x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
  wire  x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_rr; // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
  wire  x1168_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@95618.4]
  wire  x1168_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@95618.4]
  wire  x1168_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@95618.4]
  wire  x1168_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@95618.4]
  wire [22:0] x1168_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@95618.4]
  wire  x1168_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@95618.4]
  wire  x1168_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@95618.4]
  wire  x1175_inr_Foreach_sm_clock; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_reset; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_enable; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_done; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_doneLatch; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_ctrDone; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_datapathEn; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_ctrInc; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_ctrRst; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_parentAck; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_backpressure; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  x1175_inr_Foreach_sm_io_break; // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@95699.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@95699.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@95699.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@95699.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@95699.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@95739.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@95739.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@95739.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@95739.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@95739.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@95747.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@95747.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@95747.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@95747.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@95747.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_clock; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_reset; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire [20:0] x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_en_0; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire [7:0] x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_output_0; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_valid; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire [7:0] x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_bits_wdata_0; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_bits_wstrb; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire [31:0] x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_rr; // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
  wire  x1179_inr_UnitPipe_sm_clock; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_reset; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_io_enable; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_io_done; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_io_doneLatch; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_io_ctrDone; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_io_datapathEn; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_io_ctrInc; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  x1179_inr_UnitPipe_sm_io_parentAck; // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@95959.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@95959.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@95959.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@95959.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@95959.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@95967.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@95967.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@95967.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@95967.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@95967.4]
  wire  x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1_io_in_x1161_ready; // @[sm_x1179_inr_UnitPipe.scala 60:24:@95997.4]
  wire  x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x1179_inr_UnitPipe.scala 60:24:@95997.4]
  wire  _T_359; // @[package.scala 100:49:@95483.4]
  reg  _T_362; // @[package.scala 48:56:@95484.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@95517.4 package.scala 96:25:@95518.4]
  wire  _T_381; // @[package.scala 96:25:@95525.4 package.scala 96:25:@95526.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@95528.4]
  wire  _T_454; // @[package.scala 96:25:@95704.4 package.scala 96:25:@95705.4]
  wire  _T_468; // @[package.scala 96:25:@95744.4 package.scala 96:25:@95745.4]
  wire  _T_474; // @[package.scala 96:25:@95752.4 package.scala 96:25:@95753.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@95755.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@95764.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@95765.4]
  wire  _T_547; // @[package.scala 100:49:@95930.4]
  reg  _T_550; // @[package.scala 48:56:@95931.4]
  reg [31:0] _RAND_1;
  wire  x1179_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x1180_outr_UnitPipe.scala 101:57:@95937.4]
  wire  _T_563; // @[package.scala 96:25:@95964.4 package.scala 96:25:@95965.4]
  wire  _T_569; // @[package.scala 96:25:@95972.4 package.scala 96:25:@95973.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@95975.4]
  wire  x1179_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@95976.4]
  x1166_inr_UnitPipe_sm x1166_inr_UnitPipe_sm ( // @[sm_x1166_inr_UnitPipe.scala 33:18:@95455.4]
    .clock(x1166_inr_UnitPipe_sm_clock),
    .reset(x1166_inr_UnitPipe_sm_reset),
    .io_enable(x1166_inr_UnitPipe_sm_io_enable),
    .io_done(x1166_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x1166_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x1166_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x1166_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x1166_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x1166_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x1166_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@95512.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@95520.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1 x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1 ( // @[sm_x1166_inr_UnitPipe.scala 69:24:@95550.4]
    .io_in_x1159_valid(x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_valid),
    .io_in_x1159_bits_addr(x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_bits_addr),
    .io_in_x1159_bits_size(x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_bits_size),
    .io_in_x742_outdram_number(x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x742_outdram_number),
    .io_sigsIn_backpressure(x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_rr)
  );
  x1168_ctrchain x1168_ctrchain ( // @[SpatialBlocks.scala 37:22:@95618.4]
    .clock(x1168_ctrchain_clock),
    .reset(x1168_ctrchain_reset),
    .io_input_reset(x1168_ctrchain_io_input_reset),
    .io_input_enable(x1168_ctrchain_io_input_enable),
    .io_output_counts_0(x1168_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x1168_ctrchain_io_output_oobs_0),
    .io_output_done(x1168_ctrchain_io_output_done)
  );
  x1175_inr_Foreach_sm x1175_inr_Foreach_sm ( // @[sm_x1175_inr_Foreach.scala 33:18:@95671.4]
    .clock(x1175_inr_Foreach_sm_clock),
    .reset(x1175_inr_Foreach_sm_reset),
    .io_enable(x1175_inr_Foreach_sm_io_enable),
    .io_done(x1175_inr_Foreach_sm_io_done),
    .io_doneLatch(x1175_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x1175_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x1175_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x1175_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x1175_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x1175_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x1175_inr_Foreach_sm_io_backpressure),
    .io_break(x1175_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@95699.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@95739.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@95747.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1 x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1 ( // @[sm_x1175_inr_Foreach.scala 78:24:@95782.4]
    .clock(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_clock),
    .reset(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_reset),
    .io_in_x746_outbuf_0_rPort_0_ofs_0(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0),
    .io_in_x746_outbuf_0_rPort_0_en_0(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_en_0),
    .io_in_x746_outbuf_0_rPort_0_backpressure(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure),
    .io_in_x746_outbuf_0_rPort_0_output_0(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_output_0),
    .io_in_x1160_valid(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_valid),
    .io_in_x1160_bits_wdata_0(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_bits_wdata_0),
    .io_in_x1160_bits_wstrb(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_bits_wstrb),
    .io_sigsIn_backpressure(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_rr)
  );
  x1179_inr_UnitPipe_sm x1179_inr_UnitPipe_sm ( // @[sm_x1179_inr_UnitPipe.scala 32:18:@95902.4]
    .clock(x1179_inr_UnitPipe_sm_clock),
    .reset(x1179_inr_UnitPipe_sm_reset),
    .io_enable(x1179_inr_UnitPipe_sm_io_enable),
    .io_done(x1179_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x1179_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x1179_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x1179_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x1179_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x1179_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@95959.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@95967.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1 x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1 ( // @[sm_x1179_inr_UnitPipe.scala 60:24:@95997.4]
    .io_in_x1161_ready(x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1_io_in_x1161_ready),
    .io_sigsIn_datapathEn(x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x1166_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@95483.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@95517.4 package.scala 96:25:@95518.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@95525.4 package.scala 96:25:@95526.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@95528.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@95704.4 package.scala 96:25:@95705.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@95744.4 package.scala 96:25:@95745.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@95752.4 package.scala 96:25:@95753.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@95755.4]
  assign _T_479 = x1175_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@95764.4]
  assign _T_480 = ~ x1175_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@95765.4]
  assign _T_547 = x1179_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@95930.4]
  assign x1179_inr_UnitPipe_sigsIn_forwardpressure = io_in_x1161_valid | x1179_inr_UnitPipe_sm_io_doneLatch; // @[sm_x1180_outr_UnitPipe.scala 101:57:@95937.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@95964.4 package.scala 96:25:@95965.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@95972.4 package.scala 96:25:@95973.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@95975.4]
  assign x1179_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@95976.4]
  assign io_in_x746_outbuf_0_rPort_0_ofs_0 = x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@95833.4]
  assign io_in_x746_outbuf_0_rPort_0_en_0 = x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@95832.4]
  assign io_in_x746_outbuf_0_rPort_0_backpressure = x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@95831.4]
  assign io_in_x1159_valid = x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_valid; // @[sm_x1166_inr_UnitPipe.scala 49:24:@95588.4]
  assign io_in_x1159_bits_addr = x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_bits_addr; // @[sm_x1166_inr_UnitPipe.scala 49:24:@95587.4]
  assign io_in_x1159_bits_size = x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x1159_bits_size; // @[sm_x1166_inr_UnitPipe.scala 49:24:@95586.4]
  assign io_in_x1160_valid = x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_valid; // @[sm_x1175_inr_Foreach.scala 50:24:@95837.4]
  assign io_in_x1160_bits_wdata_0 = x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_bits_wdata_0; // @[sm_x1175_inr_Foreach.scala 50:24:@95836.4]
  assign io_in_x1160_bits_wstrb = x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x1160_bits_wstrb; // @[sm_x1175_inr_Foreach.scala 50:24:@95835.4]
  assign io_in_x1161_ready = x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1_io_in_x1161_ready; // @[sm_x1179_inr_UnitPipe.scala 46:24:@96033.4]
  assign io_sigsOut_smDoneIn_0 = x1166_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@95535.4]
  assign io_sigsOut_smDoneIn_1 = x1175_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@95762.4]
  assign io_sigsOut_smDoneIn_2 = x1179_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@95982.4]
  assign io_sigsOut_smCtrCopyDone_0 = x1166_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@95549.4]
  assign io_sigsOut_smCtrCopyDone_1 = x1175_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@95781.4]
  assign io_sigsOut_smCtrCopyDone_2 = x1179_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@95996.4]
  assign x1166_inr_UnitPipe_sm_clock = clock; // @[:@95456.4]
  assign x1166_inr_UnitPipe_sm_reset = reset; // @[:@95457.4]
  assign x1166_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@95532.4]
  assign x1166_inr_UnitPipe_sm_io_ctrDone = x1166_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x1180_outr_UnitPipe.scala 77:40:@95487.4]
  assign x1166_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@95534.4]
  assign x1166_inr_UnitPipe_sm_io_backpressure = io_in_x1159_ready | x1166_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@95506.4]
  assign RetimeWrapper_clock = clock; // @[:@95513.4]
  assign RetimeWrapper_reset = reset; // @[:@95514.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@95516.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@95515.4]
  assign RetimeWrapper_1_clock = clock; // @[:@95521.4]
  assign RetimeWrapper_1_reset = reset; // @[:@95522.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@95524.4]
  assign RetimeWrapper_1_io_in = x1166_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@95523.4]
  assign x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_in_x742_outdram_number = io_in_x742_outdram_number; // @[sm_x1166_inr_UnitPipe.scala 50:31:@95590.4]
  assign x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x1159_ready | x1166_inr_UnitPipe_sm_io_doneLatch; // @[sm_x1166_inr_UnitPipe.scala 74:22:@95605.4]
  assign x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x1166_inr_UnitPipe_sm_io_datapathEn; // @[sm_x1166_inr_UnitPipe.scala 74:22:@95603.4]
  assign x1166_inr_UnitPipe_kernelx1166_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x1166_inr_UnitPipe.scala 73:18:@95591.4]
  assign x1168_ctrchain_clock = clock; // @[:@95619.4]
  assign x1168_ctrchain_reset = reset; // @[:@95620.4]
  assign x1168_ctrchain_io_input_reset = x1175_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@95780.4]
  assign x1168_ctrchain_io_input_enable = x1175_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@95732.4 SpatialBlocks.scala 159:42:@95779.4]
  assign x1175_inr_Foreach_sm_clock = clock; // @[:@95672.4]
  assign x1175_inr_Foreach_sm_reset = reset; // @[:@95673.4]
  assign x1175_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@95759.4]
  assign x1175_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x1180_outr_UnitPipe.scala 90:39:@95707.4]
  assign x1175_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@95761.4]
  assign x1175_inr_Foreach_sm_io_backpressure = io_in_x1160_ready | x1175_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@95733.4]
  assign x1175_inr_Foreach_sm_io_break = 1'h0; // @[sm_x1180_outr_UnitPipe.scala 94:37:@95713.4]
  assign RetimeWrapper_2_clock = clock; // @[:@95700.4]
  assign RetimeWrapper_2_reset = reset; // @[:@95701.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@95703.4]
  assign RetimeWrapper_2_io_in = x1168_ctrchain_io_output_done; // @[package.scala 94:16:@95702.4]
  assign RetimeWrapper_3_clock = clock; // @[:@95740.4]
  assign RetimeWrapper_3_reset = reset; // @[:@95741.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@95743.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@95742.4]
  assign RetimeWrapper_4_clock = clock; // @[:@95748.4]
  assign RetimeWrapper_4_reset = reset; // @[:@95749.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@95751.4]
  assign RetimeWrapper_4_io_in = x1175_inr_Foreach_sm_io_done; // @[package.scala 94:16:@95750.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_clock = clock; // @[:@95783.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_reset = reset; // @[:@95784.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_in_x746_outbuf_0_rPort_0_output_0 = io_in_x746_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@95830.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x1160_ready | x1175_inr_Foreach_sm_io_doneLatch; // @[sm_x1175_inr_Foreach.scala 83:22:@95853.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x1175_inr_Foreach.scala 83:22:@95851.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_break = x1175_inr_Foreach_sm_io_break; // @[sm_x1175_inr_Foreach.scala 83:22:@95849.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x1168_ctrchain_io_output_counts_0[22]}},x1168_ctrchain_io_output_counts_0}; // @[sm_x1175_inr_Foreach.scala 83:22:@95844.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x1168_ctrchain_io_output_oobs_0; // @[sm_x1175_inr_Foreach.scala 83:22:@95843.4]
  assign x1175_inr_Foreach_kernelx1175_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x1175_inr_Foreach.scala 82:18:@95839.4]
  assign x1179_inr_UnitPipe_sm_clock = clock; // @[:@95903.4]
  assign x1179_inr_UnitPipe_sm_reset = reset; // @[:@95904.4]
  assign x1179_inr_UnitPipe_sm_io_enable = x1179_inr_UnitPipe_sigsIn_baseEn & x1179_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@95979.4]
  assign x1179_inr_UnitPipe_sm_io_ctrDone = x1179_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x1180_outr_UnitPipe.scala 99:40:@95934.4]
  assign x1179_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@95981.4]
  assign RetimeWrapper_5_clock = clock; // @[:@95960.4]
  assign RetimeWrapper_5_reset = reset; // @[:@95961.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@95963.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@95962.4]
  assign RetimeWrapper_6_clock = clock; // @[:@95968.4]
  assign RetimeWrapper_6_reset = reset; // @[:@95969.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@95971.4]
  assign RetimeWrapper_6_io_in = x1179_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@95970.4]
  assign x1179_inr_UnitPipe_kernelx1179_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x1179_inr_UnitPipe_sm_io_datapathEn; // @[sm_x1179_inr_UnitPipe.scala 65:22:@96046.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x1251_kernelx1251_concrete1( // @[:@96062.2]
  input          clock, // @[:@96063.4]
  input          reset, // @[:@96064.4]
  output [20:0]  io_in_x746_outbuf_0_rPort_0_ofs_0, // @[:@96065.4]
  output         io_in_x746_outbuf_0_rPort_0_en_0, // @[:@96065.4]
  output         io_in_x746_outbuf_0_rPort_0_backpressure, // @[:@96065.4]
  input  [7:0]   io_in_x746_outbuf_0_rPort_0_output_0, // @[:@96065.4]
  input          io_in_x1159_ready, // @[:@96065.4]
  output         io_in_x1159_valid, // @[:@96065.4]
  output [63:0]  io_in_x1159_bits_addr, // @[:@96065.4]
  output [31:0]  io_in_x1159_bits_size, // @[:@96065.4]
  input  [63:0]  io_in_x742_outdram_number, // @[:@96065.4]
  input          io_in_x1160_ready, // @[:@96065.4]
  output         io_in_x1160_valid, // @[:@96065.4]
  output [7:0]   io_in_x1160_bits_wdata_0, // @[:@96065.4]
  output         io_in_x1160_bits_wstrb, // @[:@96065.4]
  output         io_in_x745_TVALID, // @[:@96065.4]
  input          io_in_x745_TREADY, // @[:@96065.4]
  output [255:0] io_in_x745_TDATA, // @[:@96065.4]
  input          io_in_x744_TVALID, // @[:@96065.4]
  output         io_in_x744_TREADY, // @[:@96065.4]
  input  [255:0] io_in_x744_TDATA, // @[:@96065.4]
  input  [7:0]   io_in_x744_TID, // @[:@96065.4]
  input  [7:0]   io_in_x744_TDEST, // @[:@96065.4]
  output         io_in_x1161_ready, // @[:@96065.4]
  input          io_in_x1161_valid, // @[:@96065.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@96065.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@96065.4]
  input          io_sigsIn_smChildAcks_0, // @[:@96065.4]
  input          io_sigsIn_smChildAcks_1, // @[:@96065.4]
  output         io_sigsOut_smDoneIn_0, // @[:@96065.4]
  output         io_sigsOut_smDoneIn_1, // @[:@96065.4]
  input          io_rr // @[:@96065.4]
);
  wire  x1158_outr_UnitPipe_sm_clock; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_reset; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_enable; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_done; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_parentAck; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_childAck_0; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_childAck_1; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  x1158_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@96200.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@96200.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@96200.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@96200.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@96200.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@96208.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@96208.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@96208.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@96208.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@96208.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_clock; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_reset; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TVALID; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TREADY; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire [255:0] x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TDATA; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TVALID; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TREADY; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire [255:0] x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TDATA; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire [7:0] x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TID; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire [7:0] x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TDEST; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_rr; // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
  wire  x1180_outr_UnitPipe_sm_clock; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_reset; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_enable; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_done; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_parentAck; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_childAck_0; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_childAck_1; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_childAck_2; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  x1180_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@96489.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@96489.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@96489.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@96489.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@96489.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@96497.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@96497.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@96497.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@96497.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@96497.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_clock; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_reset; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire [20:0] x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_en_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire [7:0] x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_output_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_ready; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_valid; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire [63:0] x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_bits_addr; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire [31:0] x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_bits_size; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire [63:0] x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x742_outdram_number; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_ready; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_valid; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire [7:0] x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_bits_wdata_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_bits_wstrb; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1161_ready; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1161_valid; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_rr; // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
  wire  _T_408; // @[package.scala 96:25:@96205.4 package.scala 96:25:@96206.4]
  wire  _T_414; // @[package.scala 96:25:@96213.4 package.scala 96:25:@96214.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@96216.4]
  wire  _T_508; // @[package.scala 96:25:@96494.4 package.scala 96:25:@96495.4]
  wire  _T_514; // @[package.scala 96:25:@96502.4 package.scala 96:25:@96503.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@96505.4]
  x1158_outr_UnitPipe_sm x1158_outr_UnitPipe_sm ( // @[sm_x1158_outr_UnitPipe.scala 32:18:@96138.4]
    .clock(x1158_outr_UnitPipe_sm_clock),
    .reset(x1158_outr_UnitPipe_sm_reset),
    .io_enable(x1158_outr_UnitPipe_sm_io_enable),
    .io_done(x1158_outr_UnitPipe_sm_io_done),
    .io_parentAck(x1158_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x1158_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x1158_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x1158_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x1158_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x1158_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x1158_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x1158_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x1158_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@96200.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@96208.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1 x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1 ( // @[sm_x1158_outr_UnitPipe.scala 87:24:@96239.4]
    .clock(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_clock),
    .reset(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_reset),
    .io_in_x745_TVALID(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TVALID),
    .io_in_x745_TREADY(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TREADY),
    .io_in_x745_TDATA(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TDATA),
    .io_in_x744_TVALID(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TVALID),
    .io_in_x744_TREADY(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TREADY),
    .io_in_x744_TDATA(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TDATA),
    .io_in_x744_TID(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TID),
    .io_in_x744_TDEST(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TDEST),
    .io_sigsIn_smEnableOuts_0(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_rr)
  );
  x1180_outr_UnitPipe_sm x1180_outr_UnitPipe_sm ( // @[sm_x1180_outr_UnitPipe.scala 36:18:@96417.4]
    .clock(x1180_outr_UnitPipe_sm_clock),
    .reset(x1180_outr_UnitPipe_sm_reset),
    .io_enable(x1180_outr_UnitPipe_sm_io_enable),
    .io_done(x1180_outr_UnitPipe_sm_io_done),
    .io_parentAck(x1180_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x1180_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x1180_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x1180_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x1180_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x1180_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x1180_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x1180_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x1180_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x1180_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x1180_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x1180_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x1180_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@96489.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@96497.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1 x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1 ( // @[sm_x1180_outr_UnitPipe.scala 108:24:@96529.4]
    .clock(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_clock),
    .reset(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_reset),
    .io_in_x746_outbuf_0_rPort_0_ofs_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0),
    .io_in_x746_outbuf_0_rPort_0_en_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_en_0),
    .io_in_x746_outbuf_0_rPort_0_backpressure(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure),
    .io_in_x746_outbuf_0_rPort_0_output_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_output_0),
    .io_in_x1159_ready(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_ready),
    .io_in_x1159_valid(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_valid),
    .io_in_x1159_bits_addr(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_bits_addr),
    .io_in_x1159_bits_size(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_bits_size),
    .io_in_x742_outdram_number(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x742_outdram_number),
    .io_in_x1160_ready(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_ready),
    .io_in_x1160_valid(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_valid),
    .io_in_x1160_bits_wdata_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_bits_wdata_0),
    .io_in_x1160_bits_wstrb(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_bits_wstrb),
    .io_in_x1161_ready(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1161_ready),
    .io_in_x1161_valid(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1161_valid),
    .io_sigsIn_smEnableOuts_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@96205.4 package.scala 96:25:@96206.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@96213.4 package.scala 96:25:@96214.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@96216.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@96494.4 package.scala 96:25:@96495.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@96502.4 package.scala 96:25:@96503.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@96505.4]
  assign io_in_x746_outbuf_0_rPort_0_ofs_0 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@96612.4]
  assign io_in_x746_outbuf_0_rPort_0_en_0 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@96611.4]
  assign io_in_x746_outbuf_0_rPort_0_backpressure = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@96610.4]
  assign io_in_x1159_valid = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_valid; // @[sm_x1180_outr_UnitPipe.scala 59:24:@96616.4]
  assign io_in_x1159_bits_addr = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_bits_addr; // @[sm_x1180_outr_UnitPipe.scala 59:24:@96615.4]
  assign io_in_x1159_bits_size = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_bits_size; // @[sm_x1180_outr_UnitPipe.scala 59:24:@96614.4]
  assign io_in_x1160_valid = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_valid; // @[sm_x1180_outr_UnitPipe.scala 61:24:@96621.4]
  assign io_in_x1160_bits_wdata_0 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_bits_wdata_0; // @[sm_x1180_outr_UnitPipe.scala 61:24:@96620.4]
  assign io_in_x1160_bits_wstrb = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_bits_wstrb; // @[sm_x1180_outr_UnitPipe.scala 61:24:@96619.4]
  assign io_in_x745_TVALID = x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TVALID; // @[sm_x1158_outr_UnitPipe.scala 48:23:@96308.4]
  assign io_in_x745_TDATA = x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TDATA; // @[sm_x1158_outr_UnitPipe.scala 48:23:@96306.4]
  assign io_in_x744_TREADY = x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TREADY; // @[sm_x1158_outr_UnitPipe.scala 49:23:@96316.4]
  assign io_in_x1161_ready = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1161_ready; // @[sm_x1180_outr_UnitPipe.scala 62:24:@96625.4]
  assign io_sigsOut_smDoneIn_0 = x1158_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@96223.4]
  assign io_sigsOut_smDoneIn_1 = x1180_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@96512.4]
  assign x1158_outr_UnitPipe_sm_clock = clock; // @[:@96139.4]
  assign x1158_outr_UnitPipe_sm_reset = reset; // @[:@96140.4]
  assign x1158_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@96220.4]
  assign x1158_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@96222.4]
  assign x1158_outr_UnitPipe_sm_io_doneIn_0 = x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@96190.4]
  assign x1158_outr_UnitPipe_sm_io_doneIn_1 = x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@96191.4]
  assign x1158_outr_UnitPipe_sm_io_ctrCopyDone_0 = x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@96237.4]
  assign x1158_outr_UnitPipe_sm_io_ctrCopyDone_1 = x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@96238.4]
  assign RetimeWrapper_clock = clock; // @[:@96201.4]
  assign RetimeWrapper_reset = reset; // @[:@96202.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@96204.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@96203.4]
  assign RetimeWrapper_1_clock = clock; // @[:@96209.4]
  assign RetimeWrapper_1_reset = reset; // @[:@96210.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@96212.4]
  assign RetimeWrapper_1_io_in = x1158_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@96211.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_clock = clock; // @[:@96240.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_reset = reset; // @[:@96241.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x745_TREADY = io_in_x745_TREADY; // @[sm_x1158_outr_UnitPipe.scala 48:23:@96307.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TVALID = io_in_x744_TVALID; // @[sm_x1158_outr_UnitPipe.scala 49:23:@96317.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TDATA = io_in_x744_TDATA; // @[sm_x1158_outr_UnitPipe.scala 49:23:@96315.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TID = io_in_x744_TID; // @[sm_x1158_outr_UnitPipe.scala 49:23:@96311.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_in_x744_TDEST = io_in_x744_TDEST; // @[sm_x1158_outr_UnitPipe.scala 49:23:@96310.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x1158_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x1158_outr_UnitPipe.scala 92:22:@96333.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x1158_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x1158_outr_UnitPipe.scala 92:22:@96334.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x1158_outr_UnitPipe_sm_io_childAck_0; // @[sm_x1158_outr_UnitPipe.scala 92:22:@96329.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x1158_outr_UnitPipe_sm_io_childAck_1; // @[sm_x1158_outr_UnitPipe.scala 92:22:@96330.4]
  assign x1158_outr_UnitPipe_kernelx1158_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x1158_outr_UnitPipe.scala 91:18:@96318.4]
  assign x1180_outr_UnitPipe_sm_clock = clock; // @[:@96418.4]
  assign x1180_outr_UnitPipe_sm_reset = reset; // @[:@96419.4]
  assign x1180_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@96509.4]
  assign x1180_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@96511.4]
  assign x1180_outr_UnitPipe_sm_io_doneIn_0 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@96477.4]
  assign x1180_outr_UnitPipe_sm_io_doneIn_1 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@96478.4]
  assign x1180_outr_UnitPipe_sm_io_doneIn_2 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@96479.4]
  assign x1180_outr_UnitPipe_sm_io_ctrCopyDone_0 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@96526.4]
  assign x1180_outr_UnitPipe_sm_io_ctrCopyDone_1 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@96527.4]
  assign x1180_outr_UnitPipe_sm_io_ctrCopyDone_2 = x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@96528.4]
  assign RetimeWrapper_2_clock = clock; // @[:@96490.4]
  assign RetimeWrapper_2_reset = reset; // @[:@96491.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@96493.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@96492.4]
  assign RetimeWrapper_3_clock = clock; // @[:@96498.4]
  assign RetimeWrapper_3_reset = reset; // @[:@96499.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@96501.4]
  assign RetimeWrapper_3_io_in = x1180_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@96500.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_clock = clock; // @[:@96530.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_reset = reset; // @[:@96531.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x746_outbuf_0_rPort_0_output_0 = io_in_x746_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@96609.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1159_ready = io_in_x1159_ready; // @[sm_x1180_outr_UnitPipe.scala 59:24:@96617.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x742_outdram_number = io_in_x742_outdram_number; // @[sm_x1180_outr_UnitPipe.scala 60:31:@96618.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1160_ready = io_in_x1160_ready; // @[sm_x1180_outr_UnitPipe.scala 61:24:@96622.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_in_x1161_valid = io_in_x1161_valid; // @[sm_x1180_outr_UnitPipe.scala 62:24:@96624.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x1180_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x1180_outr_UnitPipe.scala 113:22:@96648.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x1180_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x1180_outr_UnitPipe.scala 113:22:@96649.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x1180_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x1180_outr_UnitPipe.scala 113:22:@96650.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x1180_outr_UnitPipe_sm_io_childAck_0; // @[sm_x1180_outr_UnitPipe.scala 113:22:@96642.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x1180_outr_UnitPipe_sm_io_childAck_1; // @[sm_x1180_outr_UnitPipe.scala 113:22:@96643.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x1180_outr_UnitPipe_sm_io_childAck_2; // @[sm_x1180_outr_UnitPipe.scala 113:22:@96644.4]
  assign x1180_outr_UnitPipe_kernelx1180_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x1180_outr_UnitPipe.scala 112:18:@96626.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@96678.2]
  input          clock, // @[:@96679.4]
  input          reset, // @[:@96680.4]
  input          io_in_x1159_ready, // @[:@96681.4]
  output         io_in_x1159_valid, // @[:@96681.4]
  output [63:0]  io_in_x1159_bits_addr, // @[:@96681.4]
  output [31:0]  io_in_x1159_bits_size, // @[:@96681.4]
  input  [63:0]  io_in_x742_outdram_number, // @[:@96681.4]
  input          io_in_x1160_ready, // @[:@96681.4]
  output         io_in_x1160_valid, // @[:@96681.4]
  output [7:0]   io_in_x1160_bits_wdata_0, // @[:@96681.4]
  output         io_in_x1160_bits_wstrb, // @[:@96681.4]
  output         io_in_x745_TVALID, // @[:@96681.4]
  input          io_in_x745_TREADY, // @[:@96681.4]
  output [255:0] io_in_x745_TDATA, // @[:@96681.4]
  input          io_in_x744_TVALID, // @[:@96681.4]
  output         io_in_x744_TREADY, // @[:@96681.4]
  input  [255:0] io_in_x744_TDATA, // @[:@96681.4]
  input  [7:0]   io_in_x744_TID, // @[:@96681.4]
  input  [7:0]   io_in_x744_TDEST, // @[:@96681.4]
  output         io_in_x1161_ready, // @[:@96681.4]
  input          io_in_x1161_valid, // @[:@96681.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@96681.4]
  input          io_sigsIn_smChildAcks_0, // @[:@96681.4]
  output         io_sigsOut_smDoneIn_0, // @[:@96681.4]
  input          io_rr // @[:@96681.4]
);
  wire  x746_outbuf_0_clock; // @[m_x746_outbuf_0.scala 27:17:@96691.4]
  wire  x746_outbuf_0_reset; // @[m_x746_outbuf_0.scala 27:17:@96691.4]
  wire [20:0] x746_outbuf_0_io_rPort_0_ofs_0; // @[m_x746_outbuf_0.scala 27:17:@96691.4]
  wire  x746_outbuf_0_io_rPort_0_en_0; // @[m_x746_outbuf_0.scala 27:17:@96691.4]
  wire  x746_outbuf_0_io_rPort_0_backpressure; // @[m_x746_outbuf_0.scala 27:17:@96691.4]
  wire [7:0] x746_outbuf_0_io_rPort_0_output_0; // @[m_x746_outbuf_0.scala 27:17:@96691.4]
  wire  x1251_sm_clock; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_reset; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_enable; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_done; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_ctrDone; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_ctrInc; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_parentAck; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_doneIn_0; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_doneIn_1; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_enableOut_0; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_enableOut_1; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_childAck_0; // @[sm_x1251.scala 37:18:@96749.4]
  wire  x1251_sm_io_childAck_1; // @[sm_x1251.scala 37:18:@96749.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@96816.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@96816.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@96816.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@96816.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@96816.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@96824.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@96824.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@96824.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@96824.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@96824.4]
  wire  x1251_kernelx1251_concrete1_clock; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_reset; // @[sm_x1251.scala 102:24:@96853.4]
  wire [20:0] x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_en_0; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure; // @[sm_x1251.scala 102:24:@96853.4]
  wire [7:0] x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_output_0; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x1159_ready; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x1159_valid; // @[sm_x1251.scala 102:24:@96853.4]
  wire [63:0] x1251_kernelx1251_concrete1_io_in_x1159_bits_addr; // @[sm_x1251.scala 102:24:@96853.4]
  wire [31:0] x1251_kernelx1251_concrete1_io_in_x1159_bits_size; // @[sm_x1251.scala 102:24:@96853.4]
  wire [63:0] x1251_kernelx1251_concrete1_io_in_x742_outdram_number; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x1160_ready; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x1160_valid; // @[sm_x1251.scala 102:24:@96853.4]
  wire [7:0] x1251_kernelx1251_concrete1_io_in_x1160_bits_wdata_0; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x1160_bits_wstrb; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x745_TVALID; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x745_TREADY; // @[sm_x1251.scala 102:24:@96853.4]
  wire [255:0] x1251_kernelx1251_concrete1_io_in_x745_TDATA; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x744_TVALID; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x744_TREADY; // @[sm_x1251.scala 102:24:@96853.4]
  wire [255:0] x1251_kernelx1251_concrete1_io_in_x744_TDATA; // @[sm_x1251.scala 102:24:@96853.4]
  wire [7:0] x1251_kernelx1251_concrete1_io_in_x744_TID; // @[sm_x1251.scala 102:24:@96853.4]
  wire [7:0] x1251_kernelx1251_concrete1_io_in_x744_TDEST; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x1161_ready; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_in_x1161_valid; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x1251.scala 102:24:@96853.4]
  wire  x1251_kernelx1251_concrete1_io_rr; // @[sm_x1251.scala 102:24:@96853.4]
  wire  _T_266; // @[package.scala 100:49:@96782.4]
  reg  _T_269; // @[package.scala 48:56:@96783.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@96821.4 package.scala 96:25:@96822.4]
  wire  _T_289; // @[package.scala 96:25:@96829.4 package.scala 96:25:@96830.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@96832.4]
  x746_outbuf_0 x746_outbuf_0 ( // @[m_x746_outbuf_0.scala 27:17:@96691.4]
    .clock(x746_outbuf_0_clock),
    .reset(x746_outbuf_0_reset),
    .io_rPort_0_ofs_0(x746_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x746_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x746_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x746_outbuf_0_io_rPort_0_output_0)
  );
  x1251_sm x1251_sm ( // @[sm_x1251.scala 37:18:@96749.4]
    .clock(x1251_sm_clock),
    .reset(x1251_sm_reset),
    .io_enable(x1251_sm_io_enable),
    .io_done(x1251_sm_io_done),
    .io_ctrDone(x1251_sm_io_ctrDone),
    .io_ctrInc(x1251_sm_io_ctrInc),
    .io_parentAck(x1251_sm_io_parentAck),
    .io_doneIn_0(x1251_sm_io_doneIn_0),
    .io_doneIn_1(x1251_sm_io_doneIn_1),
    .io_enableOut_0(x1251_sm_io_enableOut_0),
    .io_enableOut_1(x1251_sm_io_enableOut_1),
    .io_childAck_0(x1251_sm_io_childAck_0),
    .io_childAck_1(x1251_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@96816.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@96824.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x1251_kernelx1251_concrete1 x1251_kernelx1251_concrete1 ( // @[sm_x1251.scala 102:24:@96853.4]
    .clock(x1251_kernelx1251_concrete1_clock),
    .reset(x1251_kernelx1251_concrete1_reset),
    .io_in_x746_outbuf_0_rPort_0_ofs_0(x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0),
    .io_in_x746_outbuf_0_rPort_0_en_0(x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_en_0),
    .io_in_x746_outbuf_0_rPort_0_backpressure(x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure),
    .io_in_x746_outbuf_0_rPort_0_output_0(x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_output_0),
    .io_in_x1159_ready(x1251_kernelx1251_concrete1_io_in_x1159_ready),
    .io_in_x1159_valid(x1251_kernelx1251_concrete1_io_in_x1159_valid),
    .io_in_x1159_bits_addr(x1251_kernelx1251_concrete1_io_in_x1159_bits_addr),
    .io_in_x1159_bits_size(x1251_kernelx1251_concrete1_io_in_x1159_bits_size),
    .io_in_x742_outdram_number(x1251_kernelx1251_concrete1_io_in_x742_outdram_number),
    .io_in_x1160_ready(x1251_kernelx1251_concrete1_io_in_x1160_ready),
    .io_in_x1160_valid(x1251_kernelx1251_concrete1_io_in_x1160_valid),
    .io_in_x1160_bits_wdata_0(x1251_kernelx1251_concrete1_io_in_x1160_bits_wdata_0),
    .io_in_x1160_bits_wstrb(x1251_kernelx1251_concrete1_io_in_x1160_bits_wstrb),
    .io_in_x745_TVALID(x1251_kernelx1251_concrete1_io_in_x745_TVALID),
    .io_in_x745_TREADY(x1251_kernelx1251_concrete1_io_in_x745_TREADY),
    .io_in_x745_TDATA(x1251_kernelx1251_concrete1_io_in_x745_TDATA),
    .io_in_x744_TVALID(x1251_kernelx1251_concrete1_io_in_x744_TVALID),
    .io_in_x744_TREADY(x1251_kernelx1251_concrete1_io_in_x744_TREADY),
    .io_in_x744_TDATA(x1251_kernelx1251_concrete1_io_in_x744_TDATA),
    .io_in_x744_TID(x1251_kernelx1251_concrete1_io_in_x744_TID),
    .io_in_x744_TDEST(x1251_kernelx1251_concrete1_io_in_x744_TDEST),
    .io_in_x1161_ready(x1251_kernelx1251_concrete1_io_in_x1161_ready),
    .io_in_x1161_valid(x1251_kernelx1251_concrete1_io_in_x1161_valid),
    .io_sigsIn_smEnableOuts_0(x1251_kernelx1251_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x1251_kernelx1251_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x1251_kernelx1251_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x1251_kernelx1251_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x1251_kernelx1251_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x1251_kernelx1251_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x1251_kernelx1251_concrete1_io_rr)
  );
  assign _T_266 = x1251_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@96782.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@96821.4 package.scala 96:25:@96822.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@96829.4 package.scala 96:25:@96830.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@96832.4]
  assign io_in_x1159_valid = x1251_kernelx1251_concrete1_io_in_x1159_valid; // @[sm_x1251.scala 64:24:@96939.4]
  assign io_in_x1159_bits_addr = x1251_kernelx1251_concrete1_io_in_x1159_bits_addr; // @[sm_x1251.scala 64:24:@96938.4]
  assign io_in_x1159_bits_size = x1251_kernelx1251_concrete1_io_in_x1159_bits_size; // @[sm_x1251.scala 64:24:@96937.4]
  assign io_in_x1160_valid = x1251_kernelx1251_concrete1_io_in_x1160_valid; // @[sm_x1251.scala 66:24:@96944.4]
  assign io_in_x1160_bits_wdata_0 = x1251_kernelx1251_concrete1_io_in_x1160_bits_wdata_0; // @[sm_x1251.scala 66:24:@96943.4]
  assign io_in_x1160_bits_wstrb = x1251_kernelx1251_concrete1_io_in_x1160_bits_wstrb; // @[sm_x1251.scala 66:24:@96942.4]
  assign io_in_x745_TVALID = x1251_kernelx1251_concrete1_io_in_x745_TVALID; // @[sm_x1251.scala 67:23:@96954.4]
  assign io_in_x745_TDATA = x1251_kernelx1251_concrete1_io_in_x745_TDATA; // @[sm_x1251.scala 67:23:@96952.4]
  assign io_in_x744_TREADY = x1251_kernelx1251_concrete1_io_in_x744_TREADY; // @[sm_x1251.scala 68:23:@96962.4]
  assign io_in_x1161_ready = x1251_kernelx1251_concrete1_io_in_x1161_ready; // @[sm_x1251.scala 69:24:@96966.4]
  assign io_sigsOut_smDoneIn_0 = x1251_sm_io_done; // @[SpatialBlocks.scala 156:53:@96839.4]
  assign x746_outbuf_0_clock = clock; // @[:@96692.4]
  assign x746_outbuf_0_reset = reset; // @[:@96693.4]
  assign x746_outbuf_0_io_rPort_0_ofs_0 = x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@96935.4]
  assign x746_outbuf_0_io_rPort_0_en_0 = x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@96934.4]
  assign x746_outbuf_0_io_rPort_0_backpressure = x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@96933.4]
  assign x1251_sm_clock = clock; // @[:@96750.4]
  assign x1251_sm_reset = reset; // @[:@96751.4]
  assign x1251_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@96836.4]
  assign x1251_sm_io_ctrDone = x1251_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:27:@96786.4]
  assign x1251_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@96838.4]
  assign x1251_sm_io_doneIn_0 = x1251_kernelx1251_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@96806.4]
  assign x1251_sm_io_doneIn_1 = x1251_kernelx1251_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@96807.4]
  assign RetimeWrapper_clock = clock; // @[:@96817.4]
  assign RetimeWrapper_reset = reset; // @[:@96818.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@96820.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@96819.4]
  assign RetimeWrapper_1_clock = clock; // @[:@96825.4]
  assign RetimeWrapper_1_reset = reset; // @[:@96826.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@96828.4]
  assign RetimeWrapper_1_io_in = x1251_sm_io_done; // @[package.scala 94:16:@96827.4]
  assign x1251_kernelx1251_concrete1_clock = clock; // @[:@96854.4]
  assign x1251_kernelx1251_concrete1_reset = reset; // @[:@96855.4]
  assign x1251_kernelx1251_concrete1_io_in_x746_outbuf_0_rPort_0_output_0 = x746_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@96932.4]
  assign x1251_kernelx1251_concrete1_io_in_x1159_ready = io_in_x1159_ready; // @[sm_x1251.scala 64:24:@96940.4]
  assign x1251_kernelx1251_concrete1_io_in_x742_outdram_number = io_in_x742_outdram_number; // @[sm_x1251.scala 65:31:@96941.4]
  assign x1251_kernelx1251_concrete1_io_in_x1160_ready = io_in_x1160_ready; // @[sm_x1251.scala 66:24:@96945.4]
  assign x1251_kernelx1251_concrete1_io_in_x745_TREADY = io_in_x745_TREADY; // @[sm_x1251.scala 67:23:@96953.4]
  assign x1251_kernelx1251_concrete1_io_in_x744_TVALID = io_in_x744_TVALID; // @[sm_x1251.scala 68:23:@96963.4]
  assign x1251_kernelx1251_concrete1_io_in_x744_TDATA = io_in_x744_TDATA; // @[sm_x1251.scala 68:23:@96961.4]
  assign x1251_kernelx1251_concrete1_io_in_x744_TID = io_in_x744_TID; // @[sm_x1251.scala 68:23:@96957.4]
  assign x1251_kernelx1251_concrete1_io_in_x744_TDEST = io_in_x744_TDEST; // @[sm_x1251.scala 68:23:@96956.4]
  assign x1251_kernelx1251_concrete1_io_in_x1161_valid = io_in_x1161_valid; // @[sm_x1251.scala 69:24:@96965.4]
  assign x1251_kernelx1251_concrete1_io_sigsIn_smEnableOuts_0 = x1251_sm_io_enableOut_0; // @[sm_x1251.scala 107:22:@96977.4]
  assign x1251_kernelx1251_concrete1_io_sigsIn_smEnableOuts_1 = x1251_sm_io_enableOut_1; // @[sm_x1251.scala 107:22:@96978.4]
  assign x1251_kernelx1251_concrete1_io_sigsIn_smChildAcks_0 = x1251_sm_io_childAck_0; // @[sm_x1251.scala 107:22:@96973.4]
  assign x1251_kernelx1251_concrete1_io_sigsIn_smChildAcks_1 = x1251_sm_io_childAck_1; // @[sm_x1251.scala 107:22:@96974.4]
  assign x1251_kernelx1251_concrete1_io_rr = io_rr; // @[sm_x1251.scala 106:18:@96967.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@97000.2]
  input          clock, // @[:@97001.4]
  input          reset, // @[:@97002.4]
  input          io_enable, // @[:@97003.4]
  output         io_done, // @[:@97003.4]
  input          io_reset, // @[:@97003.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@97003.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@97003.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@97003.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@97003.4]
  output         io_memStreams_loads_0_data_ready, // @[:@97003.4]
  input          io_memStreams_loads_0_data_valid, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@97003.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@97003.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@97003.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@97003.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@97003.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@97003.4]
  input          io_memStreams_stores_0_data_ready, // @[:@97003.4]
  output         io_memStreams_stores_0_data_valid, // @[:@97003.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_0, // @[:@97003.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@97003.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@97003.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@97003.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@97003.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@97003.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@97003.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@97003.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@97003.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@97003.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@97003.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@97003.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@97003.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@97003.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@97003.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@97003.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@97003.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@97003.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@97003.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@97003.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@97003.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@97003.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@97003.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@97003.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@97003.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@97003.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@97003.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@97003.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@97003.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@97003.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@97003.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@97003.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@97003.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@97003.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@97003.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@97003.4]
  output         io_heap_0_req_valid, // @[:@97003.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@97003.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@97003.4]
  input          io_heap_0_resp_valid, // @[:@97003.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@97003.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@97003.4]
  input  [63:0]  io_argIns_0, // @[:@97003.4]
  input  [63:0]  io_argIns_1, // @[:@97003.4]
  input          io_argOuts_0_port_ready, // @[:@97003.4]
  output         io_argOuts_0_port_valid, // @[:@97003.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@97003.4]
  input  [63:0]  io_argOuts_0_echo // @[:@97003.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@97151.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@97151.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@97151.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@97151.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@97169.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@97169.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@97169.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@97169.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@97169.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@97178.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@97178.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@97178.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@97178.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@97178.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@97178.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@97217.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@97249.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@97249.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@97249.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@97249.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@97249.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x1159_ready; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x1159_valid; // @[sm_RootController.scala 91:24:@97311.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x1159_bits_addr; // @[sm_RootController.scala 91:24:@97311.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x1159_bits_size; // @[sm_RootController.scala 91:24:@97311.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x742_outdram_number; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x1160_ready; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x1160_valid; // @[sm_RootController.scala 91:24:@97311.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x1160_bits_wdata_0; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x1160_bits_wstrb; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x745_TVALID; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x745_TREADY; // @[sm_RootController.scala 91:24:@97311.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x745_TDATA; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x744_TVALID; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x744_TREADY; // @[sm_RootController.scala 91:24:@97311.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x744_TDATA; // @[sm_RootController.scala 91:24:@97311.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x744_TID; // @[sm_RootController.scala 91:24:@97311.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x744_TDEST; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x1161_ready; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_in_x1161_valid; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@97311.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@97311.4]
  wire  _T_599; // @[package.scala 96:25:@97174.4 package.scala 96:25:@97175.4]
  wire  _T_664; // @[Main.scala 46:50:@97245.4]
  wire  _T_665; // @[Main.scala 46:59:@97246.4]
  wire  _T_677; // @[package.scala 100:49:@97266.4]
  reg  _T_680; // @[package.scala 48:56:@97267.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@97151.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@97169.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@97178.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@97217.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@97249.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@97311.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x1159_ready(RootController_kernelRootController_concrete1_io_in_x1159_ready),
    .io_in_x1159_valid(RootController_kernelRootController_concrete1_io_in_x1159_valid),
    .io_in_x1159_bits_addr(RootController_kernelRootController_concrete1_io_in_x1159_bits_addr),
    .io_in_x1159_bits_size(RootController_kernelRootController_concrete1_io_in_x1159_bits_size),
    .io_in_x742_outdram_number(RootController_kernelRootController_concrete1_io_in_x742_outdram_number),
    .io_in_x1160_ready(RootController_kernelRootController_concrete1_io_in_x1160_ready),
    .io_in_x1160_valid(RootController_kernelRootController_concrete1_io_in_x1160_valid),
    .io_in_x1160_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x1160_bits_wdata_0),
    .io_in_x1160_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x1160_bits_wstrb),
    .io_in_x745_TVALID(RootController_kernelRootController_concrete1_io_in_x745_TVALID),
    .io_in_x745_TREADY(RootController_kernelRootController_concrete1_io_in_x745_TREADY),
    .io_in_x745_TDATA(RootController_kernelRootController_concrete1_io_in_x745_TDATA),
    .io_in_x744_TVALID(RootController_kernelRootController_concrete1_io_in_x744_TVALID),
    .io_in_x744_TREADY(RootController_kernelRootController_concrete1_io_in_x744_TREADY),
    .io_in_x744_TDATA(RootController_kernelRootController_concrete1_io_in_x744_TDATA),
    .io_in_x744_TID(RootController_kernelRootController_concrete1_io_in_x744_TID),
    .io_in_x744_TDEST(RootController_kernelRootController_concrete1_io_in_x744_TDEST),
    .io_in_x1161_ready(RootController_kernelRootController_concrete1_io_in_x1161_ready),
    .io_in_x1161_valid(RootController_kernelRootController_concrete1_io_in_x1161_valid),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@97174.4 package.scala 96:25:@97175.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@97245.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@97246.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@97266.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@97265.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x1159_valid; // @[sm_RootController.scala 60:24:@97374.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x1159_bits_addr; // @[sm_RootController.scala 60:24:@97373.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x1159_bits_size; // @[sm_RootController.scala 60:24:@97372.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x1160_valid; // @[sm_RootController.scala 62:24:@97379.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x1160_bits_wdata_0; // @[sm_RootController.scala 62:24:@97378.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x1160_bits_wstrb; // @[sm_RootController.scala 62:24:@97377.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x1161_ready; // @[sm_RootController.scala 65:24:@97401.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x744_TREADY; // @[sm_RootController.scala 64:23:@97397.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x745_TVALID; // @[sm_RootController.scala 63:23:@97389.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x745_TDATA; // @[sm_RootController.scala 63:23:@97387.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 63:23:@97386.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 63:23:@97385.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 63:23:@97384.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 63:23:@97383.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 63:23:@97382.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 63:23:@97381.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@97152.4]
  assign SingleCounter_reset = reset; // @[:@97153.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@97167.4]
  assign RetimeWrapper_clock = clock; // @[:@97170.4]
  assign RetimeWrapper_reset = reset; // @[:@97171.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@97173.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@97172.4]
  assign SRFF_clock = clock; // @[:@97179.4]
  assign SRFF_reset = reset; // @[:@97180.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@97429.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@97263.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@97264.4]
  assign RootController_sm_clock = clock; // @[:@97218.4]
  assign RootController_sm_reset = reset; // @[:@97219.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@97262.4 SpatialBlocks.scala 140:18:@97296.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@97290.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@97270.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@97258.4 SpatialBlocks.scala 142:21:@97298.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@97287.4]
  assign RetimeWrapper_1_clock = clock; // @[:@97250.4]
  assign RetimeWrapper_1_reset = reset; // @[:@97251.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@97253.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@97252.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@97312.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@97313.4]
  assign RootController_kernelRootController_concrete1_io_in_x1159_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 60:24:@97375.4]
  assign RootController_kernelRootController_concrete1_io_in_x742_outdram_number = io_argIns_1; // @[sm_RootController.scala 61:31:@97376.4]
  assign RootController_kernelRootController_concrete1_io_in_x1160_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 62:24:@97380.4]
  assign RootController_kernelRootController_concrete1_io_in_x745_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 63:23:@97388.4]
  assign RootController_kernelRootController_concrete1_io_in_x744_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 64:23:@97398.4]
  assign RootController_kernelRootController_concrete1_io_in_x744_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 64:23:@97396.4]
  assign RootController_kernelRootController_concrete1_io_in_x744_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 64:23:@97392.4]
  assign RootController_kernelRootController_concrete1_io_in_x744_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 64:23:@97391.4]
  assign RootController_kernelRootController_concrete1_io_in_x1161_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 65:24:@97400.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@97410.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@97408.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@97402.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@97431.2]
  input         clock, // @[:@97432.4]
  input         reset, // @[:@97433.4]
  input  [31:0] io_raddr, // @[:@97434.4]
  input         io_wen, // @[:@97434.4]
  input  [31:0] io_waddr, // @[:@97434.4]
  input  [63:0] io_wdata, // @[:@97434.4]
  output [63:0] io_rdata // @[:@97434.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@97436.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@97436.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@97436.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@97436.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@97436.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@97436.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@97436.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@97436.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@97436.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@97436.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@97436.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@97437.4]
  assign accel_reset = reset; // @[:@97438.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
