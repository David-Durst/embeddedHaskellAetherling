// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x353_TREADY(dontcare), // @[:@1298.4]
    .io_in_x353_TDATA({I_0,I_1,I_2,I_3}), // @[:@1298.4]
    .io_in_x353_TID(8'h0),
    .io_in_x353_TDEST(8'h0),
    .io_in_x354_TVALID(valid_down), // @[:@1298.4]
    .io_in_x354_TDATA({O_0,O_1,O_2,O_3}), // @[:@1298.4]
    .io_in_x354_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x361_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule


module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh48); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh48); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x355_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x724_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x647_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x356_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x357_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x361_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x387_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x696_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x367_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x387_inr_Foreach_kernelx387_inr_Foreach_concrete1( // @[:@5894.2]
  input         clock, // @[:@5895.4]
  input         reset, // @[:@5896.4]
  output        io_in_x357_fifoinpacked_0_wPort_0_en_0, // @[:@5897.4]
  input         io_in_x357_fifoinpacked_0_full, // @[:@5897.4]
  output        io_in_x357_fifoinpacked_0_active_0_in, // @[:@5897.4]
  input         io_in_x357_fifoinpacked_0_active_0_out, // @[:@5897.4]
  input         io_sigsIn_backpressure, // @[:@5897.4]
  input         io_sigsIn_datapathEn, // @[:@5897.4]
  input         io_sigsIn_break, // @[:@5897.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@5897.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5897.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5897.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@5897.4]
  input         io_rr // @[:@5897.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@5931.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@5931.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@5943.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@5943.4]
  wire  x696_sub_1_clock; // @[Math.scala 191:24:@5970.4]
  wire  x696_sub_1_reset; // @[Math.scala 191:24:@5970.4]
  wire [31:0] x696_sub_1_io_a; // @[Math.scala 191:24:@5970.4]
  wire [31:0] x696_sub_1_io_b; // @[Math.scala 191:24:@5970.4]
  wire  x696_sub_1_io_flow; // @[Math.scala 191:24:@5970.4]
  wire [31:0] x696_sub_1_io_result; // @[Math.scala 191:24:@5970.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5980.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5980.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5980.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5980.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5980.4]
  wire  x367_sum_1_clock; // @[Math.scala 150:24:@5989.4]
  wire  x367_sum_1_reset; // @[Math.scala 150:24:@5989.4]
  wire [31:0] x367_sum_1_io_a; // @[Math.scala 150:24:@5989.4]
  wire [31:0] x367_sum_1_io_b; // @[Math.scala 150:24:@5989.4]
  wire  x367_sum_1_io_flow; // @[Math.scala 150:24:@5989.4]
  wire [31:0] x367_sum_1_io_result; // @[Math.scala 150:24:@5989.4]
  wire  x368_sum_1_clock; // @[Math.scala 150:24:@6001.4]
  wire  x368_sum_1_reset; // @[Math.scala 150:24:@6001.4]
  wire [31:0] x368_sum_1_io_a; // @[Math.scala 150:24:@6001.4]
  wire [31:0] x368_sum_1_io_b; // @[Math.scala 150:24:@6001.4]
  wire  x368_sum_1_io_flow; // @[Math.scala 150:24:@6001.4]
  wire [31:0] x368_sum_1_io_result; // @[Math.scala 150:24:@6001.4]
  wire  x698_sum_1_clock; // @[Math.scala 150:24:@6016.4]
  wire  x698_sum_1_reset; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x698_sum_1_io_a; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x698_sum_1_io_b; // @[Math.scala 150:24:@6016.4]
  wire  x698_sum_1_io_flow; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x698_sum_1_io_result; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x371_1_io_b; // @[Math.scala 720:24:@6037.4]
  wire [31:0] x371_1_io_result; // @[Math.scala 720:24:@6037.4]
  wire  x372_sum_1_clock; // @[Math.scala 150:24:@6048.4]
  wire  x372_sum_1_reset; // @[Math.scala 150:24:@6048.4]
  wire [31:0] x372_sum_1_io_a; // @[Math.scala 150:24:@6048.4]
  wire [31:0] x372_sum_1_io_b; // @[Math.scala 150:24:@6048.4]
  wire  x372_sum_1_io_flow; // @[Math.scala 150:24:@6048.4]
  wire [31:0] x372_sum_1_io_result; // @[Math.scala 150:24:@6048.4]
  wire  x701_sum_1_clock; // @[Math.scala 150:24:@6063.4]
  wire  x701_sum_1_reset; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x701_sum_1_io_a; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x701_sum_1_io_b; // @[Math.scala 150:24:@6063.4]
  wire  x701_sum_1_io_flow; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x701_sum_1_io_result; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x375_1_io_b; // @[Math.scala 720:24:@6084.4]
  wire [31:0] x375_1_io_result; // @[Math.scala 720:24:@6084.4]
  wire  x376_sum_1_clock; // @[Math.scala 150:24:@6095.4]
  wire  x376_sum_1_reset; // @[Math.scala 150:24:@6095.4]
  wire [31:0] x376_sum_1_io_a; // @[Math.scala 150:24:@6095.4]
  wire [31:0] x376_sum_1_io_b; // @[Math.scala 150:24:@6095.4]
  wire  x376_sum_1_io_flow; // @[Math.scala 150:24:@6095.4]
  wire [31:0] x376_sum_1_io_result; // @[Math.scala 150:24:@6095.4]
  wire  x704_sum_1_clock; // @[Math.scala 150:24:@6110.4]
  wire  x704_sum_1_reset; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x704_sum_1_io_a; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x704_sum_1_io_b; // @[Math.scala 150:24:@6110.4]
  wire  x704_sum_1_io_flow; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x704_sum_1_io_result; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x379_1_io_b; // @[Math.scala 720:24:@6131.4]
  wire [31:0] x379_1_io_result; // @[Math.scala 720:24:@6131.4]
  wire  x380_sum_1_clock; // @[Math.scala 150:24:@6142.4]
  wire  x380_sum_1_reset; // @[Math.scala 150:24:@6142.4]
  wire [31:0] x380_sum_1_io_a; // @[Math.scala 150:24:@6142.4]
  wire [31:0] x380_sum_1_io_b; // @[Math.scala 150:24:@6142.4]
  wire  x380_sum_1_io_flow; // @[Math.scala 150:24:@6142.4]
  wire [31:0] x380_sum_1_io_result; // @[Math.scala 150:24:@6142.4]
  wire  x707_sum_1_clock; // @[Math.scala 150:24:@6157.4]
  wire  x707_sum_1_reset; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x707_sum_1_io_a; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x707_sum_1_io_b; // @[Math.scala 150:24:@6157.4]
  wire  x707_sum_1_io_flow; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x707_sum_1_io_result; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x383_1_io_b; // @[Math.scala 720:24:@6178.4]
  wire [31:0] x383_1_io_result; // @[Math.scala 720:24:@6178.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6217.4]
  wire  _T_327; // @[sm_x387_inr_Foreach.scala 62:18:@5956.4]
  wire  _T_328; // @[sm_x387_inr_Foreach.scala 62:55:@5957.4]
  wire [31:0] b362_number; // @[Math.scala 723:22:@5936.4 Math.scala 724:14:@5937.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@5961.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@5961.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@5966.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@5966.4]
  wire [31:0] x368_sum_number; // @[Math.scala 154:22:@6007.4 Math.scala 155:14:@6008.4]
  wire [33:0] _GEN_2; // @[Math.scala 461:32:@6012.4]
  wire [33:0] _T_353; // @[Math.scala 461:32:@6012.4]
  wire [31:0] x698_sum_number; // @[Math.scala 154:22:@6022.4 Math.scala 155:14:@6023.4]
  wire [31:0] _T_364; // @[Math.scala 406:49:@6029.4]
  wire [31:0] _T_366; // @[Math.scala 406:56:@6031.4]
  wire [31:0] _T_367; // @[Math.scala 406:56:@6032.4]
  wire [31:0] x372_sum_number; // @[Math.scala 154:22:@6054.4 Math.scala 155:14:@6055.4]
  wire [33:0] _GEN_3; // @[Math.scala 461:32:@6059.4]
  wire [33:0] _T_381; // @[Math.scala 461:32:@6059.4]
  wire [31:0] x701_sum_number; // @[Math.scala 154:22:@6069.4 Math.scala 155:14:@6070.4]
  wire [31:0] _T_392; // @[Math.scala 406:49:@6076.4]
  wire [31:0] _T_394; // @[Math.scala 406:56:@6078.4]
  wire [31:0] _T_395; // @[Math.scala 406:56:@6079.4]
  wire [31:0] x376_sum_number; // @[Math.scala 154:22:@6101.4 Math.scala 155:14:@6102.4]
  wire [33:0] _GEN_4; // @[Math.scala 461:32:@6106.4]
  wire [33:0] _T_409; // @[Math.scala 461:32:@6106.4]
  wire [31:0] x704_sum_number; // @[Math.scala 154:22:@6116.4 Math.scala 155:14:@6117.4]
  wire [31:0] _T_420; // @[Math.scala 406:49:@6123.4]
  wire [31:0] _T_422; // @[Math.scala 406:56:@6125.4]
  wire [31:0] _T_423; // @[Math.scala 406:56:@6126.4]
  wire [31:0] x380_sum_number; // @[Math.scala 154:22:@6148.4 Math.scala 155:14:@6149.4]
  wire [33:0] _GEN_5; // @[Math.scala 461:32:@6153.4]
  wire [33:0] _T_437; // @[Math.scala 461:32:@6153.4]
  wire [31:0] x707_sum_number; // @[Math.scala 154:22:@6163.4 Math.scala 155:14:@6164.4]
  wire [31:0] _T_448; // @[Math.scala 406:49:@6170.4]
  wire [31:0] _T_450; // @[Math.scala 406:56:@6172.4]
  wire [31:0] _T_451; // @[Math.scala 406:56:@6173.4]
  wire  _T_475; // @[sm_x387_inr_Foreach.scala 123:131:@6214.4]
  wire  _T_479; // @[package.scala 96:25:@6222.4 package.scala 96:25:@6223.4]
  wire  _T_481; // @[implicits.scala 55:10:@6224.4]
  wire  _T_482; // @[sm_x387_inr_Foreach.scala 123:148:@6225.4]
  wire  _T_484; // @[sm_x387_inr_Foreach.scala 123:236:@6227.4]
  wire  _T_485; // @[sm_x387_inr_Foreach.scala 123:255:@6228.4]
  wire  x727_b364_D4; // @[package.scala 96:25:@6202.4 package.scala 96:25:@6203.4]
  wire  _T_488; // @[sm_x387_inr_Foreach.scala 123:291:@6230.4]
  wire  x728_b365_D4; // @[package.scala 96:25:@6211.4 package.scala 96:25:@6212.4]
  _ _ ( // @[Math.scala 720:24:@5931.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@5943.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x696_sub x696_sub_1 ( // @[Math.scala 191:24:@5970.4]
    .clock(x696_sub_1_clock),
    .reset(x696_sub_1_reset),
    .io_a(x696_sub_1_io_a),
    .io_b(x696_sub_1_io_b),
    .io_flow(x696_sub_1_io_flow),
    .io_result(x696_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@5980.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x367_sum x367_sum_1 ( // @[Math.scala 150:24:@5989.4]
    .clock(x367_sum_1_clock),
    .reset(x367_sum_1_reset),
    .io_a(x367_sum_1_io_a),
    .io_b(x367_sum_1_io_b),
    .io_flow(x367_sum_1_io_flow),
    .io_result(x367_sum_1_io_result)
  );
  x367_sum x368_sum_1 ( // @[Math.scala 150:24:@6001.4]
    .clock(x368_sum_1_clock),
    .reset(x368_sum_1_reset),
    .io_a(x368_sum_1_io_a),
    .io_b(x368_sum_1_io_b),
    .io_flow(x368_sum_1_io_flow),
    .io_result(x368_sum_1_io_result)
  );
  x367_sum x698_sum_1 ( // @[Math.scala 150:24:@6016.4]
    .clock(x698_sum_1_clock),
    .reset(x698_sum_1_reset),
    .io_a(x698_sum_1_io_a),
    .io_b(x698_sum_1_io_b),
    .io_flow(x698_sum_1_io_flow),
    .io_result(x698_sum_1_io_result)
  );
  _ x371_1 ( // @[Math.scala 720:24:@6037.4]
    .io_b(x371_1_io_b),
    .io_result(x371_1_io_result)
  );
  x367_sum x372_sum_1 ( // @[Math.scala 150:24:@6048.4]
    .clock(x372_sum_1_clock),
    .reset(x372_sum_1_reset),
    .io_a(x372_sum_1_io_a),
    .io_b(x372_sum_1_io_b),
    .io_flow(x372_sum_1_io_flow),
    .io_result(x372_sum_1_io_result)
  );
  x367_sum x701_sum_1 ( // @[Math.scala 150:24:@6063.4]
    .clock(x701_sum_1_clock),
    .reset(x701_sum_1_reset),
    .io_a(x701_sum_1_io_a),
    .io_b(x701_sum_1_io_b),
    .io_flow(x701_sum_1_io_flow),
    .io_result(x701_sum_1_io_result)
  );
  _ x375_1 ( // @[Math.scala 720:24:@6084.4]
    .io_b(x375_1_io_b),
    .io_result(x375_1_io_result)
  );
  x367_sum x376_sum_1 ( // @[Math.scala 150:24:@6095.4]
    .clock(x376_sum_1_clock),
    .reset(x376_sum_1_reset),
    .io_a(x376_sum_1_io_a),
    .io_b(x376_sum_1_io_b),
    .io_flow(x376_sum_1_io_flow),
    .io_result(x376_sum_1_io_result)
  );
  x367_sum x704_sum_1 ( // @[Math.scala 150:24:@6110.4]
    .clock(x704_sum_1_clock),
    .reset(x704_sum_1_reset),
    .io_a(x704_sum_1_io_a),
    .io_b(x704_sum_1_io_b),
    .io_flow(x704_sum_1_io_flow),
    .io_result(x704_sum_1_io_result)
  );
  _ x379_1 ( // @[Math.scala 720:24:@6131.4]
    .io_b(x379_1_io_b),
    .io_result(x379_1_io_result)
  );
  x367_sum x380_sum_1 ( // @[Math.scala 150:24:@6142.4]
    .clock(x380_sum_1_clock),
    .reset(x380_sum_1_reset),
    .io_a(x380_sum_1_io_a),
    .io_b(x380_sum_1_io_b),
    .io_flow(x380_sum_1_io_flow),
    .io_result(x380_sum_1_io_result)
  );
  x367_sum x707_sum_1 ( // @[Math.scala 150:24:@6157.4]
    .clock(x707_sum_1_clock),
    .reset(x707_sum_1_reset),
    .io_a(x707_sum_1_io_a),
    .io_b(x707_sum_1_io_b),
    .io_flow(x707_sum_1_io_flow),
    .io_result(x707_sum_1_io_result)
  );
  _ x383_1 ( // @[Math.scala 720:24:@6178.4]
    .io_b(x383_1_io_b),
    .io_result(x383_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@6197.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@6206.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@6217.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x357_fifoinpacked_0_full; // @[sm_x387_inr_Foreach.scala 62:18:@5956.4]
  assign _T_328 = ~ io_in_x357_fifoinpacked_0_active_0_out; // @[sm_x387_inr_Foreach.scala 62:55:@5957.4]
  assign b362_number = __io_result; // @[Math.scala 723:22:@5936.4 Math.scala 724:14:@5937.4]
  assign _GEN_0 = {{11'd0}, b362_number}; // @[Math.scala 461:32:@5961.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@5961.4]
  assign _GEN_1 = {{7'd0}, b362_number}; // @[Math.scala 461:32:@5966.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@5966.4]
  assign x368_sum_number = x368_sum_1_io_result; // @[Math.scala 154:22:@6007.4 Math.scala 155:14:@6008.4]
  assign _GEN_2 = {{2'd0}, x368_sum_number}; // @[Math.scala 461:32:@6012.4]
  assign _T_353 = _GEN_2 << 2; // @[Math.scala 461:32:@6012.4]
  assign x698_sum_number = x698_sum_1_io_result; // @[Math.scala 154:22:@6022.4 Math.scala 155:14:@6023.4]
  assign _T_364 = $signed(x698_sum_number); // @[Math.scala 406:49:@6029.4]
  assign _T_366 = $signed(_T_364) & $signed(32'shff); // @[Math.scala 406:56:@6031.4]
  assign _T_367 = $signed(_T_366); // @[Math.scala 406:56:@6032.4]
  assign x372_sum_number = x372_sum_1_io_result; // @[Math.scala 154:22:@6054.4 Math.scala 155:14:@6055.4]
  assign _GEN_3 = {{2'd0}, x372_sum_number}; // @[Math.scala 461:32:@6059.4]
  assign _T_381 = _GEN_3 << 2; // @[Math.scala 461:32:@6059.4]
  assign x701_sum_number = x701_sum_1_io_result; // @[Math.scala 154:22:@6069.4 Math.scala 155:14:@6070.4]
  assign _T_392 = $signed(x701_sum_number); // @[Math.scala 406:49:@6076.4]
  assign _T_394 = $signed(_T_392) & $signed(32'shff); // @[Math.scala 406:56:@6078.4]
  assign _T_395 = $signed(_T_394); // @[Math.scala 406:56:@6079.4]
  assign x376_sum_number = x376_sum_1_io_result; // @[Math.scala 154:22:@6101.4 Math.scala 155:14:@6102.4]
  assign _GEN_4 = {{2'd0}, x376_sum_number}; // @[Math.scala 461:32:@6106.4]
  assign _T_409 = _GEN_4 << 2; // @[Math.scala 461:32:@6106.4]
  assign x704_sum_number = x704_sum_1_io_result; // @[Math.scala 154:22:@6116.4 Math.scala 155:14:@6117.4]
  assign _T_420 = $signed(x704_sum_number); // @[Math.scala 406:49:@6123.4]
  assign _T_422 = $signed(_T_420) & $signed(32'shff); // @[Math.scala 406:56:@6125.4]
  assign _T_423 = $signed(_T_422); // @[Math.scala 406:56:@6126.4]
  assign x380_sum_number = x380_sum_1_io_result; // @[Math.scala 154:22:@6148.4 Math.scala 155:14:@6149.4]
  assign _GEN_5 = {{2'd0}, x380_sum_number}; // @[Math.scala 461:32:@6153.4]
  assign _T_437 = _GEN_5 << 2; // @[Math.scala 461:32:@6153.4]
  assign x707_sum_number = x707_sum_1_io_result; // @[Math.scala 154:22:@6163.4 Math.scala 155:14:@6164.4]
  assign _T_448 = $signed(x707_sum_number); // @[Math.scala 406:49:@6170.4]
  assign _T_450 = $signed(_T_448) & $signed(32'shff); // @[Math.scala 406:56:@6172.4]
  assign _T_451 = $signed(_T_450); // @[Math.scala 406:56:@6173.4]
  assign _T_475 = ~ io_sigsIn_break; // @[sm_x387_inr_Foreach.scala 123:131:@6214.4]
  assign _T_479 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@6222.4 package.scala 96:25:@6223.4]
  assign _T_481 = io_rr ? _T_479 : 1'h0; // @[implicits.scala 55:10:@6224.4]
  assign _T_482 = _T_475 & _T_481; // @[sm_x387_inr_Foreach.scala 123:148:@6225.4]
  assign _T_484 = _T_482 & _T_475; // @[sm_x387_inr_Foreach.scala 123:236:@6227.4]
  assign _T_485 = _T_484 & io_sigsIn_backpressure; // @[sm_x387_inr_Foreach.scala 123:255:@6228.4]
  assign x727_b364_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6202.4 package.scala 96:25:@6203.4]
  assign _T_488 = _T_485 & x727_b364_D4; // @[sm_x387_inr_Foreach.scala 123:291:@6230.4]
  assign x728_b365_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@6211.4 package.scala 96:25:@6212.4]
  assign io_in_x357_fifoinpacked_0_wPort_0_en_0 = _T_488 & x728_b365_D4; // @[MemInterfaceType.scala 93:57:@6234.4]
  assign io_in_x357_fifoinpacked_0_active_0_in = x727_b364_D4 & x728_b365_D4; // @[MemInterfaceType.scala 147:18:@6237.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@5934.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@5946.4]
  assign x696_sub_1_clock = clock; // @[:@5971.4]
  assign x696_sub_1_reset = reset; // @[:@5972.4]
  assign x696_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@5973.4]
  assign x696_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@5974.4]
  assign x696_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@5975.4]
  assign RetimeWrapper_clock = clock; // @[:@5981.4]
  assign RetimeWrapper_reset = reset; // @[:@5982.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5984.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@5983.4]
  assign x367_sum_1_clock = clock; // @[:@5990.4]
  assign x367_sum_1_reset = reset; // @[:@5991.4]
  assign x367_sum_1_io_a = x696_sub_1_io_result; // @[Math.scala 151:17:@5992.4]
  assign x367_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@5993.4]
  assign x367_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5994.4]
  assign x368_sum_1_clock = clock; // @[:@6002.4]
  assign x368_sum_1_reset = reset; // @[:@6003.4]
  assign x368_sum_1_io_a = x367_sum_1_io_result; // @[Math.scala 151:17:@6004.4]
  assign x368_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@6005.4]
  assign x368_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6006.4]
  assign x698_sum_1_clock = clock; // @[:@6017.4]
  assign x698_sum_1_reset = reset; // @[:@6018.4]
  assign x698_sum_1_io_a = _T_353[31:0]; // @[Math.scala 151:17:@6019.4]
  assign x698_sum_1_io_b = x368_sum_1_io_result; // @[Math.scala 152:17:@6020.4]
  assign x698_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6021.4]
  assign x371_1_io_b = $unsigned(_T_367); // @[Math.scala 721:17:@6040.4]
  assign x372_sum_1_clock = clock; // @[:@6049.4]
  assign x372_sum_1_reset = reset; // @[:@6050.4]
  assign x372_sum_1_io_a = x367_sum_1_io_result; // @[Math.scala 151:17:@6051.4]
  assign x372_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@6052.4]
  assign x372_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6053.4]
  assign x701_sum_1_clock = clock; // @[:@6064.4]
  assign x701_sum_1_reset = reset; // @[:@6065.4]
  assign x701_sum_1_io_a = _T_381[31:0]; // @[Math.scala 151:17:@6066.4]
  assign x701_sum_1_io_b = x372_sum_1_io_result; // @[Math.scala 152:17:@6067.4]
  assign x701_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6068.4]
  assign x375_1_io_b = $unsigned(_T_395); // @[Math.scala 721:17:@6087.4]
  assign x376_sum_1_clock = clock; // @[:@6096.4]
  assign x376_sum_1_reset = reset; // @[:@6097.4]
  assign x376_sum_1_io_a = x367_sum_1_io_result; // @[Math.scala 151:17:@6098.4]
  assign x376_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@6099.4]
  assign x376_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6100.4]
  assign x704_sum_1_clock = clock; // @[:@6111.4]
  assign x704_sum_1_reset = reset; // @[:@6112.4]
  assign x704_sum_1_io_a = _T_409[31:0]; // @[Math.scala 151:17:@6113.4]
  assign x704_sum_1_io_b = x376_sum_1_io_result; // @[Math.scala 152:17:@6114.4]
  assign x704_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6115.4]
  assign x379_1_io_b = $unsigned(_T_423); // @[Math.scala 721:17:@6134.4]
  assign x380_sum_1_clock = clock; // @[:@6143.4]
  assign x380_sum_1_reset = reset; // @[:@6144.4]
  assign x380_sum_1_io_a = x367_sum_1_io_result; // @[Math.scala 151:17:@6145.4]
  assign x380_sum_1_io_b = 32'h4; // @[Math.scala 152:17:@6146.4]
  assign x380_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6147.4]
  assign x707_sum_1_clock = clock; // @[:@6158.4]
  assign x707_sum_1_reset = reset; // @[:@6159.4]
  assign x707_sum_1_io_a = _T_437[31:0]; // @[Math.scala 151:17:@6160.4]
  assign x707_sum_1_io_b = x380_sum_1_io_result; // @[Math.scala 152:17:@6161.4]
  assign x707_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6162.4]
  assign x383_1_io_b = $unsigned(_T_451); // @[Math.scala 721:17:@6181.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6198.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6199.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6201.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@6200.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6207.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6208.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6210.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@6209.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6218.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6219.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6221.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6220.4]
endmodule
module RetimeWrapper_48( // @[:@7355.2]
  input   clock, // @[:@7356.4]
  input   reset, // @[:@7357.4]
  input   io_flow, // @[:@7358.4]
  input   io_in, // @[:@7358.4]
  output  io_out // @[:@7358.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(73)) sr ( // @[RetimeShiftRegister.scala 15:20:@7360.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7373.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7372.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@7371.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7370.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7369.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7367.4]
endmodule
module RetimeWrapper_52( // @[:@7483.2]
  input   clock, // @[:@7484.4]
  input   reset, // @[:@7485.4]
  input   io_flow, // @[:@7486.4]
  input   io_in, // @[:@7486.4]
  output  io_out // @[:@7486.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(72)) sr ( // @[RetimeShiftRegister.scala 15:20:@7488.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7501.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7500.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@7499.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7498.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7497.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7495.4]
endmodule
module x645_inr_Foreach_SAMPLER_BOX_sm( // @[:@7503.2]
  input   clock, // @[:@7504.4]
  input   reset, // @[:@7505.4]
  input   io_enable, // @[:@7506.4]
  output  io_done, // @[:@7506.4]
  output  io_doneLatch, // @[:@7506.4]
  input   io_ctrDone, // @[:@7506.4]
  output  io_datapathEn, // @[:@7506.4]
  output  io_ctrInc, // @[:@7506.4]
  output  io_ctrRst, // @[:@7506.4]
  input   io_parentAck, // @[:@7506.4]
  input   io_backpressure, // @[:@7506.4]
  input   io_break // @[:@7506.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@7508.4]
  wire  active_reset; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@7508.4]
  wire  done_clock; // @[Controllers.scala 262:20:@7511.4]
  wire  done_reset; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@7511.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@7603.4]
  wire  _T_80; // @[Controllers.scala 264:48:@7516.4]
  wire  _T_81; // @[Controllers.scala 264:46:@7517.4]
  wire  _T_82; // @[Controllers.scala 264:62:@7518.4]
  wire  _T_83; // @[Controllers.scala 264:60:@7519.4]
  wire  _T_100; // @[package.scala 100:49:@7536.4]
  reg  _T_103; // @[package.scala 48:56:@7537.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@7550.4 package.scala 96:25:@7551.4]
  wire  _T_110; // @[package.scala 100:49:@7552.4]
  reg  _T_113; // @[package.scala 48:56:@7553.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@7555.4]
  wire  _T_118; // @[Controllers.scala 283:41:@7560.4]
  wire  _T_119; // @[Controllers.scala 283:59:@7561.4]
  wire  _T_121; // @[Controllers.scala 284:37:@7564.4]
  wire  _T_124; // @[package.scala 96:25:@7572.4 package.scala 96:25:@7573.4]
  wire  _T_126; // @[package.scala 100:49:@7574.4]
  reg  _T_129; // @[package.scala 48:56:@7575.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@7597.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@7599.4]
  reg  _T_153; // @[package.scala 48:56:@7600.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@7608.4 package.scala 96:25:@7609.4]
  wire  _T_158; // @[Controllers.scala 292:61:@7610.4]
  wire  _T_159; // @[Controllers.scala 292:24:@7611.4]
  SRFF active ( // @[Controllers.scala 261:22:@7508.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@7511.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_48 RetimeWrapper ( // @[package.scala 93:22:@7545.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_1 ( // @[package.scala 93:22:@7567.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@7579.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@7587.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@7603.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@7516.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@7517.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@7518.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@7519.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@7536.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@7550.4 package.scala 96:25:@7551.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@7552.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@7555.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@7560.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@7561.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@7564.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@7572.4 package.scala 96:25:@7573.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@7574.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@7599.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@7608.4 package.scala 96:25:@7609.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@7610.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@7611.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@7578.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@7613.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@7563.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@7566.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@7558.4]
  assign active_clock = clock; // @[:@7509.4]
  assign active_reset = reset; // @[:@7510.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@7521.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@7525.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@7526.4]
  assign done_clock = clock; // @[:@7512.4]
  assign done_reset = reset; // @[:@7513.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@7541.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@7534.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@7535.4]
  assign RetimeWrapper_clock = clock; // @[:@7546.4]
  assign RetimeWrapper_reset = reset; // @[:@7547.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@7549.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@7548.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7568.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7569.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@7571.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@7570.4]
  assign RetimeWrapper_2_clock = clock; // @[:@7580.4]
  assign RetimeWrapper_2_reset = reset; // @[:@7581.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@7583.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@7582.4]
  assign RetimeWrapper_3_clock = clock; // @[:@7588.4]
  assign RetimeWrapper_3_reset = reset; // @[:@7589.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@7591.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@7590.4]
  assign RetimeWrapper_4_clock = clock; // @[:@7604.4]
  assign RetimeWrapper_4_reset = reset; // @[:@7605.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@7607.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@7606.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_56( // @[:@7804.2]
  input          clock, // @[:@7805.4]
  input          reset, // @[:@7806.4]
  input          io_flow, // @[:@7807.4]
  input  [127:0] io_in, // @[:@7807.4]
  output [127:0] io_out // @[:@7807.4]
);
  wire [127:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire [127:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire [127:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  RetimeShiftRegister #(.WIDTH(128), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7809.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7822.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7821.4]
  assign sr_init = 128'h0; // @[RetimeShiftRegister.scala 19:16:@7820.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7819.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7818.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7816.4]
endmodule
module SRAM_1( // @[:@7840.2]
  input         clock, // @[:@7841.4]
  input         reset, // @[:@7842.4]
  input  [8:0]  io_raddr, // @[:@7843.4]
  input         io_wen, // @[:@7843.4]
  input  [8:0]  io_waddr, // @[:@7843.4]
  input  [31:0] io_wdata, // @[:@7843.4]
  output [31:0] io_rdata, // @[:@7843.4]
  input         io_backpressure // @[:@7843.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@7845.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@7845.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@7845.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@7845.4]
  wire  _T_19; // @[SRAM.scala 182:49:@7863.4]
  wire  _T_20; // @[SRAM.scala 182:37:@7864.4]
  reg  _T_23; // @[SRAM.scala 182:29:@7865.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@7867.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(320), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@7845.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@7863.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@7864.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@7872.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@7859.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@7860.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@7857.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@7862.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@7861.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@7858.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@7856.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@7855.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_57( // @[:@7886.2]
  input        clock, // @[:@7887.4]
  input        reset, // @[:@7888.4]
  input        io_flow, // @[:@7889.4]
  input  [8:0] io_in, // @[:@7889.4]
  output [8:0] io_out // @[:@7889.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7891.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7904.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7903.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@7902.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7901.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7900.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7898.4]
endmodule
module Mem1D_5( // @[:@7906.2]
  input         clock, // @[:@7907.4]
  input         reset, // @[:@7908.4]
  input  [8:0]  io_r_ofs_0, // @[:@7909.4]
  input         io_r_backpressure, // @[:@7909.4]
  input  [8:0]  io_w_ofs_0, // @[:@7909.4]
  input  [31:0] io_w_data_0, // @[:@7909.4]
  input         io_w_en_0, // @[:@7909.4]
  output [31:0] io_output // @[:@7909.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7916.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7916.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7916.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7916.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7916.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@7911.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@7913.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_57 RetimeWrapper ( // @[package.scala 93:22:@7916.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h140; // @[MemPrimitives.scala 702:32:@7911.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@7929.4]
  assign SRAM_clock = clock; // @[:@7914.4]
  assign SRAM_reset = reset; // @[:@7915.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@7923.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@7926.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@7924.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@7927.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@7928.4]
  assign RetimeWrapper_clock = clock; // @[:@7917.4]
  assign RetimeWrapper_reset = reset; // @[:@7918.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@7920.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@7919.4]
endmodule
module StickySelects_1( // @[:@10392.2]
  input   clock, // @[:@10393.4]
  input   reset, // @[:@10394.4]
  input   io_ins_0, // @[:@10395.4]
  input   io_ins_1, // @[:@10395.4]
  input   io_ins_2, // @[:@10395.4]
  input   io_ins_3, // @[:@10395.4]
  input   io_ins_4, // @[:@10395.4]
  input   io_ins_5, // @[:@10395.4]
  input   io_ins_6, // @[:@10395.4]
  input   io_ins_7, // @[:@10395.4]
  input   io_ins_8, // @[:@10395.4]
  output  io_outs_0, // @[:@10395.4]
  output  io_outs_1, // @[:@10395.4]
  output  io_outs_2, // @[:@10395.4]
  output  io_outs_3, // @[:@10395.4]
  output  io_outs_4, // @[:@10395.4]
  output  io_outs_5, // @[:@10395.4]
  output  io_outs_6, // @[:@10395.4]
  output  io_outs_7, // @[:@10395.4]
  output  io_outs_8 // @[:@10395.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@10397.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@10398.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@10399.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@10400.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@10401.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@10402.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@10403.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@10404.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@10405.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@10406.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@10407.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@10408.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@10409.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@10410.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@10411.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@10412.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@10413.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@10414.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@10416.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@10417.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@10418.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@10419.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@10420.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@10421.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@10422.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@10423.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@10424.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@10426.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@10427.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@10428.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@10429.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@10430.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@10431.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@10432.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@10433.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@10434.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@10437.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@10438.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@10439.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@10440.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@10441.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@10442.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@10443.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@10444.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@10448.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@10449.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@10450.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@10451.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@10452.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@10453.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@10454.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@10459.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@10460.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@10461.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@10462.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@10463.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@10464.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@10470.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@10471.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@10472.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@10473.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@10474.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@10481.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@10482.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@10483.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@10484.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@10492.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@10493.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@10494.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@10406.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@10407.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@10408.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@10409.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@10410.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@10411.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@10412.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@10413.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@10414.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@10416.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@10417.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@10418.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@10419.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@10420.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@10421.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@10422.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@10423.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@10424.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@10426.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@10427.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@10428.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@10429.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@10430.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@10431.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@10432.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@10433.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@10434.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@10437.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@10438.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@10439.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@10440.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@10441.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@10442.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@10443.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@10444.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@10448.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@10449.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@10450.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@10451.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@10452.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@10453.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@10454.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@10459.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@10460.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@10461.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@10462.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@10463.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@10464.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@10470.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@10471.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@10472.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@10473.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@10474.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@10481.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@10482.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@10483.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@10484.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@10492.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@10493.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@10494.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@10496.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@10497.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@10498.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@10499.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@10500.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@10501.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@10502.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@10503.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@10504.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x398_lb_0( // @[:@20040.2]
  input         clock, // @[:@20041.4]
  input         reset, // @[:@20042.4]
  input  [2:0]  io_rPort_17_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_17_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_17_ofs_0, // @[:@20043.4]
  input         io_rPort_17_en_0, // @[:@20043.4]
  input         io_rPort_17_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_17_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_16_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_16_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_16_ofs_0, // @[:@20043.4]
  input         io_rPort_16_en_0, // @[:@20043.4]
  input         io_rPort_16_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_16_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_15_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_15_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_15_ofs_0, // @[:@20043.4]
  input         io_rPort_15_en_0, // @[:@20043.4]
  input         io_rPort_15_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_15_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_14_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_14_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_14_ofs_0, // @[:@20043.4]
  input         io_rPort_14_en_0, // @[:@20043.4]
  input         io_rPort_14_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_14_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_13_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_13_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_13_ofs_0, // @[:@20043.4]
  input         io_rPort_13_en_0, // @[:@20043.4]
  input         io_rPort_13_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_13_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_12_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_12_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_12_ofs_0, // @[:@20043.4]
  input         io_rPort_12_en_0, // @[:@20043.4]
  input         io_rPort_12_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_12_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@20043.4]
  input         io_rPort_11_en_0, // @[:@20043.4]
  input         io_rPort_11_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_11_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@20043.4]
  input         io_rPort_10_en_0, // @[:@20043.4]
  input         io_rPort_10_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_10_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@20043.4]
  input         io_rPort_9_en_0, // @[:@20043.4]
  input         io_rPort_9_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_9_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@20043.4]
  input         io_rPort_8_en_0, // @[:@20043.4]
  input         io_rPort_8_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_8_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@20043.4]
  input         io_rPort_7_en_0, // @[:@20043.4]
  input         io_rPort_7_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_7_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@20043.4]
  input         io_rPort_6_en_0, // @[:@20043.4]
  input         io_rPort_6_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_6_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@20043.4]
  input         io_rPort_5_en_0, // @[:@20043.4]
  input         io_rPort_5_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_5_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@20043.4]
  input         io_rPort_4_en_0, // @[:@20043.4]
  input         io_rPort_4_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_4_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@20043.4]
  input         io_rPort_3_en_0, // @[:@20043.4]
  input         io_rPort_3_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_3_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@20043.4]
  input         io_rPort_2_en_0, // @[:@20043.4]
  input         io_rPort_2_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_2_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@20043.4]
  input         io_rPort_1_en_0, // @[:@20043.4]
  input         io_rPort_1_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_1_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@20043.4]
  input         io_rPort_0_en_0, // @[:@20043.4]
  input         io_rPort_0_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_0_output_0, // @[:@20043.4]
  input  [2:0]  io_wPort_3_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_3_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_3_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_3_data_0, // @[:@20043.4]
  input         io_wPort_3_en_0, // @[:@20043.4]
  input  [2:0]  io_wPort_2_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_2_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_2_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_2_data_0, // @[:@20043.4]
  input         io_wPort_2_en_0, // @[:@20043.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_1_data_0, // @[:@20043.4]
  input         io_wPort_1_en_0, // @[:@20043.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_0_data_0, // @[:@20043.4]
  input         io_wPort_0_en_0 // @[:@20043.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_16_clock; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_16_reset; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [8:0] Mem1D_16_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_16_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [8:0] Mem1D_16_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [31:0] Mem1D_16_io_w_data_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_16_io_w_en_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [31:0] Mem1D_16_io_output; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_17_clock; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_17_reset; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [8:0] Mem1D_17_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_17_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [8:0] Mem1D_17_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [31:0] Mem1D_17_io_w_data_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_17_io_w_en_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [31:0] Mem1D_17_io_output; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_18_clock; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_18_reset; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [8:0] Mem1D_18_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_18_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [8:0] Mem1D_18_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [31:0] Mem1D_18_io_w_data_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_18_io_w_en_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [31:0] Mem1D_18_io_output; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_19_clock; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_19_reset; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [8:0] Mem1D_19_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_19_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [8:0] Mem1D_19_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [31:0] Mem1D_19_io_w_data_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_19_io_w_en_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [31:0] Mem1D_19_io_output; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_20_clock; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_20_reset; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [8:0] Mem1D_20_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_20_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [8:0] Mem1D_20_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [31:0] Mem1D_20_io_w_data_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_20_io_w_en_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [31:0] Mem1D_20_io_output; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_21_clock; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_21_reset; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [8:0] Mem1D_21_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_21_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [8:0] Mem1D_21_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [31:0] Mem1D_21_io_w_data_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_21_io_w_en_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [31:0] Mem1D_21_io_output; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_22_clock; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_22_reset; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [8:0] Mem1D_22_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_22_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [8:0] Mem1D_22_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [31:0] Mem1D_22_io_w_data_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_22_io_w_en_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [31:0] Mem1D_22_io_output; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_23_clock; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  Mem1D_23_reset; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [8:0] Mem1D_23_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  Mem1D_23_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [8:0] Mem1D_23_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [31:0] Mem1D_23_io_w_data_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  Mem1D_23_io_w_en_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [31:0] Mem1D_23_io_output; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_6; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_7; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_8; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_6; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_7; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_8; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_6; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_7; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_8; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_6; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_7; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_8; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_8; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_8; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_8; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_8; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_16_clock; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_reset; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_0; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_1; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_2; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_3; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_4; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_5; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_6; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_7; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_8; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_0; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_1; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_2; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_3; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_4; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_5; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_6; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_7; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_8; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_17_clock; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_reset; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_0; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_1; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_2; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_3; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_4; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_5; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_6; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_7; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_8; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_0; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_1; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_2; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_3; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_4; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_5; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_6; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_7; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_8; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_18_clock; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_reset; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_0; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_1; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_2; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_3; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_4; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_5; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_6; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_7; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_8; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_0; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_1; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_2; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_3; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_4; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_5; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_6; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_7; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_8; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_19_clock; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_reset; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_0; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_1; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_2; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_3; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_4; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_5; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_6; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_7; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_8; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_0; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_1; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_2; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_3; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_4; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_5; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_6; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_7; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_8; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_20_clock; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_reset; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_0; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_1; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_2; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_3; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_4; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_5; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_6; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_7; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_8; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_0; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_1; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_2; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_3; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_4; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_5; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_6; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_7; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_8; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_21_clock; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_reset; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_0; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_1; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_2; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_3; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_4; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_5; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_6; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_7; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_8; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_0; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_1; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_2; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_3; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_4; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_5; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_6; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_7; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_8; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_22_clock; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_reset; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_0; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_1; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_2; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_3; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_4; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_5; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_6; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_7; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_8; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_0; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_1; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_2; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_3; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_4; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_5; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_6; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_7; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_8; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_23_clock; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_reset; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_0; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_1; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_2; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_3; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_4; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_5; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_6; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_7; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_8; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_0; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_1; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_2; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_3; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_4; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_5; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_6; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_7; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_8; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_io_in; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_io_out; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_io_in; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_io_out; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_io_in; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_io_out; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_io_in; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_io_out; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_io_in; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_io_out; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_io_in; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_io_out; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_io_in; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_io_out; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_io_in; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_io_out; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_io_in; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_io_out; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_io_in; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_io_out; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_io_in; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_io_out; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_io_in; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_io_out; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_io_in; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_io_out; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_io_in; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_io_out; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_io_in; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_io_out; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_io_in; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_io_out; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_io_in; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_io_out; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_io_in; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_io_out; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_io_in; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_io_out; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_io_in; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_io_out; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_io_in; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_io_out; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_io_in; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_io_out; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_io_in; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_io_out; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_io_in; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_io_out; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_io_in; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_io_out; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_io_in; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_io_out; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_io_in; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_io_out; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_io_in; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_io_out; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_io_in; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_io_out; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_io_in; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_io_out; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_io_in; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_io_out; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_io_in; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_io_out; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_io_in; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_io_out; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_io_in; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_io_out; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_io_in; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_io_out; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_198_clock; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_reset; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_io_flow; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_io_in; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_io_out; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_199_clock; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_reset; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_io_flow; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_io_in; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_io_out; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_200_clock; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_reset; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_io_flow; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_io_in; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_io_out; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_201_clock; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_reset; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_io_flow; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_io_in; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_io_out; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_202_clock; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_reset; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_io_flow; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_io_in; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_io_out; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_203_clock; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_reset; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_io_flow; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_io_in; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_io_out; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_204_clock; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_reset; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_io_flow; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_io_in; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_io_out; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_205_clock; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_reset; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_io_flow; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_io_in; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_io_out; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_206_clock; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_reset; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_io_flow; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_io_in; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_io_out; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_207_clock; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_reset; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_io_flow; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_io_in; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_io_out; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_208_clock; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_reset; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_io_flow; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_io_in; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_io_out; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_209_clock; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_reset; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_io_flow; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_io_in; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_io_out; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_210_clock; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_reset; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_io_flow; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_io_in; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_io_out; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_211_clock; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_reset; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_io_flow; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_io_in; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_io_out; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_212_clock; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_reset; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_io_flow; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_io_in; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_io_out; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_213_clock; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_reset; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_io_flow; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_io_in; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_io_out; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_214_clock; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_reset; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_io_flow; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_io_in; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_io_out; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_215_clock; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_reset; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_io_flow; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_io_in; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_io_out; // @[package.scala 93:22:@25735.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@20570.4]
  wire  _T_702; // @[MemPrimitives.scala 82:210:@20571.4]
  wire  _T_703; // @[MemPrimitives.scala 82:228:@20572.4]
  wire  _T_704; // @[MemPrimitives.scala 83:102:@20573.4]
  wire  _T_706; // @[MemPrimitives.scala 82:210:@20574.4]
  wire  _T_708; // @[MemPrimitives.scala 82:210:@20575.4]
  wire  _T_709; // @[MemPrimitives.scala 82:228:@20576.4]
  wire  _T_710; // @[MemPrimitives.scala 83:102:@20577.4]
  wire [41:0] _T_712; // @[Cat.scala 30:58:@20579.4]
  wire [41:0] _T_714; // @[Cat.scala 30:58:@20581.4]
  wire [41:0] _T_715; // @[Mux.scala 31:69:@20582.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@20589.4]
  wire  _T_722; // @[MemPrimitives.scala 82:210:@20590.4]
  wire  _T_723; // @[MemPrimitives.scala 82:228:@20591.4]
  wire  _T_724; // @[MemPrimitives.scala 83:102:@20592.4]
  wire  _T_726; // @[MemPrimitives.scala 82:210:@20593.4]
  wire  _T_728; // @[MemPrimitives.scala 82:210:@20594.4]
  wire  _T_729; // @[MemPrimitives.scala 82:228:@20595.4]
  wire  _T_730; // @[MemPrimitives.scala 83:102:@20596.4]
  wire [41:0] _T_732; // @[Cat.scala 30:58:@20598.4]
  wire [41:0] _T_734; // @[Cat.scala 30:58:@20600.4]
  wire [41:0] _T_735; // @[Mux.scala 31:69:@20601.4]
  wire  _T_742; // @[MemPrimitives.scala 82:210:@20609.4]
  wire  _T_743; // @[MemPrimitives.scala 82:228:@20610.4]
  wire  _T_744; // @[MemPrimitives.scala 83:102:@20611.4]
  wire  _T_748; // @[MemPrimitives.scala 82:210:@20613.4]
  wire  _T_749; // @[MemPrimitives.scala 82:228:@20614.4]
  wire  _T_750; // @[MemPrimitives.scala 83:102:@20615.4]
  wire [41:0] _T_752; // @[Cat.scala 30:58:@20617.4]
  wire [41:0] _T_754; // @[Cat.scala 30:58:@20619.4]
  wire [41:0] _T_755; // @[Mux.scala 31:69:@20620.4]
  wire  _T_762; // @[MemPrimitives.scala 82:210:@20628.4]
  wire  _T_763; // @[MemPrimitives.scala 82:228:@20629.4]
  wire  _T_764; // @[MemPrimitives.scala 83:102:@20630.4]
  wire  _T_768; // @[MemPrimitives.scala 82:210:@20632.4]
  wire  _T_769; // @[MemPrimitives.scala 82:228:@20633.4]
  wire  _T_770; // @[MemPrimitives.scala 83:102:@20634.4]
  wire [41:0] _T_772; // @[Cat.scala 30:58:@20636.4]
  wire [41:0] _T_774; // @[Cat.scala 30:58:@20638.4]
  wire [41:0] _T_775; // @[Mux.scala 31:69:@20639.4]
  wire  _T_782; // @[MemPrimitives.scala 82:210:@20647.4]
  wire  _T_783; // @[MemPrimitives.scala 82:228:@20648.4]
  wire  _T_784; // @[MemPrimitives.scala 83:102:@20649.4]
  wire  _T_788; // @[MemPrimitives.scala 82:210:@20651.4]
  wire  _T_789; // @[MemPrimitives.scala 82:228:@20652.4]
  wire  _T_790; // @[MemPrimitives.scala 83:102:@20653.4]
  wire [41:0] _T_792; // @[Cat.scala 30:58:@20655.4]
  wire [41:0] _T_794; // @[Cat.scala 30:58:@20657.4]
  wire [41:0] _T_795; // @[Mux.scala 31:69:@20658.4]
  wire  _T_802; // @[MemPrimitives.scala 82:210:@20666.4]
  wire  _T_803; // @[MemPrimitives.scala 82:228:@20667.4]
  wire  _T_804; // @[MemPrimitives.scala 83:102:@20668.4]
  wire  _T_808; // @[MemPrimitives.scala 82:210:@20670.4]
  wire  _T_809; // @[MemPrimitives.scala 82:228:@20671.4]
  wire  _T_810; // @[MemPrimitives.scala 83:102:@20672.4]
  wire [41:0] _T_812; // @[Cat.scala 30:58:@20674.4]
  wire [41:0] _T_814; // @[Cat.scala 30:58:@20676.4]
  wire [41:0] _T_815; // @[Mux.scala 31:69:@20677.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@20684.4]
  wire  _T_823; // @[MemPrimitives.scala 82:228:@20686.4]
  wire  _T_824; // @[MemPrimitives.scala 83:102:@20687.4]
  wire  _T_826; // @[MemPrimitives.scala 82:210:@20688.4]
  wire  _T_829; // @[MemPrimitives.scala 82:228:@20690.4]
  wire  _T_830; // @[MemPrimitives.scala 83:102:@20691.4]
  wire [41:0] _T_832; // @[Cat.scala 30:58:@20693.4]
  wire [41:0] _T_834; // @[Cat.scala 30:58:@20695.4]
  wire [41:0] _T_835; // @[Mux.scala 31:69:@20696.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@20703.4]
  wire  _T_843; // @[MemPrimitives.scala 82:228:@20705.4]
  wire  _T_844; // @[MemPrimitives.scala 83:102:@20706.4]
  wire  _T_846; // @[MemPrimitives.scala 82:210:@20707.4]
  wire  _T_849; // @[MemPrimitives.scala 82:228:@20709.4]
  wire  _T_850; // @[MemPrimitives.scala 83:102:@20710.4]
  wire [41:0] _T_852; // @[Cat.scala 30:58:@20712.4]
  wire [41:0] _T_854; // @[Cat.scala 30:58:@20714.4]
  wire [41:0] _T_855; // @[Mux.scala 31:69:@20715.4]
  wire  _T_863; // @[MemPrimitives.scala 82:228:@20724.4]
  wire  _T_864; // @[MemPrimitives.scala 83:102:@20725.4]
  wire  _T_869; // @[MemPrimitives.scala 82:228:@20728.4]
  wire  _T_870; // @[MemPrimitives.scala 83:102:@20729.4]
  wire [41:0] _T_872; // @[Cat.scala 30:58:@20731.4]
  wire [41:0] _T_874; // @[Cat.scala 30:58:@20733.4]
  wire [41:0] _T_875; // @[Mux.scala 31:69:@20734.4]
  wire  _T_883; // @[MemPrimitives.scala 82:228:@20743.4]
  wire  _T_884; // @[MemPrimitives.scala 83:102:@20744.4]
  wire  _T_889; // @[MemPrimitives.scala 82:228:@20747.4]
  wire  _T_890; // @[MemPrimitives.scala 83:102:@20748.4]
  wire [41:0] _T_892; // @[Cat.scala 30:58:@20750.4]
  wire [41:0] _T_894; // @[Cat.scala 30:58:@20752.4]
  wire [41:0] _T_895; // @[Mux.scala 31:69:@20753.4]
  wire  _T_903; // @[MemPrimitives.scala 82:228:@20762.4]
  wire  _T_904; // @[MemPrimitives.scala 83:102:@20763.4]
  wire  _T_909; // @[MemPrimitives.scala 82:228:@20766.4]
  wire  _T_910; // @[MemPrimitives.scala 83:102:@20767.4]
  wire [41:0] _T_912; // @[Cat.scala 30:58:@20769.4]
  wire [41:0] _T_914; // @[Cat.scala 30:58:@20771.4]
  wire [41:0] _T_915; // @[Mux.scala 31:69:@20772.4]
  wire  _T_923; // @[MemPrimitives.scala 82:228:@20781.4]
  wire  _T_924; // @[MemPrimitives.scala 83:102:@20782.4]
  wire  _T_929; // @[MemPrimitives.scala 82:228:@20785.4]
  wire  _T_930; // @[MemPrimitives.scala 83:102:@20786.4]
  wire [41:0] _T_932; // @[Cat.scala 30:58:@20788.4]
  wire [41:0] _T_934; // @[Cat.scala 30:58:@20790.4]
  wire [41:0] _T_935; // @[Mux.scala 31:69:@20791.4]
  wire  _T_940; // @[MemPrimitives.scala 82:210:@20798.4]
  wire  _T_943; // @[MemPrimitives.scala 82:228:@20800.4]
  wire  _T_944; // @[MemPrimitives.scala 83:102:@20801.4]
  wire  _T_946; // @[MemPrimitives.scala 82:210:@20802.4]
  wire  _T_949; // @[MemPrimitives.scala 82:228:@20804.4]
  wire  _T_950; // @[MemPrimitives.scala 83:102:@20805.4]
  wire [41:0] _T_952; // @[Cat.scala 30:58:@20807.4]
  wire [41:0] _T_954; // @[Cat.scala 30:58:@20809.4]
  wire [41:0] _T_955; // @[Mux.scala 31:69:@20810.4]
  wire  _T_960; // @[MemPrimitives.scala 82:210:@20817.4]
  wire  _T_963; // @[MemPrimitives.scala 82:228:@20819.4]
  wire  _T_964; // @[MemPrimitives.scala 83:102:@20820.4]
  wire  _T_966; // @[MemPrimitives.scala 82:210:@20821.4]
  wire  _T_969; // @[MemPrimitives.scala 82:228:@20823.4]
  wire  _T_970; // @[MemPrimitives.scala 83:102:@20824.4]
  wire [41:0] _T_972; // @[Cat.scala 30:58:@20826.4]
  wire [41:0] _T_974; // @[Cat.scala 30:58:@20828.4]
  wire [41:0] _T_975; // @[Mux.scala 31:69:@20829.4]
  wire  _T_983; // @[MemPrimitives.scala 82:228:@20838.4]
  wire  _T_984; // @[MemPrimitives.scala 83:102:@20839.4]
  wire  _T_989; // @[MemPrimitives.scala 82:228:@20842.4]
  wire  _T_990; // @[MemPrimitives.scala 83:102:@20843.4]
  wire [41:0] _T_992; // @[Cat.scala 30:58:@20845.4]
  wire [41:0] _T_994; // @[Cat.scala 30:58:@20847.4]
  wire [41:0] _T_995; // @[Mux.scala 31:69:@20848.4]
  wire  _T_1003; // @[MemPrimitives.scala 82:228:@20857.4]
  wire  _T_1004; // @[MemPrimitives.scala 83:102:@20858.4]
  wire  _T_1009; // @[MemPrimitives.scala 82:228:@20861.4]
  wire  _T_1010; // @[MemPrimitives.scala 83:102:@20862.4]
  wire [41:0] _T_1012; // @[Cat.scala 30:58:@20864.4]
  wire [41:0] _T_1014; // @[Cat.scala 30:58:@20866.4]
  wire [41:0] _T_1015; // @[Mux.scala 31:69:@20867.4]
  wire  _T_1023; // @[MemPrimitives.scala 82:228:@20876.4]
  wire  _T_1024; // @[MemPrimitives.scala 83:102:@20877.4]
  wire  _T_1029; // @[MemPrimitives.scala 82:228:@20880.4]
  wire  _T_1030; // @[MemPrimitives.scala 83:102:@20881.4]
  wire [41:0] _T_1032; // @[Cat.scala 30:58:@20883.4]
  wire [41:0] _T_1034; // @[Cat.scala 30:58:@20885.4]
  wire [41:0] _T_1035; // @[Mux.scala 31:69:@20886.4]
  wire  _T_1043; // @[MemPrimitives.scala 82:228:@20895.4]
  wire  _T_1044; // @[MemPrimitives.scala 83:102:@20896.4]
  wire  _T_1049; // @[MemPrimitives.scala 82:228:@20899.4]
  wire  _T_1050; // @[MemPrimitives.scala 83:102:@20900.4]
  wire [41:0] _T_1052; // @[Cat.scala 30:58:@20902.4]
  wire [41:0] _T_1054; // @[Cat.scala 30:58:@20904.4]
  wire [41:0] _T_1055; // @[Mux.scala 31:69:@20905.4]
  wire  _T_1060; // @[MemPrimitives.scala 82:210:@20912.4]
  wire  _T_1063; // @[MemPrimitives.scala 82:228:@20914.4]
  wire  _T_1064; // @[MemPrimitives.scala 83:102:@20915.4]
  wire  _T_1066; // @[MemPrimitives.scala 82:210:@20916.4]
  wire  _T_1069; // @[MemPrimitives.scala 82:228:@20918.4]
  wire  _T_1070; // @[MemPrimitives.scala 83:102:@20919.4]
  wire [41:0] _T_1072; // @[Cat.scala 30:58:@20921.4]
  wire [41:0] _T_1074; // @[Cat.scala 30:58:@20923.4]
  wire [41:0] _T_1075; // @[Mux.scala 31:69:@20924.4]
  wire  _T_1080; // @[MemPrimitives.scala 82:210:@20931.4]
  wire  _T_1083; // @[MemPrimitives.scala 82:228:@20933.4]
  wire  _T_1084; // @[MemPrimitives.scala 83:102:@20934.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@20935.4]
  wire  _T_1089; // @[MemPrimitives.scala 82:228:@20937.4]
  wire  _T_1090; // @[MemPrimitives.scala 83:102:@20938.4]
  wire [41:0] _T_1092; // @[Cat.scala 30:58:@20940.4]
  wire [41:0] _T_1094; // @[Cat.scala 30:58:@20942.4]
  wire [41:0] _T_1095; // @[Mux.scala 31:69:@20943.4]
  wire  _T_1103; // @[MemPrimitives.scala 82:228:@20952.4]
  wire  _T_1104; // @[MemPrimitives.scala 83:102:@20953.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:228:@20956.4]
  wire  _T_1110; // @[MemPrimitives.scala 83:102:@20957.4]
  wire [41:0] _T_1112; // @[Cat.scala 30:58:@20959.4]
  wire [41:0] _T_1114; // @[Cat.scala 30:58:@20961.4]
  wire [41:0] _T_1115; // @[Mux.scala 31:69:@20962.4]
  wire  _T_1123; // @[MemPrimitives.scala 82:228:@20971.4]
  wire  _T_1124; // @[MemPrimitives.scala 83:102:@20972.4]
  wire  _T_1129; // @[MemPrimitives.scala 82:228:@20975.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@20976.4]
  wire [41:0] _T_1132; // @[Cat.scala 30:58:@20978.4]
  wire [41:0] _T_1134; // @[Cat.scala 30:58:@20980.4]
  wire [41:0] _T_1135; // @[Mux.scala 31:69:@20981.4]
  wire  _T_1143; // @[MemPrimitives.scala 82:228:@20990.4]
  wire  _T_1144; // @[MemPrimitives.scala 83:102:@20991.4]
  wire  _T_1149; // @[MemPrimitives.scala 82:228:@20994.4]
  wire  _T_1150; // @[MemPrimitives.scala 83:102:@20995.4]
  wire [41:0] _T_1152; // @[Cat.scala 30:58:@20997.4]
  wire [41:0] _T_1154; // @[Cat.scala 30:58:@20999.4]
  wire [41:0] _T_1155; // @[Mux.scala 31:69:@21000.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:228:@21009.4]
  wire  _T_1164; // @[MemPrimitives.scala 83:102:@21010.4]
  wire  _T_1169; // @[MemPrimitives.scala 82:228:@21013.4]
  wire  _T_1170; // @[MemPrimitives.scala 83:102:@21014.4]
  wire [41:0] _T_1172; // @[Cat.scala 30:58:@21016.4]
  wire [41:0] _T_1174; // @[Cat.scala 30:58:@21018.4]
  wire [41:0] _T_1175; // @[Mux.scala 31:69:@21019.4]
  wire  _T_1180; // @[MemPrimitives.scala 110:210:@21026.4]
  wire  _T_1182; // @[MemPrimitives.scala 110:210:@21027.4]
  wire  _T_1183; // @[MemPrimitives.scala 110:228:@21028.4]
  wire  _T_1186; // @[MemPrimitives.scala 110:210:@21030.4]
  wire  _T_1188; // @[MemPrimitives.scala 110:210:@21031.4]
  wire  _T_1189; // @[MemPrimitives.scala 110:228:@21032.4]
  wire  _T_1192; // @[MemPrimitives.scala 110:210:@21034.4]
  wire  _T_1194; // @[MemPrimitives.scala 110:210:@21035.4]
  wire  _T_1195; // @[MemPrimitives.scala 110:228:@21036.4]
  wire  _T_1198; // @[MemPrimitives.scala 110:210:@21038.4]
  wire  _T_1200; // @[MemPrimitives.scala 110:210:@21039.4]
  wire  _T_1201; // @[MemPrimitives.scala 110:228:@21040.4]
  wire  _T_1204; // @[MemPrimitives.scala 110:210:@21042.4]
  wire  _T_1206; // @[MemPrimitives.scala 110:210:@21043.4]
  wire  _T_1207; // @[MemPrimitives.scala 110:228:@21044.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@21046.4]
  wire  _T_1212; // @[MemPrimitives.scala 110:210:@21047.4]
  wire  _T_1213; // @[MemPrimitives.scala 110:228:@21048.4]
  wire  _T_1216; // @[MemPrimitives.scala 110:210:@21050.4]
  wire  _T_1218; // @[MemPrimitives.scala 110:210:@21051.4]
  wire  _T_1219; // @[MemPrimitives.scala 110:228:@21052.4]
  wire  _T_1222; // @[MemPrimitives.scala 110:210:@21054.4]
  wire  _T_1224; // @[MemPrimitives.scala 110:210:@21055.4]
  wire  _T_1225; // @[MemPrimitives.scala 110:228:@21056.4]
  wire  _T_1228; // @[MemPrimitives.scala 110:210:@21058.4]
  wire  _T_1230; // @[MemPrimitives.scala 110:210:@21059.4]
  wire  _T_1231; // @[MemPrimitives.scala 110:228:@21060.4]
  wire  _T_1233; // @[MemPrimitives.scala 126:35:@21074.4]
  wire  _T_1234; // @[MemPrimitives.scala 126:35:@21075.4]
  wire  _T_1235; // @[MemPrimitives.scala 126:35:@21076.4]
  wire  _T_1236; // @[MemPrimitives.scala 126:35:@21077.4]
  wire  _T_1237; // @[MemPrimitives.scala 126:35:@21078.4]
  wire  _T_1238; // @[MemPrimitives.scala 126:35:@21079.4]
  wire  _T_1239; // @[MemPrimitives.scala 126:35:@21080.4]
  wire  _T_1240; // @[MemPrimitives.scala 126:35:@21081.4]
  wire  _T_1241; // @[MemPrimitives.scala 126:35:@21082.4]
  wire [10:0] _T_1243; // @[Cat.scala 30:58:@21084.4]
  wire [10:0] _T_1245; // @[Cat.scala 30:58:@21086.4]
  wire [10:0] _T_1247; // @[Cat.scala 30:58:@21088.4]
  wire [10:0] _T_1249; // @[Cat.scala 30:58:@21090.4]
  wire [10:0] _T_1251; // @[Cat.scala 30:58:@21092.4]
  wire [10:0] _T_1253; // @[Cat.scala 30:58:@21094.4]
  wire [10:0] _T_1255; // @[Cat.scala 30:58:@21096.4]
  wire [10:0] _T_1257; // @[Cat.scala 30:58:@21098.4]
  wire [10:0] _T_1259; // @[Cat.scala 30:58:@21100.4]
  wire [10:0] _T_1260; // @[Mux.scala 31:69:@21101.4]
  wire [10:0] _T_1261; // @[Mux.scala 31:69:@21102.4]
  wire [10:0] _T_1262; // @[Mux.scala 31:69:@21103.4]
  wire [10:0] _T_1263; // @[Mux.scala 31:69:@21104.4]
  wire [10:0] _T_1264; // @[Mux.scala 31:69:@21105.4]
  wire [10:0] _T_1265; // @[Mux.scala 31:69:@21106.4]
  wire [10:0] _T_1266; // @[Mux.scala 31:69:@21107.4]
  wire [10:0] _T_1267; // @[Mux.scala 31:69:@21108.4]
  wire  _T_1272; // @[MemPrimitives.scala 110:210:@21115.4]
  wire  _T_1274; // @[MemPrimitives.scala 110:210:@21116.4]
  wire  _T_1275; // @[MemPrimitives.scala 110:228:@21117.4]
  wire  _T_1278; // @[MemPrimitives.scala 110:210:@21119.4]
  wire  _T_1280; // @[MemPrimitives.scala 110:210:@21120.4]
  wire  _T_1281; // @[MemPrimitives.scala 110:228:@21121.4]
  wire  _T_1284; // @[MemPrimitives.scala 110:210:@21123.4]
  wire  _T_1286; // @[MemPrimitives.scala 110:210:@21124.4]
  wire  _T_1287; // @[MemPrimitives.scala 110:228:@21125.4]
  wire  _T_1290; // @[MemPrimitives.scala 110:210:@21127.4]
  wire  _T_1292; // @[MemPrimitives.scala 110:210:@21128.4]
  wire  _T_1293; // @[MemPrimitives.scala 110:228:@21129.4]
  wire  _T_1296; // @[MemPrimitives.scala 110:210:@21131.4]
  wire  _T_1298; // @[MemPrimitives.scala 110:210:@21132.4]
  wire  _T_1299; // @[MemPrimitives.scala 110:228:@21133.4]
  wire  _T_1302; // @[MemPrimitives.scala 110:210:@21135.4]
  wire  _T_1304; // @[MemPrimitives.scala 110:210:@21136.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@21137.4]
  wire  _T_1308; // @[MemPrimitives.scala 110:210:@21139.4]
  wire  _T_1310; // @[MemPrimitives.scala 110:210:@21140.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@21141.4]
  wire  _T_1314; // @[MemPrimitives.scala 110:210:@21143.4]
  wire  _T_1316; // @[MemPrimitives.scala 110:210:@21144.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@21145.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@21147.4]
  wire  _T_1322; // @[MemPrimitives.scala 110:210:@21148.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@21149.4]
  wire  _T_1325; // @[MemPrimitives.scala 126:35:@21163.4]
  wire  _T_1326; // @[MemPrimitives.scala 126:35:@21164.4]
  wire  _T_1327; // @[MemPrimitives.scala 126:35:@21165.4]
  wire  _T_1328; // @[MemPrimitives.scala 126:35:@21166.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@21167.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@21168.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@21169.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@21170.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@21171.4]
  wire [10:0] _T_1335; // @[Cat.scala 30:58:@21173.4]
  wire [10:0] _T_1337; // @[Cat.scala 30:58:@21175.4]
  wire [10:0] _T_1339; // @[Cat.scala 30:58:@21177.4]
  wire [10:0] _T_1341; // @[Cat.scala 30:58:@21179.4]
  wire [10:0] _T_1343; // @[Cat.scala 30:58:@21181.4]
  wire [10:0] _T_1345; // @[Cat.scala 30:58:@21183.4]
  wire [10:0] _T_1347; // @[Cat.scala 30:58:@21185.4]
  wire [10:0] _T_1349; // @[Cat.scala 30:58:@21187.4]
  wire [10:0] _T_1351; // @[Cat.scala 30:58:@21189.4]
  wire [10:0] _T_1352; // @[Mux.scala 31:69:@21190.4]
  wire [10:0] _T_1353; // @[Mux.scala 31:69:@21191.4]
  wire [10:0] _T_1354; // @[Mux.scala 31:69:@21192.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@21193.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@21194.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@21195.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@21196.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@21197.4]
  wire  _T_1366; // @[MemPrimitives.scala 110:210:@21205.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@21206.4]
  wire  _T_1372; // @[MemPrimitives.scala 110:210:@21209.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@21210.4]
  wire  _T_1378; // @[MemPrimitives.scala 110:210:@21213.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@21214.4]
  wire  _T_1384; // @[MemPrimitives.scala 110:210:@21217.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@21218.4]
  wire  _T_1390; // @[MemPrimitives.scala 110:210:@21221.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@21222.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@21225.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@21226.4]
  wire  _T_1402; // @[MemPrimitives.scala 110:210:@21229.4]
  wire  _T_1403; // @[MemPrimitives.scala 110:228:@21230.4]
  wire  _T_1408; // @[MemPrimitives.scala 110:210:@21233.4]
  wire  _T_1409; // @[MemPrimitives.scala 110:228:@21234.4]
  wire  _T_1414; // @[MemPrimitives.scala 110:210:@21237.4]
  wire  _T_1415; // @[MemPrimitives.scala 110:228:@21238.4]
  wire  _T_1417; // @[MemPrimitives.scala 126:35:@21252.4]
  wire  _T_1418; // @[MemPrimitives.scala 126:35:@21253.4]
  wire  _T_1419; // @[MemPrimitives.scala 126:35:@21254.4]
  wire  _T_1420; // @[MemPrimitives.scala 126:35:@21255.4]
  wire  _T_1421; // @[MemPrimitives.scala 126:35:@21256.4]
  wire  _T_1422; // @[MemPrimitives.scala 126:35:@21257.4]
  wire  _T_1423; // @[MemPrimitives.scala 126:35:@21258.4]
  wire  _T_1424; // @[MemPrimitives.scala 126:35:@21259.4]
  wire  _T_1425; // @[MemPrimitives.scala 126:35:@21260.4]
  wire [10:0] _T_1427; // @[Cat.scala 30:58:@21262.4]
  wire [10:0] _T_1429; // @[Cat.scala 30:58:@21264.4]
  wire [10:0] _T_1431; // @[Cat.scala 30:58:@21266.4]
  wire [10:0] _T_1433; // @[Cat.scala 30:58:@21268.4]
  wire [10:0] _T_1435; // @[Cat.scala 30:58:@21270.4]
  wire [10:0] _T_1437; // @[Cat.scala 30:58:@21272.4]
  wire [10:0] _T_1439; // @[Cat.scala 30:58:@21274.4]
  wire [10:0] _T_1441; // @[Cat.scala 30:58:@21276.4]
  wire [10:0] _T_1443; // @[Cat.scala 30:58:@21278.4]
  wire [10:0] _T_1444; // @[Mux.scala 31:69:@21279.4]
  wire [10:0] _T_1445; // @[Mux.scala 31:69:@21280.4]
  wire [10:0] _T_1446; // @[Mux.scala 31:69:@21281.4]
  wire [10:0] _T_1447; // @[Mux.scala 31:69:@21282.4]
  wire [10:0] _T_1448; // @[Mux.scala 31:69:@21283.4]
  wire [10:0] _T_1449; // @[Mux.scala 31:69:@21284.4]
  wire [10:0] _T_1450; // @[Mux.scala 31:69:@21285.4]
  wire [10:0] _T_1451; // @[Mux.scala 31:69:@21286.4]
  wire  _T_1458; // @[MemPrimitives.scala 110:210:@21294.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@21295.4]
  wire  _T_1464; // @[MemPrimitives.scala 110:210:@21298.4]
  wire  _T_1465; // @[MemPrimitives.scala 110:228:@21299.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@21302.4]
  wire  _T_1471; // @[MemPrimitives.scala 110:228:@21303.4]
  wire  _T_1476; // @[MemPrimitives.scala 110:210:@21306.4]
  wire  _T_1477; // @[MemPrimitives.scala 110:228:@21307.4]
  wire  _T_1482; // @[MemPrimitives.scala 110:210:@21310.4]
  wire  _T_1483; // @[MemPrimitives.scala 110:228:@21311.4]
  wire  _T_1488; // @[MemPrimitives.scala 110:210:@21314.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:228:@21315.4]
  wire  _T_1494; // @[MemPrimitives.scala 110:210:@21318.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:228:@21319.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@21322.4]
  wire  _T_1501; // @[MemPrimitives.scala 110:228:@21323.4]
  wire  _T_1506; // @[MemPrimitives.scala 110:210:@21326.4]
  wire  _T_1507; // @[MemPrimitives.scala 110:228:@21327.4]
  wire  _T_1509; // @[MemPrimitives.scala 126:35:@21341.4]
  wire  _T_1510; // @[MemPrimitives.scala 126:35:@21342.4]
  wire  _T_1511; // @[MemPrimitives.scala 126:35:@21343.4]
  wire  _T_1512; // @[MemPrimitives.scala 126:35:@21344.4]
  wire  _T_1513; // @[MemPrimitives.scala 126:35:@21345.4]
  wire  _T_1514; // @[MemPrimitives.scala 126:35:@21346.4]
  wire  _T_1515; // @[MemPrimitives.scala 126:35:@21347.4]
  wire  _T_1516; // @[MemPrimitives.scala 126:35:@21348.4]
  wire  _T_1517; // @[MemPrimitives.scala 126:35:@21349.4]
  wire [10:0] _T_1519; // @[Cat.scala 30:58:@21351.4]
  wire [10:0] _T_1521; // @[Cat.scala 30:58:@21353.4]
  wire [10:0] _T_1523; // @[Cat.scala 30:58:@21355.4]
  wire [10:0] _T_1525; // @[Cat.scala 30:58:@21357.4]
  wire [10:0] _T_1527; // @[Cat.scala 30:58:@21359.4]
  wire [10:0] _T_1529; // @[Cat.scala 30:58:@21361.4]
  wire [10:0] _T_1531; // @[Cat.scala 30:58:@21363.4]
  wire [10:0] _T_1533; // @[Cat.scala 30:58:@21365.4]
  wire [10:0] _T_1535; // @[Cat.scala 30:58:@21367.4]
  wire [10:0] _T_1536; // @[Mux.scala 31:69:@21368.4]
  wire [10:0] _T_1537; // @[Mux.scala 31:69:@21369.4]
  wire [10:0] _T_1538; // @[Mux.scala 31:69:@21370.4]
  wire [10:0] _T_1539; // @[Mux.scala 31:69:@21371.4]
  wire [10:0] _T_1540; // @[Mux.scala 31:69:@21372.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@21373.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@21374.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@21375.4]
  wire  _T_1550; // @[MemPrimitives.scala 110:210:@21383.4]
  wire  _T_1551; // @[MemPrimitives.scala 110:228:@21384.4]
  wire  _T_1556; // @[MemPrimitives.scala 110:210:@21387.4]
  wire  _T_1557; // @[MemPrimitives.scala 110:228:@21388.4]
  wire  _T_1562; // @[MemPrimitives.scala 110:210:@21391.4]
  wire  _T_1563; // @[MemPrimitives.scala 110:228:@21392.4]
  wire  _T_1568; // @[MemPrimitives.scala 110:210:@21395.4]
  wire  _T_1569; // @[MemPrimitives.scala 110:228:@21396.4]
  wire  _T_1574; // @[MemPrimitives.scala 110:210:@21399.4]
  wire  _T_1575; // @[MemPrimitives.scala 110:228:@21400.4]
  wire  _T_1580; // @[MemPrimitives.scala 110:210:@21403.4]
  wire  _T_1581; // @[MemPrimitives.scala 110:228:@21404.4]
  wire  _T_1586; // @[MemPrimitives.scala 110:210:@21407.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:228:@21408.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@21411.4]
  wire  _T_1593; // @[MemPrimitives.scala 110:228:@21412.4]
  wire  _T_1598; // @[MemPrimitives.scala 110:210:@21415.4]
  wire  _T_1599; // @[MemPrimitives.scala 110:228:@21416.4]
  wire  _T_1601; // @[MemPrimitives.scala 126:35:@21430.4]
  wire  _T_1602; // @[MemPrimitives.scala 126:35:@21431.4]
  wire  _T_1603; // @[MemPrimitives.scala 126:35:@21432.4]
  wire  _T_1604; // @[MemPrimitives.scala 126:35:@21433.4]
  wire  _T_1605; // @[MemPrimitives.scala 126:35:@21434.4]
  wire  _T_1606; // @[MemPrimitives.scala 126:35:@21435.4]
  wire  _T_1607; // @[MemPrimitives.scala 126:35:@21436.4]
  wire  _T_1608; // @[MemPrimitives.scala 126:35:@21437.4]
  wire  _T_1609; // @[MemPrimitives.scala 126:35:@21438.4]
  wire [10:0] _T_1611; // @[Cat.scala 30:58:@21440.4]
  wire [10:0] _T_1613; // @[Cat.scala 30:58:@21442.4]
  wire [10:0] _T_1615; // @[Cat.scala 30:58:@21444.4]
  wire [10:0] _T_1617; // @[Cat.scala 30:58:@21446.4]
  wire [10:0] _T_1619; // @[Cat.scala 30:58:@21448.4]
  wire [10:0] _T_1621; // @[Cat.scala 30:58:@21450.4]
  wire [10:0] _T_1623; // @[Cat.scala 30:58:@21452.4]
  wire [10:0] _T_1625; // @[Cat.scala 30:58:@21454.4]
  wire [10:0] _T_1627; // @[Cat.scala 30:58:@21456.4]
  wire [10:0] _T_1628; // @[Mux.scala 31:69:@21457.4]
  wire [10:0] _T_1629; // @[Mux.scala 31:69:@21458.4]
  wire [10:0] _T_1630; // @[Mux.scala 31:69:@21459.4]
  wire [10:0] _T_1631; // @[Mux.scala 31:69:@21460.4]
  wire [10:0] _T_1632; // @[Mux.scala 31:69:@21461.4]
  wire [10:0] _T_1633; // @[Mux.scala 31:69:@21462.4]
  wire [10:0] _T_1634; // @[Mux.scala 31:69:@21463.4]
  wire [10:0] _T_1635; // @[Mux.scala 31:69:@21464.4]
  wire  _T_1642; // @[MemPrimitives.scala 110:210:@21472.4]
  wire  _T_1643; // @[MemPrimitives.scala 110:228:@21473.4]
  wire  _T_1648; // @[MemPrimitives.scala 110:210:@21476.4]
  wire  _T_1649; // @[MemPrimitives.scala 110:228:@21477.4]
  wire  _T_1654; // @[MemPrimitives.scala 110:210:@21480.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:228:@21481.4]
  wire  _T_1660; // @[MemPrimitives.scala 110:210:@21484.4]
  wire  _T_1661; // @[MemPrimitives.scala 110:228:@21485.4]
  wire  _T_1666; // @[MemPrimitives.scala 110:210:@21488.4]
  wire  _T_1667; // @[MemPrimitives.scala 110:228:@21489.4]
  wire  _T_1672; // @[MemPrimitives.scala 110:210:@21492.4]
  wire  _T_1673; // @[MemPrimitives.scala 110:228:@21493.4]
  wire  _T_1678; // @[MemPrimitives.scala 110:210:@21496.4]
  wire  _T_1679; // @[MemPrimitives.scala 110:228:@21497.4]
  wire  _T_1684; // @[MemPrimitives.scala 110:210:@21500.4]
  wire  _T_1685; // @[MemPrimitives.scala 110:228:@21501.4]
  wire  _T_1690; // @[MemPrimitives.scala 110:210:@21504.4]
  wire  _T_1691; // @[MemPrimitives.scala 110:228:@21505.4]
  wire  _T_1693; // @[MemPrimitives.scala 126:35:@21519.4]
  wire  _T_1694; // @[MemPrimitives.scala 126:35:@21520.4]
  wire  _T_1695; // @[MemPrimitives.scala 126:35:@21521.4]
  wire  _T_1696; // @[MemPrimitives.scala 126:35:@21522.4]
  wire  _T_1697; // @[MemPrimitives.scala 126:35:@21523.4]
  wire  _T_1698; // @[MemPrimitives.scala 126:35:@21524.4]
  wire  _T_1699; // @[MemPrimitives.scala 126:35:@21525.4]
  wire  _T_1700; // @[MemPrimitives.scala 126:35:@21526.4]
  wire  _T_1701; // @[MemPrimitives.scala 126:35:@21527.4]
  wire [10:0] _T_1703; // @[Cat.scala 30:58:@21529.4]
  wire [10:0] _T_1705; // @[Cat.scala 30:58:@21531.4]
  wire [10:0] _T_1707; // @[Cat.scala 30:58:@21533.4]
  wire [10:0] _T_1709; // @[Cat.scala 30:58:@21535.4]
  wire [10:0] _T_1711; // @[Cat.scala 30:58:@21537.4]
  wire [10:0] _T_1713; // @[Cat.scala 30:58:@21539.4]
  wire [10:0] _T_1715; // @[Cat.scala 30:58:@21541.4]
  wire [10:0] _T_1717; // @[Cat.scala 30:58:@21543.4]
  wire [10:0] _T_1719; // @[Cat.scala 30:58:@21545.4]
  wire [10:0] _T_1720; // @[Mux.scala 31:69:@21546.4]
  wire [10:0] _T_1721; // @[Mux.scala 31:69:@21547.4]
  wire [10:0] _T_1722; // @[Mux.scala 31:69:@21548.4]
  wire [10:0] _T_1723; // @[Mux.scala 31:69:@21549.4]
  wire [10:0] _T_1724; // @[Mux.scala 31:69:@21550.4]
  wire [10:0] _T_1725; // @[Mux.scala 31:69:@21551.4]
  wire [10:0] _T_1726; // @[Mux.scala 31:69:@21552.4]
  wire [10:0] _T_1727; // @[Mux.scala 31:69:@21553.4]
  wire  _T_1732; // @[MemPrimitives.scala 110:210:@21560.4]
  wire  _T_1735; // @[MemPrimitives.scala 110:228:@21562.4]
  wire  _T_1738; // @[MemPrimitives.scala 110:210:@21564.4]
  wire  _T_1741; // @[MemPrimitives.scala 110:228:@21566.4]
  wire  _T_1744; // @[MemPrimitives.scala 110:210:@21568.4]
  wire  _T_1747; // @[MemPrimitives.scala 110:228:@21570.4]
  wire  _T_1750; // @[MemPrimitives.scala 110:210:@21572.4]
  wire  _T_1753; // @[MemPrimitives.scala 110:228:@21574.4]
  wire  _T_1756; // @[MemPrimitives.scala 110:210:@21576.4]
  wire  _T_1759; // @[MemPrimitives.scala 110:228:@21578.4]
  wire  _T_1762; // @[MemPrimitives.scala 110:210:@21580.4]
  wire  _T_1765; // @[MemPrimitives.scala 110:228:@21582.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@21584.4]
  wire  _T_1771; // @[MemPrimitives.scala 110:228:@21586.4]
  wire  _T_1774; // @[MemPrimitives.scala 110:210:@21588.4]
  wire  _T_1777; // @[MemPrimitives.scala 110:228:@21590.4]
  wire  _T_1780; // @[MemPrimitives.scala 110:210:@21592.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:228:@21594.4]
  wire  _T_1785; // @[MemPrimitives.scala 126:35:@21608.4]
  wire  _T_1786; // @[MemPrimitives.scala 126:35:@21609.4]
  wire  _T_1787; // @[MemPrimitives.scala 126:35:@21610.4]
  wire  _T_1788; // @[MemPrimitives.scala 126:35:@21611.4]
  wire  _T_1789; // @[MemPrimitives.scala 126:35:@21612.4]
  wire  _T_1790; // @[MemPrimitives.scala 126:35:@21613.4]
  wire  _T_1791; // @[MemPrimitives.scala 126:35:@21614.4]
  wire  _T_1792; // @[MemPrimitives.scala 126:35:@21615.4]
  wire  _T_1793; // @[MemPrimitives.scala 126:35:@21616.4]
  wire [10:0] _T_1795; // @[Cat.scala 30:58:@21618.4]
  wire [10:0] _T_1797; // @[Cat.scala 30:58:@21620.4]
  wire [10:0] _T_1799; // @[Cat.scala 30:58:@21622.4]
  wire [10:0] _T_1801; // @[Cat.scala 30:58:@21624.4]
  wire [10:0] _T_1803; // @[Cat.scala 30:58:@21626.4]
  wire [10:0] _T_1805; // @[Cat.scala 30:58:@21628.4]
  wire [10:0] _T_1807; // @[Cat.scala 30:58:@21630.4]
  wire [10:0] _T_1809; // @[Cat.scala 30:58:@21632.4]
  wire [10:0] _T_1811; // @[Cat.scala 30:58:@21634.4]
  wire [10:0] _T_1812; // @[Mux.scala 31:69:@21635.4]
  wire [10:0] _T_1813; // @[Mux.scala 31:69:@21636.4]
  wire [10:0] _T_1814; // @[Mux.scala 31:69:@21637.4]
  wire [10:0] _T_1815; // @[Mux.scala 31:69:@21638.4]
  wire [10:0] _T_1816; // @[Mux.scala 31:69:@21639.4]
  wire [10:0] _T_1817; // @[Mux.scala 31:69:@21640.4]
  wire [10:0] _T_1818; // @[Mux.scala 31:69:@21641.4]
  wire [10:0] _T_1819; // @[Mux.scala 31:69:@21642.4]
  wire  _T_1824; // @[MemPrimitives.scala 110:210:@21649.4]
  wire  _T_1827; // @[MemPrimitives.scala 110:228:@21651.4]
  wire  _T_1830; // @[MemPrimitives.scala 110:210:@21653.4]
  wire  _T_1833; // @[MemPrimitives.scala 110:228:@21655.4]
  wire  _T_1836; // @[MemPrimitives.scala 110:210:@21657.4]
  wire  _T_1839; // @[MemPrimitives.scala 110:228:@21659.4]
  wire  _T_1842; // @[MemPrimitives.scala 110:210:@21661.4]
  wire  _T_1845; // @[MemPrimitives.scala 110:228:@21663.4]
  wire  _T_1848; // @[MemPrimitives.scala 110:210:@21665.4]
  wire  _T_1851; // @[MemPrimitives.scala 110:228:@21667.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@21669.4]
  wire  _T_1857; // @[MemPrimitives.scala 110:228:@21671.4]
  wire  _T_1860; // @[MemPrimitives.scala 110:210:@21673.4]
  wire  _T_1863; // @[MemPrimitives.scala 110:228:@21675.4]
  wire  _T_1866; // @[MemPrimitives.scala 110:210:@21677.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:228:@21679.4]
  wire  _T_1872; // @[MemPrimitives.scala 110:210:@21681.4]
  wire  _T_1875; // @[MemPrimitives.scala 110:228:@21683.4]
  wire  _T_1877; // @[MemPrimitives.scala 126:35:@21697.4]
  wire  _T_1878; // @[MemPrimitives.scala 126:35:@21698.4]
  wire  _T_1879; // @[MemPrimitives.scala 126:35:@21699.4]
  wire  _T_1880; // @[MemPrimitives.scala 126:35:@21700.4]
  wire  _T_1881; // @[MemPrimitives.scala 126:35:@21701.4]
  wire  _T_1882; // @[MemPrimitives.scala 126:35:@21702.4]
  wire  _T_1883; // @[MemPrimitives.scala 126:35:@21703.4]
  wire  _T_1884; // @[MemPrimitives.scala 126:35:@21704.4]
  wire  _T_1885; // @[MemPrimitives.scala 126:35:@21705.4]
  wire [10:0] _T_1887; // @[Cat.scala 30:58:@21707.4]
  wire [10:0] _T_1889; // @[Cat.scala 30:58:@21709.4]
  wire [10:0] _T_1891; // @[Cat.scala 30:58:@21711.4]
  wire [10:0] _T_1893; // @[Cat.scala 30:58:@21713.4]
  wire [10:0] _T_1895; // @[Cat.scala 30:58:@21715.4]
  wire [10:0] _T_1897; // @[Cat.scala 30:58:@21717.4]
  wire [10:0] _T_1899; // @[Cat.scala 30:58:@21719.4]
  wire [10:0] _T_1901; // @[Cat.scala 30:58:@21721.4]
  wire [10:0] _T_1903; // @[Cat.scala 30:58:@21723.4]
  wire [10:0] _T_1904; // @[Mux.scala 31:69:@21724.4]
  wire [10:0] _T_1905; // @[Mux.scala 31:69:@21725.4]
  wire [10:0] _T_1906; // @[Mux.scala 31:69:@21726.4]
  wire [10:0] _T_1907; // @[Mux.scala 31:69:@21727.4]
  wire [10:0] _T_1908; // @[Mux.scala 31:69:@21728.4]
  wire [10:0] _T_1909; // @[Mux.scala 31:69:@21729.4]
  wire [10:0] _T_1910; // @[Mux.scala 31:69:@21730.4]
  wire [10:0] _T_1911; // @[Mux.scala 31:69:@21731.4]
  wire  _T_1919; // @[MemPrimitives.scala 110:228:@21740.4]
  wire  _T_1925; // @[MemPrimitives.scala 110:228:@21744.4]
  wire  _T_1931; // @[MemPrimitives.scala 110:228:@21748.4]
  wire  _T_1937; // @[MemPrimitives.scala 110:228:@21752.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:228:@21756.4]
  wire  _T_1949; // @[MemPrimitives.scala 110:228:@21760.4]
  wire  _T_1955; // @[MemPrimitives.scala 110:228:@21764.4]
  wire  _T_1961; // @[MemPrimitives.scala 110:228:@21768.4]
  wire  _T_1967; // @[MemPrimitives.scala 110:228:@21772.4]
  wire  _T_1969; // @[MemPrimitives.scala 126:35:@21786.4]
  wire  _T_1970; // @[MemPrimitives.scala 126:35:@21787.4]
  wire  _T_1971; // @[MemPrimitives.scala 126:35:@21788.4]
  wire  _T_1972; // @[MemPrimitives.scala 126:35:@21789.4]
  wire  _T_1973; // @[MemPrimitives.scala 126:35:@21790.4]
  wire  _T_1974; // @[MemPrimitives.scala 126:35:@21791.4]
  wire  _T_1975; // @[MemPrimitives.scala 126:35:@21792.4]
  wire  _T_1976; // @[MemPrimitives.scala 126:35:@21793.4]
  wire  _T_1977; // @[MemPrimitives.scala 126:35:@21794.4]
  wire [10:0] _T_1979; // @[Cat.scala 30:58:@21796.4]
  wire [10:0] _T_1981; // @[Cat.scala 30:58:@21798.4]
  wire [10:0] _T_1983; // @[Cat.scala 30:58:@21800.4]
  wire [10:0] _T_1985; // @[Cat.scala 30:58:@21802.4]
  wire [10:0] _T_1987; // @[Cat.scala 30:58:@21804.4]
  wire [10:0] _T_1989; // @[Cat.scala 30:58:@21806.4]
  wire [10:0] _T_1991; // @[Cat.scala 30:58:@21808.4]
  wire [10:0] _T_1993; // @[Cat.scala 30:58:@21810.4]
  wire [10:0] _T_1995; // @[Cat.scala 30:58:@21812.4]
  wire [10:0] _T_1996; // @[Mux.scala 31:69:@21813.4]
  wire [10:0] _T_1997; // @[Mux.scala 31:69:@21814.4]
  wire [10:0] _T_1998; // @[Mux.scala 31:69:@21815.4]
  wire [10:0] _T_1999; // @[Mux.scala 31:69:@21816.4]
  wire [10:0] _T_2000; // @[Mux.scala 31:69:@21817.4]
  wire [10:0] _T_2001; // @[Mux.scala 31:69:@21818.4]
  wire [10:0] _T_2002; // @[Mux.scala 31:69:@21819.4]
  wire [10:0] _T_2003; // @[Mux.scala 31:69:@21820.4]
  wire  _T_2011; // @[MemPrimitives.scala 110:228:@21829.4]
  wire  _T_2017; // @[MemPrimitives.scala 110:228:@21833.4]
  wire  _T_2023; // @[MemPrimitives.scala 110:228:@21837.4]
  wire  _T_2029; // @[MemPrimitives.scala 110:228:@21841.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:228:@21845.4]
  wire  _T_2041; // @[MemPrimitives.scala 110:228:@21849.4]
  wire  _T_2047; // @[MemPrimitives.scala 110:228:@21853.4]
  wire  _T_2053; // @[MemPrimitives.scala 110:228:@21857.4]
  wire  _T_2059; // @[MemPrimitives.scala 110:228:@21861.4]
  wire  _T_2061; // @[MemPrimitives.scala 126:35:@21875.4]
  wire  _T_2062; // @[MemPrimitives.scala 126:35:@21876.4]
  wire  _T_2063; // @[MemPrimitives.scala 126:35:@21877.4]
  wire  _T_2064; // @[MemPrimitives.scala 126:35:@21878.4]
  wire  _T_2065; // @[MemPrimitives.scala 126:35:@21879.4]
  wire  _T_2066; // @[MemPrimitives.scala 126:35:@21880.4]
  wire  _T_2067; // @[MemPrimitives.scala 126:35:@21881.4]
  wire  _T_2068; // @[MemPrimitives.scala 126:35:@21882.4]
  wire  _T_2069; // @[MemPrimitives.scala 126:35:@21883.4]
  wire [10:0] _T_2071; // @[Cat.scala 30:58:@21885.4]
  wire [10:0] _T_2073; // @[Cat.scala 30:58:@21887.4]
  wire [10:0] _T_2075; // @[Cat.scala 30:58:@21889.4]
  wire [10:0] _T_2077; // @[Cat.scala 30:58:@21891.4]
  wire [10:0] _T_2079; // @[Cat.scala 30:58:@21893.4]
  wire [10:0] _T_2081; // @[Cat.scala 30:58:@21895.4]
  wire [10:0] _T_2083; // @[Cat.scala 30:58:@21897.4]
  wire [10:0] _T_2085; // @[Cat.scala 30:58:@21899.4]
  wire [10:0] _T_2087; // @[Cat.scala 30:58:@21901.4]
  wire [10:0] _T_2088; // @[Mux.scala 31:69:@21902.4]
  wire [10:0] _T_2089; // @[Mux.scala 31:69:@21903.4]
  wire [10:0] _T_2090; // @[Mux.scala 31:69:@21904.4]
  wire [10:0] _T_2091; // @[Mux.scala 31:69:@21905.4]
  wire [10:0] _T_2092; // @[Mux.scala 31:69:@21906.4]
  wire [10:0] _T_2093; // @[Mux.scala 31:69:@21907.4]
  wire [10:0] _T_2094; // @[Mux.scala 31:69:@21908.4]
  wire [10:0] _T_2095; // @[Mux.scala 31:69:@21909.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:228:@21918.4]
  wire  _T_2109; // @[MemPrimitives.scala 110:228:@21922.4]
  wire  _T_2115; // @[MemPrimitives.scala 110:228:@21926.4]
  wire  _T_2121; // @[MemPrimitives.scala 110:228:@21930.4]
  wire  _T_2127; // @[MemPrimitives.scala 110:228:@21934.4]
  wire  _T_2133; // @[MemPrimitives.scala 110:228:@21938.4]
  wire  _T_2139; // @[MemPrimitives.scala 110:228:@21942.4]
  wire  _T_2145; // @[MemPrimitives.scala 110:228:@21946.4]
  wire  _T_2151; // @[MemPrimitives.scala 110:228:@21950.4]
  wire  _T_2153; // @[MemPrimitives.scala 126:35:@21964.4]
  wire  _T_2154; // @[MemPrimitives.scala 126:35:@21965.4]
  wire  _T_2155; // @[MemPrimitives.scala 126:35:@21966.4]
  wire  _T_2156; // @[MemPrimitives.scala 126:35:@21967.4]
  wire  _T_2157; // @[MemPrimitives.scala 126:35:@21968.4]
  wire  _T_2158; // @[MemPrimitives.scala 126:35:@21969.4]
  wire  _T_2159; // @[MemPrimitives.scala 126:35:@21970.4]
  wire  _T_2160; // @[MemPrimitives.scala 126:35:@21971.4]
  wire  _T_2161; // @[MemPrimitives.scala 126:35:@21972.4]
  wire [10:0] _T_2163; // @[Cat.scala 30:58:@21974.4]
  wire [10:0] _T_2165; // @[Cat.scala 30:58:@21976.4]
  wire [10:0] _T_2167; // @[Cat.scala 30:58:@21978.4]
  wire [10:0] _T_2169; // @[Cat.scala 30:58:@21980.4]
  wire [10:0] _T_2171; // @[Cat.scala 30:58:@21982.4]
  wire [10:0] _T_2173; // @[Cat.scala 30:58:@21984.4]
  wire [10:0] _T_2175; // @[Cat.scala 30:58:@21986.4]
  wire [10:0] _T_2177; // @[Cat.scala 30:58:@21988.4]
  wire [10:0] _T_2179; // @[Cat.scala 30:58:@21990.4]
  wire [10:0] _T_2180; // @[Mux.scala 31:69:@21991.4]
  wire [10:0] _T_2181; // @[Mux.scala 31:69:@21992.4]
  wire [10:0] _T_2182; // @[Mux.scala 31:69:@21993.4]
  wire [10:0] _T_2183; // @[Mux.scala 31:69:@21994.4]
  wire [10:0] _T_2184; // @[Mux.scala 31:69:@21995.4]
  wire [10:0] _T_2185; // @[Mux.scala 31:69:@21996.4]
  wire [10:0] _T_2186; // @[Mux.scala 31:69:@21997.4]
  wire [10:0] _T_2187; // @[Mux.scala 31:69:@21998.4]
  wire  _T_2195; // @[MemPrimitives.scala 110:228:@22007.4]
  wire  _T_2201; // @[MemPrimitives.scala 110:228:@22011.4]
  wire  _T_2207; // @[MemPrimitives.scala 110:228:@22015.4]
  wire  _T_2213; // @[MemPrimitives.scala 110:228:@22019.4]
  wire  _T_2219; // @[MemPrimitives.scala 110:228:@22023.4]
  wire  _T_2225; // @[MemPrimitives.scala 110:228:@22027.4]
  wire  _T_2231; // @[MemPrimitives.scala 110:228:@22031.4]
  wire  _T_2237; // @[MemPrimitives.scala 110:228:@22035.4]
  wire  _T_2243; // @[MemPrimitives.scala 110:228:@22039.4]
  wire  _T_2245; // @[MemPrimitives.scala 126:35:@22053.4]
  wire  _T_2246; // @[MemPrimitives.scala 126:35:@22054.4]
  wire  _T_2247; // @[MemPrimitives.scala 126:35:@22055.4]
  wire  _T_2248; // @[MemPrimitives.scala 126:35:@22056.4]
  wire  _T_2249; // @[MemPrimitives.scala 126:35:@22057.4]
  wire  _T_2250; // @[MemPrimitives.scala 126:35:@22058.4]
  wire  _T_2251; // @[MemPrimitives.scala 126:35:@22059.4]
  wire  _T_2252; // @[MemPrimitives.scala 126:35:@22060.4]
  wire  _T_2253; // @[MemPrimitives.scala 126:35:@22061.4]
  wire [10:0] _T_2255; // @[Cat.scala 30:58:@22063.4]
  wire [10:0] _T_2257; // @[Cat.scala 30:58:@22065.4]
  wire [10:0] _T_2259; // @[Cat.scala 30:58:@22067.4]
  wire [10:0] _T_2261; // @[Cat.scala 30:58:@22069.4]
  wire [10:0] _T_2263; // @[Cat.scala 30:58:@22071.4]
  wire [10:0] _T_2265; // @[Cat.scala 30:58:@22073.4]
  wire [10:0] _T_2267; // @[Cat.scala 30:58:@22075.4]
  wire [10:0] _T_2269; // @[Cat.scala 30:58:@22077.4]
  wire [10:0] _T_2271; // @[Cat.scala 30:58:@22079.4]
  wire [10:0] _T_2272; // @[Mux.scala 31:69:@22080.4]
  wire [10:0] _T_2273; // @[Mux.scala 31:69:@22081.4]
  wire [10:0] _T_2274; // @[Mux.scala 31:69:@22082.4]
  wire [10:0] _T_2275; // @[Mux.scala 31:69:@22083.4]
  wire [10:0] _T_2276; // @[Mux.scala 31:69:@22084.4]
  wire [10:0] _T_2277; // @[Mux.scala 31:69:@22085.4]
  wire [10:0] _T_2278; // @[Mux.scala 31:69:@22086.4]
  wire [10:0] _T_2279; // @[Mux.scala 31:69:@22087.4]
  wire  _T_2284; // @[MemPrimitives.scala 110:210:@22094.4]
  wire  _T_2287; // @[MemPrimitives.scala 110:228:@22096.4]
  wire  _T_2290; // @[MemPrimitives.scala 110:210:@22098.4]
  wire  _T_2293; // @[MemPrimitives.scala 110:228:@22100.4]
  wire  _T_2296; // @[MemPrimitives.scala 110:210:@22102.4]
  wire  _T_2299; // @[MemPrimitives.scala 110:228:@22104.4]
  wire  _T_2302; // @[MemPrimitives.scala 110:210:@22106.4]
  wire  _T_2305; // @[MemPrimitives.scala 110:228:@22108.4]
  wire  _T_2308; // @[MemPrimitives.scala 110:210:@22110.4]
  wire  _T_2311; // @[MemPrimitives.scala 110:228:@22112.4]
  wire  _T_2314; // @[MemPrimitives.scala 110:210:@22114.4]
  wire  _T_2317; // @[MemPrimitives.scala 110:228:@22116.4]
  wire  _T_2320; // @[MemPrimitives.scala 110:210:@22118.4]
  wire  _T_2323; // @[MemPrimitives.scala 110:228:@22120.4]
  wire  _T_2326; // @[MemPrimitives.scala 110:210:@22122.4]
  wire  _T_2329; // @[MemPrimitives.scala 110:228:@22124.4]
  wire  _T_2332; // @[MemPrimitives.scala 110:210:@22126.4]
  wire  _T_2335; // @[MemPrimitives.scala 110:228:@22128.4]
  wire  _T_2337; // @[MemPrimitives.scala 126:35:@22142.4]
  wire  _T_2338; // @[MemPrimitives.scala 126:35:@22143.4]
  wire  _T_2339; // @[MemPrimitives.scala 126:35:@22144.4]
  wire  _T_2340; // @[MemPrimitives.scala 126:35:@22145.4]
  wire  _T_2341; // @[MemPrimitives.scala 126:35:@22146.4]
  wire  _T_2342; // @[MemPrimitives.scala 126:35:@22147.4]
  wire  _T_2343; // @[MemPrimitives.scala 126:35:@22148.4]
  wire  _T_2344; // @[MemPrimitives.scala 126:35:@22149.4]
  wire  _T_2345; // @[MemPrimitives.scala 126:35:@22150.4]
  wire [10:0] _T_2347; // @[Cat.scala 30:58:@22152.4]
  wire [10:0] _T_2349; // @[Cat.scala 30:58:@22154.4]
  wire [10:0] _T_2351; // @[Cat.scala 30:58:@22156.4]
  wire [10:0] _T_2353; // @[Cat.scala 30:58:@22158.4]
  wire [10:0] _T_2355; // @[Cat.scala 30:58:@22160.4]
  wire [10:0] _T_2357; // @[Cat.scala 30:58:@22162.4]
  wire [10:0] _T_2359; // @[Cat.scala 30:58:@22164.4]
  wire [10:0] _T_2361; // @[Cat.scala 30:58:@22166.4]
  wire [10:0] _T_2363; // @[Cat.scala 30:58:@22168.4]
  wire [10:0] _T_2364; // @[Mux.scala 31:69:@22169.4]
  wire [10:0] _T_2365; // @[Mux.scala 31:69:@22170.4]
  wire [10:0] _T_2366; // @[Mux.scala 31:69:@22171.4]
  wire [10:0] _T_2367; // @[Mux.scala 31:69:@22172.4]
  wire [10:0] _T_2368; // @[Mux.scala 31:69:@22173.4]
  wire [10:0] _T_2369; // @[Mux.scala 31:69:@22174.4]
  wire [10:0] _T_2370; // @[Mux.scala 31:69:@22175.4]
  wire [10:0] _T_2371; // @[Mux.scala 31:69:@22176.4]
  wire  _T_2376; // @[MemPrimitives.scala 110:210:@22183.4]
  wire  _T_2379; // @[MemPrimitives.scala 110:228:@22185.4]
  wire  _T_2382; // @[MemPrimitives.scala 110:210:@22187.4]
  wire  _T_2385; // @[MemPrimitives.scala 110:228:@22189.4]
  wire  _T_2388; // @[MemPrimitives.scala 110:210:@22191.4]
  wire  _T_2391; // @[MemPrimitives.scala 110:228:@22193.4]
  wire  _T_2394; // @[MemPrimitives.scala 110:210:@22195.4]
  wire  _T_2397; // @[MemPrimitives.scala 110:228:@22197.4]
  wire  _T_2400; // @[MemPrimitives.scala 110:210:@22199.4]
  wire  _T_2403; // @[MemPrimitives.scala 110:228:@22201.4]
  wire  _T_2406; // @[MemPrimitives.scala 110:210:@22203.4]
  wire  _T_2409; // @[MemPrimitives.scala 110:228:@22205.4]
  wire  _T_2412; // @[MemPrimitives.scala 110:210:@22207.4]
  wire  _T_2415; // @[MemPrimitives.scala 110:228:@22209.4]
  wire  _T_2418; // @[MemPrimitives.scala 110:210:@22211.4]
  wire  _T_2421; // @[MemPrimitives.scala 110:228:@22213.4]
  wire  _T_2424; // @[MemPrimitives.scala 110:210:@22215.4]
  wire  _T_2427; // @[MemPrimitives.scala 110:228:@22217.4]
  wire  _T_2429; // @[MemPrimitives.scala 126:35:@22231.4]
  wire  _T_2430; // @[MemPrimitives.scala 126:35:@22232.4]
  wire  _T_2431; // @[MemPrimitives.scala 126:35:@22233.4]
  wire  _T_2432; // @[MemPrimitives.scala 126:35:@22234.4]
  wire  _T_2433; // @[MemPrimitives.scala 126:35:@22235.4]
  wire  _T_2434; // @[MemPrimitives.scala 126:35:@22236.4]
  wire  _T_2435; // @[MemPrimitives.scala 126:35:@22237.4]
  wire  _T_2436; // @[MemPrimitives.scala 126:35:@22238.4]
  wire  _T_2437; // @[MemPrimitives.scala 126:35:@22239.4]
  wire [10:0] _T_2439; // @[Cat.scala 30:58:@22241.4]
  wire [10:0] _T_2441; // @[Cat.scala 30:58:@22243.4]
  wire [10:0] _T_2443; // @[Cat.scala 30:58:@22245.4]
  wire [10:0] _T_2445; // @[Cat.scala 30:58:@22247.4]
  wire [10:0] _T_2447; // @[Cat.scala 30:58:@22249.4]
  wire [10:0] _T_2449; // @[Cat.scala 30:58:@22251.4]
  wire [10:0] _T_2451; // @[Cat.scala 30:58:@22253.4]
  wire [10:0] _T_2453; // @[Cat.scala 30:58:@22255.4]
  wire [10:0] _T_2455; // @[Cat.scala 30:58:@22257.4]
  wire [10:0] _T_2456; // @[Mux.scala 31:69:@22258.4]
  wire [10:0] _T_2457; // @[Mux.scala 31:69:@22259.4]
  wire [10:0] _T_2458; // @[Mux.scala 31:69:@22260.4]
  wire [10:0] _T_2459; // @[Mux.scala 31:69:@22261.4]
  wire [10:0] _T_2460; // @[Mux.scala 31:69:@22262.4]
  wire [10:0] _T_2461; // @[Mux.scala 31:69:@22263.4]
  wire [10:0] _T_2462; // @[Mux.scala 31:69:@22264.4]
  wire [10:0] _T_2463; // @[Mux.scala 31:69:@22265.4]
  wire  _T_2471; // @[MemPrimitives.scala 110:228:@22274.4]
  wire  _T_2477; // @[MemPrimitives.scala 110:228:@22278.4]
  wire  _T_2483; // @[MemPrimitives.scala 110:228:@22282.4]
  wire  _T_2489; // @[MemPrimitives.scala 110:228:@22286.4]
  wire  _T_2495; // @[MemPrimitives.scala 110:228:@22290.4]
  wire  _T_2501; // @[MemPrimitives.scala 110:228:@22294.4]
  wire  _T_2507; // @[MemPrimitives.scala 110:228:@22298.4]
  wire  _T_2513; // @[MemPrimitives.scala 110:228:@22302.4]
  wire  _T_2519; // @[MemPrimitives.scala 110:228:@22306.4]
  wire  _T_2521; // @[MemPrimitives.scala 126:35:@22320.4]
  wire  _T_2522; // @[MemPrimitives.scala 126:35:@22321.4]
  wire  _T_2523; // @[MemPrimitives.scala 126:35:@22322.4]
  wire  _T_2524; // @[MemPrimitives.scala 126:35:@22323.4]
  wire  _T_2525; // @[MemPrimitives.scala 126:35:@22324.4]
  wire  _T_2526; // @[MemPrimitives.scala 126:35:@22325.4]
  wire  _T_2527; // @[MemPrimitives.scala 126:35:@22326.4]
  wire  _T_2528; // @[MemPrimitives.scala 126:35:@22327.4]
  wire  _T_2529; // @[MemPrimitives.scala 126:35:@22328.4]
  wire [10:0] _T_2531; // @[Cat.scala 30:58:@22330.4]
  wire [10:0] _T_2533; // @[Cat.scala 30:58:@22332.4]
  wire [10:0] _T_2535; // @[Cat.scala 30:58:@22334.4]
  wire [10:0] _T_2537; // @[Cat.scala 30:58:@22336.4]
  wire [10:0] _T_2539; // @[Cat.scala 30:58:@22338.4]
  wire [10:0] _T_2541; // @[Cat.scala 30:58:@22340.4]
  wire [10:0] _T_2543; // @[Cat.scala 30:58:@22342.4]
  wire [10:0] _T_2545; // @[Cat.scala 30:58:@22344.4]
  wire [10:0] _T_2547; // @[Cat.scala 30:58:@22346.4]
  wire [10:0] _T_2548; // @[Mux.scala 31:69:@22347.4]
  wire [10:0] _T_2549; // @[Mux.scala 31:69:@22348.4]
  wire [10:0] _T_2550; // @[Mux.scala 31:69:@22349.4]
  wire [10:0] _T_2551; // @[Mux.scala 31:69:@22350.4]
  wire [10:0] _T_2552; // @[Mux.scala 31:69:@22351.4]
  wire [10:0] _T_2553; // @[Mux.scala 31:69:@22352.4]
  wire [10:0] _T_2554; // @[Mux.scala 31:69:@22353.4]
  wire [10:0] _T_2555; // @[Mux.scala 31:69:@22354.4]
  wire  _T_2563; // @[MemPrimitives.scala 110:228:@22363.4]
  wire  _T_2569; // @[MemPrimitives.scala 110:228:@22367.4]
  wire  _T_2575; // @[MemPrimitives.scala 110:228:@22371.4]
  wire  _T_2581; // @[MemPrimitives.scala 110:228:@22375.4]
  wire  _T_2587; // @[MemPrimitives.scala 110:228:@22379.4]
  wire  _T_2593; // @[MemPrimitives.scala 110:228:@22383.4]
  wire  _T_2599; // @[MemPrimitives.scala 110:228:@22387.4]
  wire  _T_2605; // @[MemPrimitives.scala 110:228:@22391.4]
  wire  _T_2611; // @[MemPrimitives.scala 110:228:@22395.4]
  wire  _T_2613; // @[MemPrimitives.scala 126:35:@22409.4]
  wire  _T_2614; // @[MemPrimitives.scala 126:35:@22410.4]
  wire  _T_2615; // @[MemPrimitives.scala 126:35:@22411.4]
  wire  _T_2616; // @[MemPrimitives.scala 126:35:@22412.4]
  wire  _T_2617; // @[MemPrimitives.scala 126:35:@22413.4]
  wire  _T_2618; // @[MemPrimitives.scala 126:35:@22414.4]
  wire  _T_2619; // @[MemPrimitives.scala 126:35:@22415.4]
  wire  _T_2620; // @[MemPrimitives.scala 126:35:@22416.4]
  wire  _T_2621; // @[MemPrimitives.scala 126:35:@22417.4]
  wire [10:0] _T_2623; // @[Cat.scala 30:58:@22419.4]
  wire [10:0] _T_2625; // @[Cat.scala 30:58:@22421.4]
  wire [10:0] _T_2627; // @[Cat.scala 30:58:@22423.4]
  wire [10:0] _T_2629; // @[Cat.scala 30:58:@22425.4]
  wire [10:0] _T_2631; // @[Cat.scala 30:58:@22427.4]
  wire [10:0] _T_2633; // @[Cat.scala 30:58:@22429.4]
  wire [10:0] _T_2635; // @[Cat.scala 30:58:@22431.4]
  wire [10:0] _T_2637; // @[Cat.scala 30:58:@22433.4]
  wire [10:0] _T_2639; // @[Cat.scala 30:58:@22435.4]
  wire [10:0] _T_2640; // @[Mux.scala 31:69:@22436.4]
  wire [10:0] _T_2641; // @[Mux.scala 31:69:@22437.4]
  wire [10:0] _T_2642; // @[Mux.scala 31:69:@22438.4]
  wire [10:0] _T_2643; // @[Mux.scala 31:69:@22439.4]
  wire [10:0] _T_2644; // @[Mux.scala 31:69:@22440.4]
  wire [10:0] _T_2645; // @[Mux.scala 31:69:@22441.4]
  wire [10:0] _T_2646; // @[Mux.scala 31:69:@22442.4]
  wire [10:0] _T_2647; // @[Mux.scala 31:69:@22443.4]
  wire  _T_2655; // @[MemPrimitives.scala 110:228:@22452.4]
  wire  _T_2661; // @[MemPrimitives.scala 110:228:@22456.4]
  wire  _T_2667; // @[MemPrimitives.scala 110:228:@22460.4]
  wire  _T_2673; // @[MemPrimitives.scala 110:228:@22464.4]
  wire  _T_2679; // @[MemPrimitives.scala 110:228:@22468.4]
  wire  _T_2685; // @[MemPrimitives.scala 110:228:@22472.4]
  wire  _T_2691; // @[MemPrimitives.scala 110:228:@22476.4]
  wire  _T_2697; // @[MemPrimitives.scala 110:228:@22480.4]
  wire  _T_2703; // @[MemPrimitives.scala 110:228:@22484.4]
  wire  _T_2705; // @[MemPrimitives.scala 126:35:@22498.4]
  wire  _T_2706; // @[MemPrimitives.scala 126:35:@22499.4]
  wire  _T_2707; // @[MemPrimitives.scala 126:35:@22500.4]
  wire  _T_2708; // @[MemPrimitives.scala 126:35:@22501.4]
  wire  _T_2709; // @[MemPrimitives.scala 126:35:@22502.4]
  wire  _T_2710; // @[MemPrimitives.scala 126:35:@22503.4]
  wire  _T_2711; // @[MemPrimitives.scala 126:35:@22504.4]
  wire  _T_2712; // @[MemPrimitives.scala 126:35:@22505.4]
  wire  _T_2713; // @[MemPrimitives.scala 126:35:@22506.4]
  wire [10:0] _T_2715; // @[Cat.scala 30:58:@22508.4]
  wire [10:0] _T_2717; // @[Cat.scala 30:58:@22510.4]
  wire [10:0] _T_2719; // @[Cat.scala 30:58:@22512.4]
  wire [10:0] _T_2721; // @[Cat.scala 30:58:@22514.4]
  wire [10:0] _T_2723; // @[Cat.scala 30:58:@22516.4]
  wire [10:0] _T_2725; // @[Cat.scala 30:58:@22518.4]
  wire [10:0] _T_2727; // @[Cat.scala 30:58:@22520.4]
  wire [10:0] _T_2729; // @[Cat.scala 30:58:@22522.4]
  wire [10:0] _T_2731; // @[Cat.scala 30:58:@22524.4]
  wire [10:0] _T_2732; // @[Mux.scala 31:69:@22525.4]
  wire [10:0] _T_2733; // @[Mux.scala 31:69:@22526.4]
  wire [10:0] _T_2734; // @[Mux.scala 31:69:@22527.4]
  wire [10:0] _T_2735; // @[Mux.scala 31:69:@22528.4]
  wire [10:0] _T_2736; // @[Mux.scala 31:69:@22529.4]
  wire [10:0] _T_2737; // @[Mux.scala 31:69:@22530.4]
  wire [10:0] _T_2738; // @[Mux.scala 31:69:@22531.4]
  wire [10:0] _T_2739; // @[Mux.scala 31:69:@22532.4]
  wire  _T_2747; // @[MemPrimitives.scala 110:228:@22541.4]
  wire  _T_2753; // @[MemPrimitives.scala 110:228:@22545.4]
  wire  _T_2759; // @[MemPrimitives.scala 110:228:@22549.4]
  wire  _T_2765; // @[MemPrimitives.scala 110:228:@22553.4]
  wire  _T_2771; // @[MemPrimitives.scala 110:228:@22557.4]
  wire  _T_2777; // @[MemPrimitives.scala 110:228:@22561.4]
  wire  _T_2783; // @[MemPrimitives.scala 110:228:@22565.4]
  wire  _T_2789; // @[MemPrimitives.scala 110:228:@22569.4]
  wire  _T_2795; // @[MemPrimitives.scala 110:228:@22573.4]
  wire  _T_2797; // @[MemPrimitives.scala 126:35:@22587.4]
  wire  _T_2798; // @[MemPrimitives.scala 126:35:@22588.4]
  wire  _T_2799; // @[MemPrimitives.scala 126:35:@22589.4]
  wire  _T_2800; // @[MemPrimitives.scala 126:35:@22590.4]
  wire  _T_2801; // @[MemPrimitives.scala 126:35:@22591.4]
  wire  _T_2802; // @[MemPrimitives.scala 126:35:@22592.4]
  wire  _T_2803; // @[MemPrimitives.scala 126:35:@22593.4]
  wire  _T_2804; // @[MemPrimitives.scala 126:35:@22594.4]
  wire  _T_2805; // @[MemPrimitives.scala 126:35:@22595.4]
  wire [10:0] _T_2807; // @[Cat.scala 30:58:@22597.4]
  wire [10:0] _T_2809; // @[Cat.scala 30:58:@22599.4]
  wire [10:0] _T_2811; // @[Cat.scala 30:58:@22601.4]
  wire [10:0] _T_2813; // @[Cat.scala 30:58:@22603.4]
  wire [10:0] _T_2815; // @[Cat.scala 30:58:@22605.4]
  wire [10:0] _T_2817; // @[Cat.scala 30:58:@22607.4]
  wire [10:0] _T_2819; // @[Cat.scala 30:58:@22609.4]
  wire [10:0] _T_2821; // @[Cat.scala 30:58:@22611.4]
  wire [10:0] _T_2823; // @[Cat.scala 30:58:@22613.4]
  wire [10:0] _T_2824; // @[Mux.scala 31:69:@22614.4]
  wire [10:0] _T_2825; // @[Mux.scala 31:69:@22615.4]
  wire [10:0] _T_2826; // @[Mux.scala 31:69:@22616.4]
  wire [10:0] _T_2827; // @[Mux.scala 31:69:@22617.4]
  wire [10:0] _T_2828; // @[Mux.scala 31:69:@22618.4]
  wire [10:0] _T_2829; // @[Mux.scala 31:69:@22619.4]
  wire [10:0] _T_2830; // @[Mux.scala 31:69:@22620.4]
  wire [10:0] _T_2831; // @[Mux.scala 31:69:@22621.4]
  wire  _T_2836; // @[MemPrimitives.scala 110:210:@22628.4]
  wire  _T_2839; // @[MemPrimitives.scala 110:228:@22630.4]
  wire  _T_2842; // @[MemPrimitives.scala 110:210:@22632.4]
  wire  _T_2845; // @[MemPrimitives.scala 110:228:@22634.4]
  wire  _T_2848; // @[MemPrimitives.scala 110:210:@22636.4]
  wire  _T_2851; // @[MemPrimitives.scala 110:228:@22638.4]
  wire  _T_2854; // @[MemPrimitives.scala 110:210:@22640.4]
  wire  _T_2857; // @[MemPrimitives.scala 110:228:@22642.4]
  wire  _T_2860; // @[MemPrimitives.scala 110:210:@22644.4]
  wire  _T_2863; // @[MemPrimitives.scala 110:228:@22646.4]
  wire  _T_2866; // @[MemPrimitives.scala 110:210:@22648.4]
  wire  _T_2869; // @[MemPrimitives.scala 110:228:@22650.4]
  wire  _T_2872; // @[MemPrimitives.scala 110:210:@22652.4]
  wire  _T_2875; // @[MemPrimitives.scala 110:228:@22654.4]
  wire  _T_2878; // @[MemPrimitives.scala 110:210:@22656.4]
  wire  _T_2881; // @[MemPrimitives.scala 110:228:@22658.4]
  wire  _T_2884; // @[MemPrimitives.scala 110:210:@22660.4]
  wire  _T_2887; // @[MemPrimitives.scala 110:228:@22662.4]
  wire  _T_2889; // @[MemPrimitives.scala 126:35:@22676.4]
  wire  _T_2890; // @[MemPrimitives.scala 126:35:@22677.4]
  wire  _T_2891; // @[MemPrimitives.scala 126:35:@22678.4]
  wire  _T_2892; // @[MemPrimitives.scala 126:35:@22679.4]
  wire  _T_2893; // @[MemPrimitives.scala 126:35:@22680.4]
  wire  _T_2894; // @[MemPrimitives.scala 126:35:@22681.4]
  wire  _T_2895; // @[MemPrimitives.scala 126:35:@22682.4]
  wire  _T_2896; // @[MemPrimitives.scala 126:35:@22683.4]
  wire  _T_2897; // @[MemPrimitives.scala 126:35:@22684.4]
  wire [10:0] _T_2899; // @[Cat.scala 30:58:@22686.4]
  wire [10:0] _T_2901; // @[Cat.scala 30:58:@22688.4]
  wire [10:0] _T_2903; // @[Cat.scala 30:58:@22690.4]
  wire [10:0] _T_2905; // @[Cat.scala 30:58:@22692.4]
  wire [10:0] _T_2907; // @[Cat.scala 30:58:@22694.4]
  wire [10:0] _T_2909; // @[Cat.scala 30:58:@22696.4]
  wire [10:0] _T_2911; // @[Cat.scala 30:58:@22698.4]
  wire [10:0] _T_2913; // @[Cat.scala 30:58:@22700.4]
  wire [10:0] _T_2915; // @[Cat.scala 30:58:@22702.4]
  wire [10:0] _T_2916; // @[Mux.scala 31:69:@22703.4]
  wire [10:0] _T_2917; // @[Mux.scala 31:69:@22704.4]
  wire [10:0] _T_2918; // @[Mux.scala 31:69:@22705.4]
  wire [10:0] _T_2919; // @[Mux.scala 31:69:@22706.4]
  wire [10:0] _T_2920; // @[Mux.scala 31:69:@22707.4]
  wire [10:0] _T_2921; // @[Mux.scala 31:69:@22708.4]
  wire [10:0] _T_2922; // @[Mux.scala 31:69:@22709.4]
  wire [10:0] _T_2923; // @[Mux.scala 31:69:@22710.4]
  wire  _T_2928; // @[MemPrimitives.scala 110:210:@22717.4]
  wire  _T_2931; // @[MemPrimitives.scala 110:228:@22719.4]
  wire  _T_2934; // @[MemPrimitives.scala 110:210:@22721.4]
  wire  _T_2937; // @[MemPrimitives.scala 110:228:@22723.4]
  wire  _T_2940; // @[MemPrimitives.scala 110:210:@22725.4]
  wire  _T_2943; // @[MemPrimitives.scala 110:228:@22727.4]
  wire  _T_2946; // @[MemPrimitives.scala 110:210:@22729.4]
  wire  _T_2949; // @[MemPrimitives.scala 110:228:@22731.4]
  wire  _T_2952; // @[MemPrimitives.scala 110:210:@22733.4]
  wire  _T_2955; // @[MemPrimitives.scala 110:228:@22735.4]
  wire  _T_2958; // @[MemPrimitives.scala 110:210:@22737.4]
  wire  _T_2961; // @[MemPrimitives.scala 110:228:@22739.4]
  wire  _T_2964; // @[MemPrimitives.scala 110:210:@22741.4]
  wire  _T_2967; // @[MemPrimitives.scala 110:228:@22743.4]
  wire  _T_2970; // @[MemPrimitives.scala 110:210:@22745.4]
  wire  _T_2973; // @[MemPrimitives.scala 110:228:@22747.4]
  wire  _T_2976; // @[MemPrimitives.scala 110:210:@22749.4]
  wire  _T_2979; // @[MemPrimitives.scala 110:228:@22751.4]
  wire  _T_2981; // @[MemPrimitives.scala 126:35:@22765.4]
  wire  _T_2982; // @[MemPrimitives.scala 126:35:@22766.4]
  wire  _T_2983; // @[MemPrimitives.scala 126:35:@22767.4]
  wire  _T_2984; // @[MemPrimitives.scala 126:35:@22768.4]
  wire  _T_2985; // @[MemPrimitives.scala 126:35:@22769.4]
  wire  _T_2986; // @[MemPrimitives.scala 126:35:@22770.4]
  wire  _T_2987; // @[MemPrimitives.scala 126:35:@22771.4]
  wire  _T_2988; // @[MemPrimitives.scala 126:35:@22772.4]
  wire  _T_2989; // @[MemPrimitives.scala 126:35:@22773.4]
  wire [10:0] _T_2991; // @[Cat.scala 30:58:@22775.4]
  wire [10:0] _T_2993; // @[Cat.scala 30:58:@22777.4]
  wire [10:0] _T_2995; // @[Cat.scala 30:58:@22779.4]
  wire [10:0] _T_2997; // @[Cat.scala 30:58:@22781.4]
  wire [10:0] _T_2999; // @[Cat.scala 30:58:@22783.4]
  wire [10:0] _T_3001; // @[Cat.scala 30:58:@22785.4]
  wire [10:0] _T_3003; // @[Cat.scala 30:58:@22787.4]
  wire [10:0] _T_3005; // @[Cat.scala 30:58:@22789.4]
  wire [10:0] _T_3007; // @[Cat.scala 30:58:@22791.4]
  wire [10:0] _T_3008; // @[Mux.scala 31:69:@22792.4]
  wire [10:0] _T_3009; // @[Mux.scala 31:69:@22793.4]
  wire [10:0] _T_3010; // @[Mux.scala 31:69:@22794.4]
  wire [10:0] _T_3011; // @[Mux.scala 31:69:@22795.4]
  wire [10:0] _T_3012; // @[Mux.scala 31:69:@22796.4]
  wire [10:0] _T_3013; // @[Mux.scala 31:69:@22797.4]
  wire [10:0] _T_3014; // @[Mux.scala 31:69:@22798.4]
  wire [10:0] _T_3015; // @[Mux.scala 31:69:@22799.4]
  wire  _T_3023; // @[MemPrimitives.scala 110:228:@22808.4]
  wire  _T_3029; // @[MemPrimitives.scala 110:228:@22812.4]
  wire  _T_3035; // @[MemPrimitives.scala 110:228:@22816.4]
  wire  _T_3041; // @[MemPrimitives.scala 110:228:@22820.4]
  wire  _T_3047; // @[MemPrimitives.scala 110:228:@22824.4]
  wire  _T_3053; // @[MemPrimitives.scala 110:228:@22828.4]
  wire  _T_3059; // @[MemPrimitives.scala 110:228:@22832.4]
  wire  _T_3065; // @[MemPrimitives.scala 110:228:@22836.4]
  wire  _T_3071; // @[MemPrimitives.scala 110:228:@22840.4]
  wire  _T_3073; // @[MemPrimitives.scala 126:35:@22854.4]
  wire  _T_3074; // @[MemPrimitives.scala 126:35:@22855.4]
  wire  _T_3075; // @[MemPrimitives.scala 126:35:@22856.4]
  wire  _T_3076; // @[MemPrimitives.scala 126:35:@22857.4]
  wire  _T_3077; // @[MemPrimitives.scala 126:35:@22858.4]
  wire  _T_3078; // @[MemPrimitives.scala 126:35:@22859.4]
  wire  _T_3079; // @[MemPrimitives.scala 126:35:@22860.4]
  wire  _T_3080; // @[MemPrimitives.scala 126:35:@22861.4]
  wire  _T_3081; // @[MemPrimitives.scala 126:35:@22862.4]
  wire [10:0] _T_3083; // @[Cat.scala 30:58:@22864.4]
  wire [10:0] _T_3085; // @[Cat.scala 30:58:@22866.4]
  wire [10:0] _T_3087; // @[Cat.scala 30:58:@22868.4]
  wire [10:0] _T_3089; // @[Cat.scala 30:58:@22870.4]
  wire [10:0] _T_3091; // @[Cat.scala 30:58:@22872.4]
  wire [10:0] _T_3093; // @[Cat.scala 30:58:@22874.4]
  wire [10:0] _T_3095; // @[Cat.scala 30:58:@22876.4]
  wire [10:0] _T_3097; // @[Cat.scala 30:58:@22878.4]
  wire [10:0] _T_3099; // @[Cat.scala 30:58:@22880.4]
  wire [10:0] _T_3100; // @[Mux.scala 31:69:@22881.4]
  wire [10:0] _T_3101; // @[Mux.scala 31:69:@22882.4]
  wire [10:0] _T_3102; // @[Mux.scala 31:69:@22883.4]
  wire [10:0] _T_3103; // @[Mux.scala 31:69:@22884.4]
  wire [10:0] _T_3104; // @[Mux.scala 31:69:@22885.4]
  wire [10:0] _T_3105; // @[Mux.scala 31:69:@22886.4]
  wire [10:0] _T_3106; // @[Mux.scala 31:69:@22887.4]
  wire [10:0] _T_3107; // @[Mux.scala 31:69:@22888.4]
  wire  _T_3115; // @[MemPrimitives.scala 110:228:@22897.4]
  wire  _T_3121; // @[MemPrimitives.scala 110:228:@22901.4]
  wire  _T_3127; // @[MemPrimitives.scala 110:228:@22905.4]
  wire  _T_3133; // @[MemPrimitives.scala 110:228:@22909.4]
  wire  _T_3139; // @[MemPrimitives.scala 110:228:@22913.4]
  wire  _T_3145; // @[MemPrimitives.scala 110:228:@22917.4]
  wire  _T_3151; // @[MemPrimitives.scala 110:228:@22921.4]
  wire  _T_3157; // @[MemPrimitives.scala 110:228:@22925.4]
  wire  _T_3163; // @[MemPrimitives.scala 110:228:@22929.4]
  wire  _T_3165; // @[MemPrimitives.scala 126:35:@22943.4]
  wire  _T_3166; // @[MemPrimitives.scala 126:35:@22944.4]
  wire  _T_3167; // @[MemPrimitives.scala 126:35:@22945.4]
  wire  _T_3168; // @[MemPrimitives.scala 126:35:@22946.4]
  wire  _T_3169; // @[MemPrimitives.scala 126:35:@22947.4]
  wire  _T_3170; // @[MemPrimitives.scala 126:35:@22948.4]
  wire  _T_3171; // @[MemPrimitives.scala 126:35:@22949.4]
  wire  _T_3172; // @[MemPrimitives.scala 126:35:@22950.4]
  wire  _T_3173; // @[MemPrimitives.scala 126:35:@22951.4]
  wire [10:0] _T_3175; // @[Cat.scala 30:58:@22953.4]
  wire [10:0] _T_3177; // @[Cat.scala 30:58:@22955.4]
  wire [10:0] _T_3179; // @[Cat.scala 30:58:@22957.4]
  wire [10:0] _T_3181; // @[Cat.scala 30:58:@22959.4]
  wire [10:0] _T_3183; // @[Cat.scala 30:58:@22961.4]
  wire [10:0] _T_3185; // @[Cat.scala 30:58:@22963.4]
  wire [10:0] _T_3187; // @[Cat.scala 30:58:@22965.4]
  wire [10:0] _T_3189; // @[Cat.scala 30:58:@22967.4]
  wire [10:0] _T_3191; // @[Cat.scala 30:58:@22969.4]
  wire [10:0] _T_3192; // @[Mux.scala 31:69:@22970.4]
  wire [10:0] _T_3193; // @[Mux.scala 31:69:@22971.4]
  wire [10:0] _T_3194; // @[Mux.scala 31:69:@22972.4]
  wire [10:0] _T_3195; // @[Mux.scala 31:69:@22973.4]
  wire [10:0] _T_3196; // @[Mux.scala 31:69:@22974.4]
  wire [10:0] _T_3197; // @[Mux.scala 31:69:@22975.4]
  wire [10:0] _T_3198; // @[Mux.scala 31:69:@22976.4]
  wire [10:0] _T_3199; // @[Mux.scala 31:69:@22977.4]
  wire  _T_3207; // @[MemPrimitives.scala 110:228:@22986.4]
  wire  _T_3213; // @[MemPrimitives.scala 110:228:@22990.4]
  wire  _T_3219; // @[MemPrimitives.scala 110:228:@22994.4]
  wire  _T_3225; // @[MemPrimitives.scala 110:228:@22998.4]
  wire  _T_3231; // @[MemPrimitives.scala 110:228:@23002.4]
  wire  _T_3237; // @[MemPrimitives.scala 110:228:@23006.4]
  wire  _T_3243; // @[MemPrimitives.scala 110:228:@23010.4]
  wire  _T_3249; // @[MemPrimitives.scala 110:228:@23014.4]
  wire  _T_3255; // @[MemPrimitives.scala 110:228:@23018.4]
  wire  _T_3257; // @[MemPrimitives.scala 126:35:@23032.4]
  wire  _T_3258; // @[MemPrimitives.scala 126:35:@23033.4]
  wire  _T_3259; // @[MemPrimitives.scala 126:35:@23034.4]
  wire  _T_3260; // @[MemPrimitives.scala 126:35:@23035.4]
  wire  _T_3261; // @[MemPrimitives.scala 126:35:@23036.4]
  wire  _T_3262; // @[MemPrimitives.scala 126:35:@23037.4]
  wire  _T_3263; // @[MemPrimitives.scala 126:35:@23038.4]
  wire  _T_3264; // @[MemPrimitives.scala 126:35:@23039.4]
  wire  _T_3265; // @[MemPrimitives.scala 126:35:@23040.4]
  wire [10:0] _T_3267; // @[Cat.scala 30:58:@23042.4]
  wire [10:0] _T_3269; // @[Cat.scala 30:58:@23044.4]
  wire [10:0] _T_3271; // @[Cat.scala 30:58:@23046.4]
  wire [10:0] _T_3273; // @[Cat.scala 30:58:@23048.4]
  wire [10:0] _T_3275; // @[Cat.scala 30:58:@23050.4]
  wire [10:0] _T_3277; // @[Cat.scala 30:58:@23052.4]
  wire [10:0] _T_3279; // @[Cat.scala 30:58:@23054.4]
  wire [10:0] _T_3281; // @[Cat.scala 30:58:@23056.4]
  wire [10:0] _T_3283; // @[Cat.scala 30:58:@23058.4]
  wire [10:0] _T_3284; // @[Mux.scala 31:69:@23059.4]
  wire [10:0] _T_3285; // @[Mux.scala 31:69:@23060.4]
  wire [10:0] _T_3286; // @[Mux.scala 31:69:@23061.4]
  wire [10:0] _T_3287; // @[Mux.scala 31:69:@23062.4]
  wire [10:0] _T_3288; // @[Mux.scala 31:69:@23063.4]
  wire [10:0] _T_3289; // @[Mux.scala 31:69:@23064.4]
  wire [10:0] _T_3290; // @[Mux.scala 31:69:@23065.4]
  wire [10:0] _T_3291; // @[Mux.scala 31:69:@23066.4]
  wire  _T_3299; // @[MemPrimitives.scala 110:228:@23075.4]
  wire  _T_3305; // @[MemPrimitives.scala 110:228:@23079.4]
  wire  _T_3311; // @[MemPrimitives.scala 110:228:@23083.4]
  wire  _T_3317; // @[MemPrimitives.scala 110:228:@23087.4]
  wire  _T_3323; // @[MemPrimitives.scala 110:228:@23091.4]
  wire  _T_3329; // @[MemPrimitives.scala 110:228:@23095.4]
  wire  _T_3335; // @[MemPrimitives.scala 110:228:@23099.4]
  wire  _T_3341; // @[MemPrimitives.scala 110:228:@23103.4]
  wire  _T_3347; // @[MemPrimitives.scala 110:228:@23107.4]
  wire  _T_3349; // @[MemPrimitives.scala 126:35:@23121.4]
  wire  _T_3350; // @[MemPrimitives.scala 126:35:@23122.4]
  wire  _T_3351; // @[MemPrimitives.scala 126:35:@23123.4]
  wire  _T_3352; // @[MemPrimitives.scala 126:35:@23124.4]
  wire  _T_3353; // @[MemPrimitives.scala 126:35:@23125.4]
  wire  _T_3354; // @[MemPrimitives.scala 126:35:@23126.4]
  wire  _T_3355; // @[MemPrimitives.scala 126:35:@23127.4]
  wire  _T_3356; // @[MemPrimitives.scala 126:35:@23128.4]
  wire  _T_3357; // @[MemPrimitives.scala 126:35:@23129.4]
  wire [10:0] _T_3359; // @[Cat.scala 30:58:@23131.4]
  wire [10:0] _T_3361; // @[Cat.scala 30:58:@23133.4]
  wire [10:0] _T_3363; // @[Cat.scala 30:58:@23135.4]
  wire [10:0] _T_3365; // @[Cat.scala 30:58:@23137.4]
  wire [10:0] _T_3367; // @[Cat.scala 30:58:@23139.4]
  wire [10:0] _T_3369; // @[Cat.scala 30:58:@23141.4]
  wire [10:0] _T_3371; // @[Cat.scala 30:58:@23143.4]
  wire [10:0] _T_3373; // @[Cat.scala 30:58:@23145.4]
  wire [10:0] _T_3375; // @[Cat.scala 30:58:@23147.4]
  wire [10:0] _T_3376; // @[Mux.scala 31:69:@23148.4]
  wire [10:0] _T_3377; // @[Mux.scala 31:69:@23149.4]
  wire [10:0] _T_3378; // @[Mux.scala 31:69:@23150.4]
  wire [10:0] _T_3379; // @[Mux.scala 31:69:@23151.4]
  wire [10:0] _T_3380; // @[Mux.scala 31:69:@23152.4]
  wire [10:0] _T_3381; // @[Mux.scala 31:69:@23153.4]
  wire [10:0] _T_3382; // @[Mux.scala 31:69:@23154.4]
  wire [10:0] _T_3383; // @[Mux.scala 31:69:@23155.4]
  wire  _T_3479; // @[package.scala 96:25:@23284.4 package.scala 96:25:@23285.4]
  wire [31:0] _T_3483; // @[Mux.scala 31:69:@23294.4]
  wire  _T_3476; // @[package.scala 96:25:@23276.4 package.scala 96:25:@23277.4]
  wire [31:0] _T_3484; // @[Mux.scala 31:69:@23295.4]
  wire  _T_3473; // @[package.scala 96:25:@23268.4 package.scala 96:25:@23269.4]
  wire [31:0] _T_3485; // @[Mux.scala 31:69:@23296.4]
  wire  _T_3470; // @[package.scala 96:25:@23260.4 package.scala 96:25:@23261.4]
  wire [31:0] _T_3486; // @[Mux.scala 31:69:@23297.4]
  wire  _T_3467; // @[package.scala 96:25:@23252.4 package.scala 96:25:@23253.4]
  wire [31:0] _T_3487; // @[Mux.scala 31:69:@23298.4]
  wire  _T_3464; // @[package.scala 96:25:@23244.4 package.scala 96:25:@23245.4]
  wire [31:0] _T_3488; // @[Mux.scala 31:69:@23299.4]
  wire  _T_3461; // @[package.scala 96:25:@23236.4 package.scala 96:25:@23237.4]
  wire [31:0] _T_3489; // @[Mux.scala 31:69:@23300.4]
  wire  _T_3458; // @[package.scala 96:25:@23228.4 package.scala 96:25:@23229.4]
  wire [31:0] _T_3490; // @[Mux.scala 31:69:@23301.4]
  wire  _T_3455; // @[package.scala 96:25:@23220.4 package.scala 96:25:@23221.4]
  wire [31:0] _T_3491; // @[Mux.scala 31:69:@23302.4]
  wire  _T_3452; // @[package.scala 96:25:@23212.4 package.scala 96:25:@23213.4]
  wire [31:0] _T_3492; // @[Mux.scala 31:69:@23303.4]
  wire  _T_3449; // @[package.scala 96:25:@23204.4 package.scala 96:25:@23205.4]
  wire  _T_3586; // @[package.scala 96:25:@23428.4 package.scala 96:25:@23429.4]
  wire [31:0] _T_3590; // @[Mux.scala 31:69:@23438.4]
  wire  _T_3583; // @[package.scala 96:25:@23420.4 package.scala 96:25:@23421.4]
  wire [31:0] _T_3591; // @[Mux.scala 31:69:@23439.4]
  wire  _T_3580; // @[package.scala 96:25:@23412.4 package.scala 96:25:@23413.4]
  wire [31:0] _T_3592; // @[Mux.scala 31:69:@23440.4]
  wire  _T_3577; // @[package.scala 96:25:@23404.4 package.scala 96:25:@23405.4]
  wire [31:0] _T_3593; // @[Mux.scala 31:69:@23441.4]
  wire  _T_3574; // @[package.scala 96:25:@23396.4 package.scala 96:25:@23397.4]
  wire [31:0] _T_3594; // @[Mux.scala 31:69:@23442.4]
  wire  _T_3571; // @[package.scala 96:25:@23388.4 package.scala 96:25:@23389.4]
  wire [31:0] _T_3595; // @[Mux.scala 31:69:@23443.4]
  wire  _T_3568; // @[package.scala 96:25:@23380.4 package.scala 96:25:@23381.4]
  wire [31:0] _T_3596; // @[Mux.scala 31:69:@23444.4]
  wire  _T_3565; // @[package.scala 96:25:@23372.4 package.scala 96:25:@23373.4]
  wire [31:0] _T_3597; // @[Mux.scala 31:69:@23445.4]
  wire  _T_3562; // @[package.scala 96:25:@23364.4 package.scala 96:25:@23365.4]
  wire [31:0] _T_3598; // @[Mux.scala 31:69:@23446.4]
  wire  _T_3559; // @[package.scala 96:25:@23356.4 package.scala 96:25:@23357.4]
  wire [31:0] _T_3599; // @[Mux.scala 31:69:@23447.4]
  wire  _T_3556; // @[package.scala 96:25:@23348.4 package.scala 96:25:@23349.4]
  wire  _T_3693; // @[package.scala 96:25:@23572.4 package.scala 96:25:@23573.4]
  wire [31:0] _T_3697; // @[Mux.scala 31:69:@23582.4]
  wire  _T_3690; // @[package.scala 96:25:@23564.4 package.scala 96:25:@23565.4]
  wire [31:0] _T_3698; // @[Mux.scala 31:69:@23583.4]
  wire  _T_3687; // @[package.scala 96:25:@23556.4 package.scala 96:25:@23557.4]
  wire [31:0] _T_3699; // @[Mux.scala 31:69:@23584.4]
  wire  _T_3684; // @[package.scala 96:25:@23548.4 package.scala 96:25:@23549.4]
  wire [31:0] _T_3700; // @[Mux.scala 31:69:@23585.4]
  wire  _T_3681; // @[package.scala 96:25:@23540.4 package.scala 96:25:@23541.4]
  wire [31:0] _T_3701; // @[Mux.scala 31:69:@23586.4]
  wire  _T_3678; // @[package.scala 96:25:@23532.4 package.scala 96:25:@23533.4]
  wire [31:0] _T_3702; // @[Mux.scala 31:69:@23587.4]
  wire  _T_3675; // @[package.scala 96:25:@23524.4 package.scala 96:25:@23525.4]
  wire [31:0] _T_3703; // @[Mux.scala 31:69:@23588.4]
  wire  _T_3672; // @[package.scala 96:25:@23516.4 package.scala 96:25:@23517.4]
  wire [31:0] _T_3704; // @[Mux.scala 31:69:@23589.4]
  wire  _T_3669; // @[package.scala 96:25:@23508.4 package.scala 96:25:@23509.4]
  wire [31:0] _T_3705; // @[Mux.scala 31:69:@23590.4]
  wire  _T_3666; // @[package.scala 96:25:@23500.4 package.scala 96:25:@23501.4]
  wire [31:0] _T_3706; // @[Mux.scala 31:69:@23591.4]
  wire  _T_3663; // @[package.scala 96:25:@23492.4 package.scala 96:25:@23493.4]
  wire  _T_3800; // @[package.scala 96:25:@23716.4 package.scala 96:25:@23717.4]
  wire [31:0] _T_3804; // @[Mux.scala 31:69:@23726.4]
  wire  _T_3797; // @[package.scala 96:25:@23708.4 package.scala 96:25:@23709.4]
  wire [31:0] _T_3805; // @[Mux.scala 31:69:@23727.4]
  wire  _T_3794; // @[package.scala 96:25:@23700.4 package.scala 96:25:@23701.4]
  wire [31:0] _T_3806; // @[Mux.scala 31:69:@23728.4]
  wire  _T_3791; // @[package.scala 96:25:@23692.4 package.scala 96:25:@23693.4]
  wire [31:0] _T_3807; // @[Mux.scala 31:69:@23729.4]
  wire  _T_3788; // @[package.scala 96:25:@23684.4 package.scala 96:25:@23685.4]
  wire [31:0] _T_3808; // @[Mux.scala 31:69:@23730.4]
  wire  _T_3785; // @[package.scala 96:25:@23676.4 package.scala 96:25:@23677.4]
  wire [31:0] _T_3809; // @[Mux.scala 31:69:@23731.4]
  wire  _T_3782; // @[package.scala 96:25:@23668.4 package.scala 96:25:@23669.4]
  wire [31:0] _T_3810; // @[Mux.scala 31:69:@23732.4]
  wire  _T_3779; // @[package.scala 96:25:@23660.4 package.scala 96:25:@23661.4]
  wire [31:0] _T_3811; // @[Mux.scala 31:69:@23733.4]
  wire  _T_3776; // @[package.scala 96:25:@23652.4 package.scala 96:25:@23653.4]
  wire [31:0] _T_3812; // @[Mux.scala 31:69:@23734.4]
  wire  _T_3773; // @[package.scala 96:25:@23644.4 package.scala 96:25:@23645.4]
  wire [31:0] _T_3813; // @[Mux.scala 31:69:@23735.4]
  wire  _T_3770; // @[package.scala 96:25:@23636.4 package.scala 96:25:@23637.4]
  wire  _T_3907; // @[package.scala 96:25:@23860.4 package.scala 96:25:@23861.4]
  wire [31:0] _T_3911; // @[Mux.scala 31:69:@23870.4]
  wire  _T_3904; // @[package.scala 96:25:@23852.4 package.scala 96:25:@23853.4]
  wire [31:0] _T_3912; // @[Mux.scala 31:69:@23871.4]
  wire  _T_3901; // @[package.scala 96:25:@23844.4 package.scala 96:25:@23845.4]
  wire [31:0] _T_3913; // @[Mux.scala 31:69:@23872.4]
  wire  _T_3898; // @[package.scala 96:25:@23836.4 package.scala 96:25:@23837.4]
  wire [31:0] _T_3914; // @[Mux.scala 31:69:@23873.4]
  wire  _T_3895; // @[package.scala 96:25:@23828.4 package.scala 96:25:@23829.4]
  wire [31:0] _T_3915; // @[Mux.scala 31:69:@23874.4]
  wire  _T_3892; // @[package.scala 96:25:@23820.4 package.scala 96:25:@23821.4]
  wire [31:0] _T_3916; // @[Mux.scala 31:69:@23875.4]
  wire  _T_3889; // @[package.scala 96:25:@23812.4 package.scala 96:25:@23813.4]
  wire [31:0] _T_3917; // @[Mux.scala 31:69:@23876.4]
  wire  _T_3886; // @[package.scala 96:25:@23804.4 package.scala 96:25:@23805.4]
  wire [31:0] _T_3918; // @[Mux.scala 31:69:@23877.4]
  wire  _T_3883; // @[package.scala 96:25:@23796.4 package.scala 96:25:@23797.4]
  wire [31:0] _T_3919; // @[Mux.scala 31:69:@23878.4]
  wire  _T_3880; // @[package.scala 96:25:@23788.4 package.scala 96:25:@23789.4]
  wire [31:0] _T_3920; // @[Mux.scala 31:69:@23879.4]
  wire  _T_3877; // @[package.scala 96:25:@23780.4 package.scala 96:25:@23781.4]
  wire  _T_4014; // @[package.scala 96:25:@24004.4 package.scala 96:25:@24005.4]
  wire [31:0] _T_4018; // @[Mux.scala 31:69:@24014.4]
  wire  _T_4011; // @[package.scala 96:25:@23996.4 package.scala 96:25:@23997.4]
  wire [31:0] _T_4019; // @[Mux.scala 31:69:@24015.4]
  wire  _T_4008; // @[package.scala 96:25:@23988.4 package.scala 96:25:@23989.4]
  wire [31:0] _T_4020; // @[Mux.scala 31:69:@24016.4]
  wire  _T_4005; // @[package.scala 96:25:@23980.4 package.scala 96:25:@23981.4]
  wire [31:0] _T_4021; // @[Mux.scala 31:69:@24017.4]
  wire  _T_4002; // @[package.scala 96:25:@23972.4 package.scala 96:25:@23973.4]
  wire [31:0] _T_4022; // @[Mux.scala 31:69:@24018.4]
  wire  _T_3999; // @[package.scala 96:25:@23964.4 package.scala 96:25:@23965.4]
  wire [31:0] _T_4023; // @[Mux.scala 31:69:@24019.4]
  wire  _T_3996; // @[package.scala 96:25:@23956.4 package.scala 96:25:@23957.4]
  wire [31:0] _T_4024; // @[Mux.scala 31:69:@24020.4]
  wire  _T_3993; // @[package.scala 96:25:@23948.4 package.scala 96:25:@23949.4]
  wire [31:0] _T_4025; // @[Mux.scala 31:69:@24021.4]
  wire  _T_3990; // @[package.scala 96:25:@23940.4 package.scala 96:25:@23941.4]
  wire [31:0] _T_4026; // @[Mux.scala 31:69:@24022.4]
  wire  _T_3987; // @[package.scala 96:25:@23932.4 package.scala 96:25:@23933.4]
  wire [31:0] _T_4027; // @[Mux.scala 31:69:@24023.4]
  wire  _T_3984; // @[package.scala 96:25:@23924.4 package.scala 96:25:@23925.4]
  wire  _T_4121; // @[package.scala 96:25:@24148.4 package.scala 96:25:@24149.4]
  wire [31:0] _T_4125; // @[Mux.scala 31:69:@24158.4]
  wire  _T_4118; // @[package.scala 96:25:@24140.4 package.scala 96:25:@24141.4]
  wire [31:0] _T_4126; // @[Mux.scala 31:69:@24159.4]
  wire  _T_4115; // @[package.scala 96:25:@24132.4 package.scala 96:25:@24133.4]
  wire [31:0] _T_4127; // @[Mux.scala 31:69:@24160.4]
  wire  _T_4112; // @[package.scala 96:25:@24124.4 package.scala 96:25:@24125.4]
  wire [31:0] _T_4128; // @[Mux.scala 31:69:@24161.4]
  wire  _T_4109; // @[package.scala 96:25:@24116.4 package.scala 96:25:@24117.4]
  wire [31:0] _T_4129; // @[Mux.scala 31:69:@24162.4]
  wire  _T_4106; // @[package.scala 96:25:@24108.4 package.scala 96:25:@24109.4]
  wire [31:0] _T_4130; // @[Mux.scala 31:69:@24163.4]
  wire  _T_4103; // @[package.scala 96:25:@24100.4 package.scala 96:25:@24101.4]
  wire [31:0] _T_4131; // @[Mux.scala 31:69:@24164.4]
  wire  _T_4100; // @[package.scala 96:25:@24092.4 package.scala 96:25:@24093.4]
  wire [31:0] _T_4132; // @[Mux.scala 31:69:@24165.4]
  wire  _T_4097; // @[package.scala 96:25:@24084.4 package.scala 96:25:@24085.4]
  wire [31:0] _T_4133; // @[Mux.scala 31:69:@24166.4]
  wire  _T_4094; // @[package.scala 96:25:@24076.4 package.scala 96:25:@24077.4]
  wire [31:0] _T_4134; // @[Mux.scala 31:69:@24167.4]
  wire  _T_4091; // @[package.scala 96:25:@24068.4 package.scala 96:25:@24069.4]
  wire  _T_4228; // @[package.scala 96:25:@24292.4 package.scala 96:25:@24293.4]
  wire [31:0] _T_4232; // @[Mux.scala 31:69:@24302.4]
  wire  _T_4225; // @[package.scala 96:25:@24284.4 package.scala 96:25:@24285.4]
  wire [31:0] _T_4233; // @[Mux.scala 31:69:@24303.4]
  wire  _T_4222; // @[package.scala 96:25:@24276.4 package.scala 96:25:@24277.4]
  wire [31:0] _T_4234; // @[Mux.scala 31:69:@24304.4]
  wire  _T_4219; // @[package.scala 96:25:@24268.4 package.scala 96:25:@24269.4]
  wire [31:0] _T_4235; // @[Mux.scala 31:69:@24305.4]
  wire  _T_4216; // @[package.scala 96:25:@24260.4 package.scala 96:25:@24261.4]
  wire [31:0] _T_4236; // @[Mux.scala 31:69:@24306.4]
  wire  _T_4213; // @[package.scala 96:25:@24252.4 package.scala 96:25:@24253.4]
  wire [31:0] _T_4237; // @[Mux.scala 31:69:@24307.4]
  wire  _T_4210; // @[package.scala 96:25:@24244.4 package.scala 96:25:@24245.4]
  wire [31:0] _T_4238; // @[Mux.scala 31:69:@24308.4]
  wire  _T_4207; // @[package.scala 96:25:@24236.4 package.scala 96:25:@24237.4]
  wire [31:0] _T_4239; // @[Mux.scala 31:69:@24309.4]
  wire  _T_4204; // @[package.scala 96:25:@24228.4 package.scala 96:25:@24229.4]
  wire [31:0] _T_4240; // @[Mux.scala 31:69:@24310.4]
  wire  _T_4201; // @[package.scala 96:25:@24220.4 package.scala 96:25:@24221.4]
  wire [31:0] _T_4241; // @[Mux.scala 31:69:@24311.4]
  wire  _T_4198; // @[package.scala 96:25:@24212.4 package.scala 96:25:@24213.4]
  wire  _T_4335; // @[package.scala 96:25:@24436.4 package.scala 96:25:@24437.4]
  wire [31:0] _T_4339; // @[Mux.scala 31:69:@24446.4]
  wire  _T_4332; // @[package.scala 96:25:@24428.4 package.scala 96:25:@24429.4]
  wire [31:0] _T_4340; // @[Mux.scala 31:69:@24447.4]
  wire  _T_4329; // @[package.scala 96:25:@24420.4 package.scala 96:25:@24421.4]
  wire [31:0] _T_4341; // @[Mux.scala 31:69:@24448.4]
  wire  _T_4326; // @[package.scala 96:25:@24412.4 package.scala 96:25:@24413.4]
  wire [31:0] _T_4342; // @[Mux.scala 31:69:@24449.4]
  wire  _T_4323; // @[package.scala 96:25:@24404.4 package.scala 96:25:@24405.4]
  wire [31:0] _T_4343; // @[Mux.scala 31:69:@24450.4]
  wire  _T_4320; // @[package.scala 96:25:@24396.4 package.scala 96:25:@24397.4]
  wire [31:0] _T_4344; // @[Mux.scala 31:69:@24451.4]
  wire  _T_4317; // @[package.scala 96:25:@24388.4 package.scala 96:25:@24389.4]
  wire [31:0] _T_4345; // @[Mux.scala 31:69:@24452.4]
  wire  _T_4314; // @[package.scala 96:25:@24380.4 package.scala 96:25:@24381.4]
  wire [31:0] _T_4346; // @[Mux.scala 31:69:@24453.4]
  wire  _T_4311; // @[package.scala 96:25:@24372.4 package.scala 96:25:@24373.4]
  wire [31:0] _T_4347; // @[Mux.scala 31:69:@24454.4]
  wire  _T_4308; // @[package.scala 96:25:@24364.4 package.scala 96:25:@24365.4]
  wire [31:0] _T_4348; // @[Mux.scala 31:69:@24455.4]
  wire  _T_4305; // @[package.scala 96:25:@24356.4 package.scala 96:25:@24357.4]
  wire  _T_4442; // @[package.scala 96:25:@24580.4 package.scala 96:25:@24581.4]
  wire [31:0] _T_4446; // @[Mux.scala 31:69:@24590.4]
  wire  _T_4439; // @[package.scala 96:25:@24572.4 package.scala 96:25:@24573.4]
  wire [31:0] _T_4447; // @[Mux.scala 31:69:@24591.4]
  wire  _T_4436; // @[package.scala 96:25:@24564.4 package.scala 96:25:@24565.4]
  wire [31:0] _T_4448; // @[Mux.scala 31:69:@24592.4]
  wire  _T_4433; // @[package.scala 96:25:@24556.4 package.scala 96:25:@24557.4]
  wire [31:0] _T_4449; // @[Mux.scala 31:69:@24593.4]
  wire  _T_4430; // @[package.scala 96:25:@24548.4 package.scala 96:25:@24549.4]
  wire [31:0] _T_4450; // @[Mux.scala 31:69:@24594.4]
  wire  _T_4427; // @[package.scala 96:25:@24540.4 package.scala 96:25:@24541.4]
  wire [31:0] _T_4451; // @[Mux.scala 31:69:@24595.4]
  wire  _T_4424; // @[package.scala 96:25:@24532.4 package.scala 96:25:@24533.4]
  wire [31:0] _T_4452; // @[Mux.scala 31:69:@24596.4]
  wire  _T_4421; // @[package.scala 96:25:@24524.4 package.scala 96:25:@24525.4]
  wire [31:0] _T_4453; // @[Mux.scala 31:69:@24597.4]
  wire  _T_4418; // @[package.scala 96:25:@24516.4 package.scala 96:25:@24517.4]
  wire [31:0] _T_4454; // @[Mux.scala 31:69:@24598.4]
  wire  _T_4415; // @[package.scala 96:25:@24508.4 package.scala 96:25:@24509.4]
  wire [31:0] _T_4455; // @[Mux.scala 31:69:@24599.4]
  wire  _T_4412; // @[package.scala 96:25:@24500.4 package.scala 96:25:@24501.4]
  wire  _T_4549; // @[package.scala 96:25:@24724.4 package.scala 96:25:@24725.4]
  wire [31:0] _T_4553; // @[Mux.scala 31:69:@24734.4]
  wire  _T_4546; // @[package.scala 96:25:@24716.4 package.scala 96:25:@24717.4]
  wire [31:0] _T_4554; // @[Mux.scala 31:69:@24735.4]
  wire  _T_4543; // @[package.scala 96:25:@24708.4 package.scala 96:25:@24709.4]
  wire [31:0] _T_4555; // @[Mux.scala 31:69:@24736.4]
  wire  _T_4540; // @[package.scala 96:25:@24700.4 package.scala 96:25:@24701.4]
  wire [31:0] _T_4556; // @[Mux.scala 31:69:@24737.4]
  wire  _T_4537; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  wire [31:0] _T_4557; // @[Mux.scala 31:69:@24738.4]
  wire  _T_4534; // @[package.scala 96:25:@24684.4 package.scala 96:25:@24685.4]
  wire [31:0] _T_4558; // @[Mux.scala 31:69:@24739.4]
  wire  _T_4531; // @[package.scala 96:25:@24676.4 package.scala 96:25:@24677.4]
  wire [31:0] _T_4559; // @[Mux.scala 31:69:@24740.4]
  wire  _T_4528; // @[package.scala 96:25:@24668.4 package.scala 96:25:@24669.4]
  wire [31:0] _T_4560; // @[Mux.scala 31:69:@24741.4]
  wire  _T_4525; // @[package.scala 96:25:@24660.4 package.scala 96:25:@24661.4]
  wire [31:0] _T_4561; // @[Mux.scala 31:69:@24742.4]
  wire  _T_4522; // @[package.scala 96:25:@24652.4 package.scala 96:25:@24653.4]
  wire [31:0] _T_4562; // @[Mux.scala 31:69:@24743.4]
  wire  _T_4519; // @[package.scala 96:25:@24644.4 package.scala 96:25:@24645.4]
  wire  _T_4656; // @[package.scala 96:25:@24868.4 package.scala 96:25:@24869.4]
  wire [31:0] _T_4660; // @[Mux.scala 31:69:@24878.4]
  wire  _T_4653; // @[package.scala 96:25:@24860.4 package.scala 96:25:@24861.4]
  wire [31:0] _T_4661; // @[Mux.scala 31:69:@24879.4]
  wire  _T_4650; // @[package.scala 96:25:@24852.4 package.scala 96:25:@24853.4]
  wire [31:0] _T_4662; // @[Mux.scala 31:69:@24880.4]
  wire  _T_4647; // @[package.scala 96:25:@24844.4 package.scala 96:25:@24845.4]
  wire [31:0] _T_4663; // @[Mux.scala 31:69:@24881.4]
  wire  _T_4644; // @[package.scala 96:25:@24836.4 package.scala 96:25:@24837.4]
  wire [31:0] _T_4664; // @[Mux.scala 31:69:@24882.4]
  wire  _T_4641; // @[package.scala 96:25:@24828.4 package.scala 96:25:@24829.4]
  wire [31:0] _T_4665; // @[Mux.scala 31:69:@24883.4]
  wire  _T_4638; // @[package.scala 96:25:@24820.4 package.scala 96:25:@24821.4]
  wire [31:0] _T_4666; // @[Mux.scala 31:69:@24884.4]
  wire  _T_4635; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  wire [31:0] _T_4667; // @[Mux.scala 31:69:@24885.4]
  wire  _T_4632; // @[package.scala 96:25:@24804.4 package.scala 96:25:@24805.4]
  wire [31:0] _T_4668; // @[Mux.scala 31:69:@24886.4]
  wire  _T_4629; // @[package.scala 96:25:@24796.4 package.scala 96:25:@24797.4]
  wire [31:0] _T_4669; // @[Mux.scala 31:69:@24887.4]
  wire  _T_4626; // @[package.scala 96:25:@24788.4 package.scala 96:25:@24789.4]
  wire  _T_4763; // @[package.scala 96:25:@25012.4 package.scala 96:25:@25013.4]
  wire [31:0] _T_4767; // @[Mux.scala 31:69:@25022.4]
  wire  _T_4760; // @[package.scala 96:25:@25004.4 package.scala 96:25:@25005.4]
  wire [31:0] _T_4768; // @[Mux.scala 31:69:@25023.4]
  wire  _T_4757; // @[package.scala 96:25:@24996.4 package.scala 96:25:@24997.4]
  wire [31:0] _T_4769; // @[Mux.scala 31:69:@25024.4]
  wire  _T_4754; // @[package.scala 96:25:@24988.4 package.scala 96:25:@24989.4]
  wire [31:0] _T_4770; // @[Mux.scala 31:69:@25025.4]
  wire  _T_4751; // @[package.scala 96:25:@24980.4 package.scala 96:25:@24981.4]
  wire [31:0] _T_4771; // @[Mux.scala 31:69:@25026.4]
  wire  _T_4748; // @[package.scala 96:25:@24972.4 package.scala 96:25:@24973.4]
  wire [31:0] _T_4772; // @[Mux.scala 31:69:@25027.4]
  wire  _T_4745; // @[package.scala 96:25:@24964.4 package.scala 96:25:@24965.4]
  wire [31:0] _T_4773; // @[Mux.scala 31:69:@25028.4]
  wire  _T_4742; // @[package.scala 96:25:@24956.4 package.scala 96:25:@24957.4]
  wire [31:0] _T_4774; // @[Mux.scala 31:69:@25029.4]
  wire  _T_4739; // @[package.scala 96:25:@24948.4 package.scala 96:25:@24949.4]
  wire [31:0] _T_4775; // @[Mux.scala 31:69:@25030.4]
  wire  _T_4736; // @[package.scala 96:25:@24940.4 package.scala 96:25:@24941.4]
  wire [31:0] _T_4776; // @[Mux.scala 31:69:@25031.4]
  wire  _T_4733; // @[package.scala 96:25:@24932.4 package.scala 96:25:@24933.4]
  wire  _T_4870; // @[package.scala 96:25:@25156.4 package.scala 96:25:@25157.4]
  wire [31:0] _T_4874; // @[Mux.scala 31:69:@25166.4]
  wire  _T_4867; // @[package.scala 96:25:@25148.4 package.scala 96:25:@25149.4]
  wire [31:0] _T_4875; // @[Mux.scala 31:69:@25167.4]
  wire  _T_4864; // @[package.scala 96:25:@25140.4 package.scala 96:25:@25141.4]
  wire [31:0] _T_4876; // @[Mux.scala 31:69:@25168.4]
  wire  _T_4861; // @[package.scala 96:25:@25132.4 package.scala 96:25:@25133.4]
  wire [31:0] _T_4877; // @[Mux.scala 31:69:@25169.4]
  wire  _T_4858; // @[package.scala 96:25:@25124.4 package.scala 96:25:@25125.4]
  wire [31:0] _T_4878; // @[Mux.scala 31:69:@25170.4]
  wire  _T_4855; // @[package.scala 96:25:@25116.4 package.scala 96:25:@25117.4]
  wire [31:0] _T_4879; // @[Mux.scala 31:69:@25171.4]
  wire  _T_4852; // @[package.scala 96:25:@25108.4 package.scala 96:25:@25109.4]
  wire [31:0] _T_4880; // @[Mux.scala 31:69:@25172.4]
  wire  _T_4849; // @[package.scala 96:25:@25100.4 package.scala 96:25:@25101.4]
  wire [31:0] _T_4881; // @[Mux.scala 31:69:@25173.4]
  wire  _T_4846; // @[package.scala 96:25:@25092.4 package.scala 96:25:@25093.4]
  wire [31:0] _T_4882; // @[Mux.scala 31:69:@25174.4]
  wire  _T_4843; // @[package.scala 96:25:@25084.4 package.scala 96:25:@25085.4]
  wire [31:0] _T_4883; // @[Mux.scala 31:69:@25175.4]
  wire  _T_4840; // @[package.scala 96:25:@25076.4 package.scala 96:25:@25077.4]
  wire  _T_4977; // @[package.scala 96:25:@25300.4 package.scala 96:25:@25301.4]
  wire [31:0] _T_4981; // @[Mux.scala 31:69:@25310.4]
  wire  _T_4974; // @[package.scala 96:25:@25292.4 package.scala 96:25:@25293.4]
  wire [31:0] _T_4982; // @[Mux.scala 31:69:@25311.4]
  wire  _T_4971; // @[package.scala 96:25:@25284.4 package.scala 96:25:@25285.4]
  wire [31:0] _T_4983; // @[Mux.scala 31:69:@25312.4]
  wire  _T_4968; // @[package.scala 96:25:@25276.4 package.scala 96:25:@25277.4]
  wire [31:0] _T_4984; // @[Mux.scala 31:69:@25313.4]
  wire  _T_4965; // @[package.scala 96:25:@25268.4 package.scala 96:25:@25269.4]
  wire [31:0] _T_4985; // @[Mux.scala 31:69:@25314.4]
  wire  _T_4962; // @[package.scala 96:25:@25260.4 package.scala 96:25:@25261.4]
  wire [31:0] _T_4986; // @[Mux.scala 31:69:@25315.4]
  wire  _T_4959; // @[package.scala 96:25:@25252.4 package.scala 96:25:@25253.4]
  wire [31:0] _T_4987; // @[Mux.scala 31:69:@25316.4]
  wire  _T_4956; // @[package.scala 96:25:@25244.4 package.scala 96:25:@25245.4]
  wire [31:0] _T_4988; // @[Mux.scala 31:69:@25317.4]
  wire  _T_4953; // @[package.scala 96:25:@25236.4 package.scala 96:25:@25237.4]
  wire [31:0] _T_4989; // @[Mux.scala 31:69:@25318.4]
  wire  _T_4950; // @[package.scala 96:25:@25228.4 package.scala 96:25:@25229.4]
  wire [31:0] _T_4990; // @[Mux.scala 31:69:@25319.4]
  wire  _T_4947; // @[package.scala 96:25:@25220.4 package.scala 96:25:@25221.4]
  wire  _T_5084; // @[package.scala 96:25:@25444.4 package.scala 96:25:@25445.4]
  wire [31:0] _T_5088; // @[Mux.scala 31:69:@25454.4]
  wire  _T_5081; // @[package.scala 96:25:@25436.4 package.scala 96:25:@25437.4]
  wire [31:0] _T_5089; // @[Mux.scala 31:69:@25455.4]
  wire  _T_5078; // @[package.scala 96:25:@25428.4 package.scala 96:25:@25429.4]
  wire [31:0] _T_5090; // @[Mux.scala 31:69:@25456.4]
  wire  _T_5075; // @[package.scala 96:25:@25420.4 package.scala 96:25:@25421.4]
  wire [31:0] _T_5091; // @[Mux.scala 31:69:@25457.4]
  wire  _T_5072; // @[package.scala 96:25:@25412.4 package.scala 96:25:@25413.4]
  wire [31:0] _T_5092; // @[Mux.scala 31:69:@25458.4]
  wire  _T_5069; // @[package.scala 96:25:@25404.4 package.scala 96:25:@25405.4]
  wire [31:0] _T_5093; // @[Mux.scala 31:69:@25459.4]
  wire  _T_5066; // @[package.scala 96:25:@25396.4 package.scala 96:25:@25397.4]
  wire [31:0] _T_5094; // @[Mux.scala 31:69:@25460.4]
  wire  _T_5063; // @[package.scala 96:25:@25388.4 package.scala 96:25:@25389.4]
  wire [31:0] _T_5095; // @[Mux.scala 31:69:@25461.4]
  wire  _T_5060; // @[package.scala 96:25:@25380.4 package.scala 96:25:@25381.4]
  wire [31:0] _T_5096; // @[Mux.scala 31:69:@25462.4]
  wire  _T_5057; // @[package.scala 96:25:@25372.4 package.scala 96:25:@25373.4]
  wire [31:0] _T_5097; // @[Mux.scala 31:69:@25463.4]
  wire  _T_5054; // @[package.scala 96:25:@25364.4 package.scala 96:25:@25365.4]
  wire  _T_5191; // @[package.scala 96:25:@25588.4 package.scala 96:25:@25589.4]
  wire [31:0] _T_5195; // @[Mux.scala 31:69:@25598.4]
  wire  _T_5188; // @[package.scala 96:25:@25580.4 package.scala 96:25:@25581.4]
  wire [31:0] _T_5196; // @[Mux.scala 31:69:@25599.4]
  wire  _T_5185; // @[package.scala 96:25:@25572.4 package.scala 96:25:@25573.4]
  wire [31:0] _T_5197; // @[Mux.scala 31:69:@25600.4]
  wire  _T_5182; // @[package.scala 96:25:@25564.4 package.scala 96:25:@25565.4]
  wire [31:0] _T_5198; // @[Mux.scala 31:69:@25601.4]
  wire  _T_5179; // @[package.scala 96:25:@25556.4 package.scala 96:25:@25557.4]
  wire [31:0] _T_5199; // @[Mux.scala 31:69:@25602.4]
  wire  _T_5176; // @[package.scala 96:25:@25548.4 package.scala 96:25:@25549.4]
  wire [31:0] _T_5200; // @[Mux.scala 31:69:@25603.4]
  wire  _T_5173; // @[package.scala 96:25:@25540.4 package.scala 96:25:@25541.4]
  wire [31:0] _T_5201; // @[Mux.scala 31:69:@25604.4]
  wire  _T_5170; // @[package.scala 96:25:@25532.4 package.scala 96:25:@25533.4]
  wire [31:0] _T_5202; // @[Mux.scala 31:69:@25605.4]
  wire  _T_5167; // @[package.scala 96:25:@25524.4 package.scala 96:25:@25525.4]
  wire [31:0] _T_5203; // @[Mux.scala 31:69:@25606.4]
  wire  _T_5164; // @[package.scala 96:25:@25516.4 package.scala 96:25:@25517.4]
  wire [31:0] _T_5204; // @[Mux.scala 31:69:@25607.4]
  wire  _T_5161; // @[package.scala 96:25:@25508.4 package.scala 96:25:@25509.4]
  wire  _T_5298; // @[package.scala 96:25:@25732.4 package.scala 96:25:@25733.4]
  wire [31:0] _T_5302; // @[Mux.scala 31:69:@25742.4]
  wire  _T_5295; // @[package.scala 96:25:@25724.4 package.scala 96:25:@25725.4]
  wire [31:0] _T_5303; // @[Mux.scala 31:69:@25743.4]
  wire  _T_5292; // @[package.scala 96:25:@25716.4 package.scala 96:25:@25717.4]
  wire [31:0] _T_5304; // @[Mux.scala 31:69:@25744.4]
  wire  _T_5289; // @[package.scala 96:25:@25708.4 package.scala 96:25:@25709.4]
  wire [31:0] _T_5305; // @[Mux.scala 31:69:@25745.4]
  wire  _T_5286; // @[package.scala 96:25:@25700.4 package.scala 96:25:@25701.4]
  wire [31:0] _T_5306; // @[Mux.scala 31:69:@25746.4]
  wire  _T_5283; // @[package.scala 96:25:@25692.4 package.scala 96:25:@25693.4]
  wire [31:0] _T_5307; // @[Mux.scala 31:69:@25747.4]
  wire  _T_5280; // @[package.scala 96:25:@25684.4 package.scala 96:25:@25685.4]
  wire [31:0] _T_5308; // @[Mux.scala 31:69:@25748.4]
  wire  _T_5277; // @[package.scala 96:25:@25676.4 package.scala 96:25:@25677.4]
  wire [31:0] _T_5309; // @[Mux.scala 31:69:@25749.4]
  wire  _T_5274; // @[package.scala 96:25:@25668.4 package.scala 96:25:@25669.4]
  wire [31:0] _T_5310; // @[Mux.scala 31:69:@25750.4]
  wire  _T_5271; // @[package.scala 96:25:@25660.4 package.scala 96:25:@25661.4]
  wire [31:0] _T_5311; // @[Mux.scala 31:69:@25751.4]
  wire  _T_5268; // @[package.scala 96:25:@25652.4 package.scala 96:25:@25653.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@20186.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@20202.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@20218.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@20234.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@20250.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@20266.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@20282.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@20298.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@20314.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@20330.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@20346.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@20362.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@20378.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@20394.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@20410.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@20426.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  Mem1D_5 Mem1D_16 ( // @[MemPrimitives.scala 64:21:@20442.4]
    .clock(Mem1D_16_clock),
    .reset(Mem1D_16_reset),
    .io_r_ofs_0(Mem1D_16_io_r_ofs_0),
    .io_r_backpressure(Mem1D_16_io_r_backpressure),
    .io_w_ofs_0(Mem1D_16_io_w_ofs_0),
    .io_w_data_0(Mem1D_16_io_w_data_0),
    .io_w_en_0(Mem1D_16_io_w_en_0),
    .io_output(Mem1D_16_io_output)
  );
  Mem1D_5 Mem1D_17 ( // @[MemPrimitives.scala 64:21:@20458.4]
    .clock(Mem1D_17_clock),
    .reset(Mem1D_17_reset),
    .io_r_ofs_0(Mem1D_17_io_r_ofs_0),
    .io_r_backpressure(Mem1D_17_io_r_backpressure),
    .io_w_ofs_0(Mem1D_17_io_w_ofs_0),
    .io_w_data_0(Mem1D_17_io_w_data_0),
    .io_w_en_0(Mem1D_17_io_w_en_0),
    .io_output(Mem1D_17_io_output)
  );
  Mem1D_5 Mem1D_18 ( // @[MemPrimitives.scala 64:21:@20474.4]
    .clock(Mem1D_18_clock),
    .reset(Mem1D_18_reset),
    .io_r_ofs_0(Mem1D_18_io_r_ofs_0),
    .io_r_backpressure(Mem1D_18_io_r_backpressure),
    .io_w_ofs_0(Mem1D_18_io_w_ofs_0),
    .io_w_data_0(Mem1D_18_io_w_data_0),
    .io_w_en_0(Mem1D_18_io_w_en_0),
    .io_output(Mem1D_18_io_output)
  );
  Mem1D_5 Mem1D_19 ( // @[MemPrimitives.scala 64:21:@20490.4]
    .clock(Mem1D_19_clock),
    .reset(Mem1D_19_reset),
    .io_r_ofs_0(Mem1D_19_io_r_ofs_0),
    .io_r_backpressure(Mem1D_19_io_r_backpressure),
    .io_w_ofs_0(Mem1D_19_io_w_ofs_0),
    .io_w_data_0(Mem1D_19_io_w_data_0),
    .io_w_en_0(Mem1D_19_io_w_en_0),
    .io_output(Mem1D_19_io_output)
  );
  Mem1D_5 Mem1D_20 ( // @[MemPrimitives.scala 64:21:@20506.4]
    .clock(Mem1D_20_clock),
    .reset(Mem1D_20_reset),
    .io_r_ofs_0(Mem1D_20_io_r_ofs_0),
    .io_r_backpressure(Mem1D_20_io_r_backpressure),
    .io_w_ofs_0(Mem1D_20_io_w_ofs_0),
    .io_w_data_0(Mem1D_20_io_w_data_0),
    .io_w_en_0(Mem1D_20_io_w_en_0),
    .io_output(Mem1D_20_io_output)
  );
  Mem1D_5 Mem1D_21 ( // @[MemPrimitives.scala 64:21:@20522.4]
    .clock(Mem1D_21_clock),
    .reset(Mem1D_21_reset),
    .io_r_ofs_0(Mem1D_21_io_r_ofs_0),
    .io_r_backpressure(Mem1D_21_io_r_backpressure),
    .io_w_ofs_0(Mem1D_21_io_w_ofs_0),
    .io_w_data_0(Mem1D_21_io_w_data_0),
    .io_w_en_0(Mem1D_21_io_w_en_0),
    .io_output(Mem1D_21_io_output)
  );
  Mem1D_5 Mem1D_22 ( // @[MemPrimitives.scala 64:21:@20538.4]
    .clock(Mem1D_22_clock),
    .reset(Mem1D_22_reset),
    .io_r_ofs_0(Mem1D_22_io_r_ofs_0),
    .io_r_backpressure(Mem1D_22_io_r_backpressure),
    .io_w_ofs_0(Mem1D_22_io_w_ofs_0),
    .io_w_data_0(Mem1D_22_io_w_data_0),
    .io_w_en_0(Mem1D_22_io_w_en_0),
    .io_output(Mem1D_22_io_output)
  );
  Mem1D_5 Mem1D_23 ( // @[MemPrimitives.scala 64:21:@20554.4]
    .clock(Mem1D_23_clock),
    .reset(Mem1D_23_reset),
    .io_r_ofs_0(Mem1D_23_io_r_ofs_0),
    .io_r_backpressure(Mem1D_23_io_r_backpressure),
    .io_w_ofs_0(Mem1D_23_io_w_ofs_0),
    .io_w_data_0(Mem1D_23_io_w_data_0),
    .io_w_en_0(Mem1D_23_io_w_en_0),
    .io_output(Mem1D_23_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@21062.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@21151.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@21240.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@21329.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@21418.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@21507.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@21596.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@21685.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@21774.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@21863.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@21952.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@22041.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@22130.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_ins_6(StickySelects_12_io_ins_6),
    .io_ins_7(StickySelects_12_io_ins_7),
    .io_ins_8(StickySelects_12_io_ins_8),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5),
    .io_outs_6(StickySelects_12_io_outs_6),
    .io_outs_7(StickySelects_12_io_outs_7),
    .io_outs_8(StickySelects_12_io_outs_8)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@22219.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_ins_6(StickySelects_13_io_ins_6),
    .io_ins_7(StickySelects_13_io_ins_7),
    .io_ins_8(StickySelects_13_io_ins_8),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5),
    .io_outs_6(StickySelects_13_io_outs_6),
    .io_outs_7(StickySelects_13_io_outs_7),
    .io_outs_8(StickySelects_13_io_outs_8)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@22308.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_ins_8(StickySelects_14_io_ins_8),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7),
    .io_outs_8(StickySelects_14_io_outs_8)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@22397.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_ins_8(StickySelects_15_io_ins_8),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7),
    .io_outs_8(StickySelects_15_io_outs_8)
  );
  StickySelects_1 StickySelects_16 ( // @[MemPrimitives.scala 124:33:@22486.4]
    .clock(StickySelects_16_clock),
    .reset(StickySelects_16_reset),
    .io_ins_0(StickySelects_16_io_ins_0),
    .io_ins_1(StickySelects_16_io_ins_1),
    .io_ins_2(StickySelects_16_io_ins_2),
    .io_ins_3(StickySelects_16_io_ins_3),
    .io_ins_4(StickySelects_16_io_ins_4),
    .io_ins_5(StickySelects_16_io_ins_5),
    .io_ins_6(StickySelects_16_io_ins_6),
    .io_ins_7(StickySelects_16_io_ins_7),
    .io_ins_8(StickySelects_16_io_ins_8),
    .io_outs_0(StickySelects_16_io_outs_0),
    .io_outs_1(StickySelects_16_io_outs_1),
    .io_outs_2(StickySelects_16_io_outs_2),
    .io_outs_3(StickySelects_16_io_outs_3),
    .io_outs_4(StickySelects_16_io_outs_4),
    .io_outs_5(StickySelects_16_io_outs_5),
    .io_outs_6(StickySelects_16_io_outs_6),
    .io_outs_7(StickySelects_16_io_outs_7),
    .io_outs_8(StickySelects_16_io_outs_8)
  );
  StickySelects_1 StickySelects_17 ( // @[MemPrimitives.scala 124:33:@22575.4]
    .clock(StickySelects_17_clock),
    .reset(StickySelects_17_reset),
    .io_ins_0(StickySelects_17_io_ins_0),
    .io_ins_1(StickySelects_17_io_ins_1),
    .io_ins_2(StickySelects_17_io_ins_2),
    .io_ins_3(StickySelects_17_io_ins_3),
    .io_ins_4(StickySelects_17_io_ins_4),
    .io_ins_5(StickySelects_17_io_ins_5),
    .io_ins_6(StickySelects_17_io_ins_6),
    .io_ins_7(StickySelects_17_io_ins_7),
    .io_ins_8(StickySelects_17_io_ins_8),
    .io_outs_0(StickySelects_17_io_outs_0),
    .io_outs_1(StickySelects_17_io_outs_1),
    .io_outs_2(StickySelects_17_io_outs_2),
    .io_outs_3(StickySelects_17_io_outs_3),
    .io_outs_4(StickySelects_17_io_outs_4),
    .io_outs_5(StickySelects_17_io_outs_5),
    .io_outs_6(StickySelects_17_io_outs_6),
    .io_outs_7(StickySelects_17_io_outs_7),
    .io_outs_8(StickySelects_17_io_outs_8)
  );
  StickySelects_1 StickySelects_18 ( // @[MemPrimitives.scala 124:33:@22664.4]
    .clock(StickySelects_18_clock),
    .reset(StickySelects_18_reset),
    .io_ins_0(StickySelects_18_io_ins_0),
    .io_ins_1(StickySelects_18_io_ins_1),
    .io_ins_2(StickySelects_18_io_ins_2),
    .io_ins_3(StickySelects_18_io_ins_3),
    .io_ins_4(StickySelects_18_io_ins_4),
    .io_ins_5(StickySelects_18_io_ins_5),
    .io_ins_6(StickySelects_18_io_ins_6),
    .io_ins_7(StickySelects_18_io_ins_7),
    .io_ins_8(StickySelects_18_io_ins_8),
    .io_outs_0(StickySelects_18_io_outs_0),
    .io_outs_1(StickySelects_18_io_outs_1),
    .io_outs_2(StickySelects_18_io_outs_2),
    .io_outs_3(StickySelects_18_io_outs_3),
    .io_outs_4(StickySelects_18_io_outs_4),
    .io_outs_5(StickySelects_18_io_outs_5),
    .io_outs_6(StickySelects_18_io_outs_6),
    .io_outs_7(StickySelects_18_io_outs_7),
    .io_outs_8(StickySelects_18_io_outs_8)
  );
  StickySelects_1 StickySelects_19 ( // @[MemPrimitives.scala 124:33:@22753.4]
    .clock(StickySelects_19_clock),
    .reset(StickySelects_19_reset),
    .io_ins_0(StickySelects_19_io_ins_0),
    .io_ins_1(StickySelects_19_io_ins_1),
    .io_ins_2(StickySelects_19_io_ins_2),
    .io_ins_3(StickySelects_19_io_ins_3),
    .io_ins_4(StickySelects_19_io_ins_4),
    .io_ins_5(StickySelects_19_io_ins_5),
    .io_ins_6(StickySelects_19_io_ins_6),
    .io_ins_7(StickySelects_19_io_ins_7),
    .io_ins_8(StickySelects_19_io_ins_8),
    .io_outs_0(StickySelects_19_io_outs_0),
    .io_outs_1(StickySelects_19_io_outs_1),
    .io_outs_2(StickySelects_19_io_outs_2),
    .io_outs_3(StickySelects_19_io_outs_3),
    .io_outs_4(StickySelects_19_io_outs_4),
    .io_outs_5(StickySelects_19_io_outs_5),
    .io_outs_6(StickySelects_19_io_outs_6),
    .io_outs_7(StickySelects_19_io_outs_7),
    .io_outs_8(StickySelects_19_io_outs_8)
  );
  StickySelects_1 StickySelects_20 ( // @[MemPrimitives.scala 124:33:@22842.4]
    .clock(StickySelects_20_clock),
    .reset(StickySelects_20_reset),
    .io_ins_0(StickySelects_20_io_ins_0),
    .io_ins_1(StickySelects_20_io_ins_1),
    .io_ins_2(StickySelects_20_io_ins_2),
    .io_ins_3(StickySelects_20_io_ins_3),
    .io_ins_4(StickySelects_20_io_ins_4),
    .io_ins_5(StickySelects_20_io_ins_5),
    .io_ins_6(StickySelects_20_io_ins_6),
    .io_ins_7(StickySelects_20_io_ins_7),
    .io_ins_8(StickySelects_20_io_ins_8),
    .io_outs_0(StickySelects_20_io_outs_0),
    .io_outs_1(StickySelects_20_io_outs_1),
    .io_outs_2(StickySelects_20_io_outs_2),
    .io_outs_3(StickySelects_20_io_outs_3),
    .io_outs_4(StickySelects_20_io_outs_4),
    .io_outs_5(StickySelects_20_io_outs_5),
    .io_outs_6(StickySelects_20_io_outs_6),
    .io_outs_7(StickySelects_20_io_outs_7),
    .io_outs_8(StickySelects_20_io_outs_8)
  );
  StickySelects_1 StickySelects_21 ( // @[MemPrimitives.scala 124:33:@22931.4]
    .clock(StickySelects_21_clock),
    .reset(StickySelects_21_reset),
    .io_ins_0(StickySelects_21_io_ins_0),
    .io_ins_1(StickySelects_21_io_ins_1),
    .io_ins_2(StickySelects_21_io_ins_2),
    .io_ins_3(StickySelects_21_io_ins_3),
    .io_ins_4(StickySelects_21_io_ins_4),
    .io_ins_5(StickySelects_21_io_ins_5),
    .io_ins_6(StickySelects_21_io_ins_6),
    .io_ins_7(StickySelects_21_io_ins_7),
    .io_ins_8(StickySelects_21_io_ins_8),
    .io_outs_0(StickySelects_21_io_outs_0),
    .io_outs_1(StickySelects_21_io_outs_1),
    .io_outs_2(StickySelects_21_io_outs_2),
    .io_outs_3(StickySelects_21_io_outs_3),
    .io_outs_4(StickySelects_21_io_outs_4),
    .io_outs_5(StickySelects_21_io_outs_5),
    .io_outs_6(StickySelects_21_io_outs_6),
    .io_outs_7(StickySelects_21_io_outs_7),
    .io_outs_8(StickySelects_21_io_outs_8)
  );
  StickySelects_1 StickySelects_22 ( // @[MemPrimitives.scala 124:33:@23020.4]
    .clock(StickySelects_22_clock),
    .reset(StickySelects_22_reset),
    .io_ins_0(StickySelects_22_io_ins_0),
    .io_ins_1(StickySelects_22_io_ins_1),
    .io_ins_2(StickySelects_22_io_ins_2),
    .io_ins_3(StickySelects_22_io_ins_3),
    .io_ins_4(StickySelects_22_io_ins_4),
    .io_ins_5(StickySelects_22_io_ins_5),
    .io_ins_6(StickySelects_22_io_ins_6),
    .io_ins_7(StickySelects_22_io_ins_7),
    .io_ins_8(StickySelects_22_io_ins_8),
    .io_outs_0(StickySelects_22_io_outs_0),
    .io_outs_1(StickySelects_22_io_outs_1),
    .io_outs_2(StickySelects_22_io_outs_2),
    .io_outs_3(StickySelects_22_io_outs_3),
    .io_outs_4(StickySelects_22_io_outs_4),
    .io_outs_5(StickySelects_22_io_outs_5),
    .io_outs_6(StickySelects_22_io_outs_6),
    .io_outs_7(StickySelects_22_io_outs_7),
    .io_outs_8(StickySelects_22_io_outs_8)
  );
  StickySelects_1 StickySelects_23 ( // @[MemPrimitives.scala 124:33:@23109.4]
    .clock(StickySelects_23_clock),
    .reset(StickySelects_23_reset),
    .io_ins_0(StickySelects_23_io_ins_0),
    .io_ins_1(StickySelects_23_io_ins_1),
    .io_ins_2(StickySelects_23_io_ins_2),
    .io_ins_3(StickySelects_23_io_ins_3),
    .io_ins_4(StickySelects_23_io_ins_4),
    .io_ins_5(StickySelects_23_io_ins_5),
    .io_ins_6(StickySelects_23_io_ins_6),
    .io_ins_7(StickySelects_23_io_ins_7),
    .io_ins_8(StickySelects_23_io_ins_8),
    .io_outs_0(StickySelects_23_io_outs_0),
    .io_outs_1(StickySelects_23_io_outs_1),
    .io_outs_2(StickySelects_23_io_outs_2),
    .io_outs_3(StickySelects_23_io_outs_3),
    .io_outs_4(StickySelects_23_io_outs_4),
    .io_outs_5(StickySelects_23_io_outs_5),
    .io_outs_6(StickySelects_23_io_outs_6),
    .io_outs_7(StickySelects_23_io_outs_7),
    .io_outs_8(StickySelects_23_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@23199.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@23207.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@23215.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@23223.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@23231.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@23239.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@23247.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@23255.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@23263.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@23271.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@23279.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@23287.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@23343.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@23351.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@23359.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@23367.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@23375.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@23383.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@23391.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@23399.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@23407.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@23415.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@23423.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@23431.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@23487.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@23495.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@23503.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@23511.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@23519.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@23527.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@23535.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@23543.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@23551.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@23559.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@23567.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@23575.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@23631.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@23639.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@23647.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@23655.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@23663.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@23671.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@23679.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@23687.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@23695.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@23703.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@23711.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@23719.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@23775.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@23783.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@23791.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@23799.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@23807.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@23815.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@23823.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@23831.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@23839.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@23847.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@23855.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@23863.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@23919.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@23927.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@23935.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@23943.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@23951.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@23959.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@23967.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@23975.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@23983.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@23991.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@23999.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@24007.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@24063.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@24071.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@24079.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@24087.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@24095.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@24103.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@24111.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@24119.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@24127.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@24135.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@24143.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@24151.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@24207.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@24215.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@24223.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@24231.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@24239.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@24247.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@24255.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@24263.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@24271.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@24279.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@24287.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@24295.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@24351.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@24359.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@24367.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@24375.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@24383.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@24391.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@24399.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@24407.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@24415.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@24423.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@24431.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@24439.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_108 ( // @[package.scala 93:22:@24495.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_109 ( // @[package.scala 93:22:@24503.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_110 ( // @[package.scala 93:22:@24511.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_111 ( // @[package.scala 93:22:@24519.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_112 ( // @[package.scala 93:22:@24527.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_113 ( // @[package.scala 93:22:@24535.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_114 ( // @[package.scala 93:22:@24543.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_115 ( // @[package.scala 93:22:@24551.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_116 ( // @[package.scala 93:22:@24559.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_117 ( // @[package.scala 93:22:@24567.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_118 ( // @[package.scala 93:22:@24575.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_119 ( // @[package.scala 93:22:@24583.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_120 ( // @[package.scala 93:22:@24639.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_121 ( // @[package.scala 93:22:@24647.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_122 ( // @[package.scala 93:22:@24655.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_123 ( // @[package.scala 93:22:@24663.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_124 ( // @[package.scala 93:22:@24671.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_125 ( // @[package.scala 93:22:@24679.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_126 ( // @[package.scala 93:22:@24687.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_127 ( // @[package.scala 93:22:@24695.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_128 ( // @[package.scala 93:22:@24703.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_129 ( // @[package.scala 93:22:@24711.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_130 ( // @[package.scala 93:22:@24719.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_131 ( // @[package.scala 93:22:@24727.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_132 ( // @[package.scala 93:22:@24783.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_133 ( // @[package.scala 93:22:@24791.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_134 ( // @[package.scala 93:22:@24799.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_135 ( // @[package.scala 93:22:@24807.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_136 ( // @[package.scala 93:22:@24815.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_137 ( // @[package.scala 93:22:@24823.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_138 ( // @[package.scala 93:22:@24831.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_139 ( // @[package.scala 93:22:@24839.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_140 ( // @[package.scala 93:22:@24847.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_141 ( // @[package.scala 93:22:@24855.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_142 ( // @[package.scala 93:22:@24863.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_143 ( // @[package.scala 93:22:@24871.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_144 ( // @[package.scala 93:22:@24927.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_145 ( // @[package.scala 93:22:@24935.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_146 ( // @[package.scala 93:22:@24943.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_147 ( // @[package.scala 93:22:@24951.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_148 ( // @[package.scala 93:22:@24959.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_149 ( // @[package.scala 93:22:@24967.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_150 ( // @[package.scala 93:22:@24975.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_151 ( // @[package.scala 93:22:@24983.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_152 ( // @[package.scala 93:22:@24991.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_153 ( // @[package.scala 93:22:@24999.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_154 ( // @[package.scala 93:22:@25007.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_155 ( // @[package.scala 93:22:@25015.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_156 ( // @[package.scala 93:22:@25071.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_157 ( // @[package.scala 93:22:@25079.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_158 ( // @[package.scala 93:22:@25087.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_159 ( // @[package.scala 93:22:@25095.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_160 ( // @[package.scala 93:22:@25103.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_161 ( // @[package.scala 93:22:@25111.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_162 ( // @[package.scala 93:22:@25119.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_163 ( // @[package.scala 93:22:@25127.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_164 ( // @[package.scala 93:22:@25135.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_165 ( // @[package.scala 93:22:@25143.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_166 ( // @[package.scala 93:22:@25151.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_167 ( // @[package.scala 93:22:@25159.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_168 ( // @[package.scala 93:22:@25215.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_169 ( // @[package.scala 93:22:@25223.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_170 ( // @[package.scala 93:22:@25231.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_171 ( // @[package.scala 93:22:@25239.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_172 ( // @[package.scala 93:22:@25247.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_173 ( // @[package.scala 93:22:@25255.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_174 ( // @[package.scala 93:22:@25263.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_175 ( // @[package.scala 93:22:@25271.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_176 ( // @[package.scala 93:22:@25279.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_177 ( // @[package.scala 93:22:@25287.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_178 ( // @[package.scala 93:22:@25295.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_179 ( // @[package.scala 93:22:@25303.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_180 ( // @[package.scala 93:22:@25359.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_181 ( // @[package.scala 93:22:@25367.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_182 ( // @[package.scala 93:22:@25375.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_183 ( // @[package.scala 93:22:@25383.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_184 ( // @[package.scala 93:22:@25391.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_185 ( // @[package.scala 93:22:@25399.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_186 ( // @[package.scala 93:22:@25407.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_187 ( // @[package.scala 93:22:@25415.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_188 ( // @[package.scala 93:22:@25423.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_189 ( // @[package.scala 93:22:@25431.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_190 ( // @[package.scala 93:22:@25439.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_191 ( // @[package.scala 93:22:@25447.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_192 ( // @[package.scala 93:22:@25503.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_193 ( // @[package.scala 93:22:@25511.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_194 ( // @[package.scala 93:22:@25519.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_195 ( // @[package.scala 93:22:@25527.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_196 ( // @[package.scala 93:22:@25535.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_197 ( // @[package.scala 93:22:@25543.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_198 ( // @[package.scala 93:22:@25551.4]
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_199 ( // @[package.scala 93:22:@25559.4]
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_200 ( // @[package.scala 93:22:@25567.4]
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_201 ( // @[package.scala 93:22:@25575.4]
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_202 ( // @[package.scala 93:22:@25583.4]
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_203 ( // @[package.scala 93:22:@25591.4]
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_204 ( // @[package.scala 93:22:@25647.4]
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_205 ( // @[package.scala 93:22:@25655.4]
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_206 ( // @[package.scala 93:22:@25663.4]
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_207 ( // @[package.scala 93:22:@25671.4]
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_208 ( // @[package.scala 93:22:@25679.4]
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_209 ( // @[package.scala 93:22:@25687.4]
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_210 ( // @[package.scala 93:22:@25695.4]
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_211 ( // @[package.scala 93:22:@25703.4]
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_212 ( // @[package.scala 93:22:@25711.4]
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_213 ( // @[package.scala 93:22:@25719.4]
    .clock(RetimeWrapper_213_clock),
    .reset(RetimeWrapper_213_reset),
    .io_flow(RetimeWrapper_213_io_flow),
    .io_in(RetimeWrapper_213_io_in),
    .io_out(RetimeWrapper_213_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_214 ( // @[package.scala 93:22:@25727.4]
    .clock(RetimeWrapper_214_clock),
    .reset(RetimeWrapper_214_reset),
    .io_flow(RetimeWrapper_214_io_flow),
    .io_in(RetimeWrapper_214_io_in),
    .io_out(RetimeWrapper_214_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_215 ( // @[package.scala 93:22:@25735.4]
    .clock(RetimeWrapper_215_clock),
    .reset(RetimeWrapper_215_reset),
    .io_flow(RetimeWrapper_215_io_flow),
    .io_in(RetimeWrapper_215_io_in),
    .io_out(RetimeWrapper_215_io_out)
  );
  assign _T_700 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20570.4]
  assign _T_702 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@20571.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 82:228:@20572.4]
  assign _T_704 = io_wPort_0_en_0 & _T_703; // @[MemPrimitives.scala 83:102:@20573.4]
  assign _T_706 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20574.4]
  assign _T_708 = io_wPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@20575.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 82:228:@20576.4]
  assign _T_710 = io_wPort_2_en_0 & _T_709; // @[MemPrimitives.scala 83:102:@20577.4]
  assign _T_712 = {_T_704,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20579.4]
  assign _T_714 = {_T_710,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20581.4]
  assign _T_715 = _T_704 ? _T_712 : _T_714; // @[Mux.scala 31:69:@20582.4]
  assign _T_720 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20589.4]
  assign _T_722 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@20590.4]
  assign _T_723 = _T_720 & _T_722; // @[MemPrimitives.scala 82:228:@20591.4]
  assign _T_724 = io_wPort_1_en_0 & _T_723; // @[MemPrimitives.scala 83:102:@20592.4]
  assign _T_726 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20593.4]
  assign _T_728 = io_wPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@20594.4]
  assign _T_729 = _T_726 & _T_728; // @[MemPrimitives.scala 82:228:@20595.4]
  assign _T_730 = io_wPort_3_en_0 & _T_729; // @[MemPrimitives.scala 83:102:@20596.4]
  assign _T_732 = {_T_724,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20598.4]
  assign _T_734 = {_T_730,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20600.4]
  assign _T_735 = _T_724 ? _T_732 : _T_734; // @[Mux.scala 31:69:@20601.4]
  assign _T_742 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@20609.4]
  assign _T_743 = _T_700 & _T_742; // @[MemPrimitives.scala 82:228:@20610.4]
  assign _T_744 = io_wPort_0_en_0 & _T_743; // @[MemPrimitives.scala 83:102:@20611.4]
  assign _T_748 = io_wPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@20613.4]
  assign _T_749 = _T_706 & _T_748; // @[MemPrimitives.scala 82:228:@20614.4]
  assign _T_750 = io_wPort_2_en_0 & _T_749; // @[MemPrimitives.scala 83:102:@20615.4]
  assign _T_752 = {_T_744,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20617.4]
  assign _T_754 = {_T_750,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20619.4]
  assign _T_755 = _T_744 ? _T_752 : _T_754; // @[Mux.scala 31:69:@20620.4]
  assign _T_762 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@20628.4]
  assign _T_763 = _T_720 & _T_762; // @[MemPrimitives.scala 82:228:@20629.4]
  assign _T_764 = io_wPort_1_en_0 & _T_763; // @[MemPrimitives.scala 83:102:@20630.4]
  assign _T_768 = io_wPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@20632.4]
  assign _T_769 = _T_726 & _T_768; // @[MemPrimitives.scala 82:228:@20633.4]
  assign _T_770 = io_wPort_3_en_0 & _T_769; // @[MemPrimitives.scala 83:102:@20634.4]
  assign _T_772 = {_T_764,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20636.4]
  assign _T_774 = {_T_770,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20638.4]
  assign _T_775 = _T_764 ? _T_772 : _T_774; // @[Mux.scala 31:69:@20639.4]
  assign _T_782 = io_wPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@20647.4]
  assign _T_783 = _T_700 & _T_782; // @[MemPrimitives.scala 82:228:@20648.4]
  assign _T_784 = io_wPort_0_en_0 & _T_783; // @[MemPrimitives.scala 83:102:@20649.4]
  assign _T_788 = io_wPort_2_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@20651.4]
  assign _T_789 = _T_706 & _T_788; // @[MemPrimitives.scala 82:228:@20652.4]
  assign _T_790 = io_wPort_2_en_0 & _T_789; // @[MemPrimitives.scala 83:102:@20653.4]
  assign _T_792 = {_T_784,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20655.4]
  assign _T_794 = {_T_790,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20657.4]
  assign _T_795 = _T_784 ? _T_792 : _T_794; // @[Mux.scala 31:69:@20658.4]
  assign _T_802 = io_wPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@20666.4]
  assign _T_803 = _T_720 & _T_802; // @[MemPrimitives.scala 82:228:@20667.4]
  assign _T_804 = io_wPort_1_en_0 & _T_803; // @[MemPrimitives.scala 83:102:@20668.4]
  assign _T_808 = io_wPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@20670.4]
  assign _T_809 = _T_726 & _T_808; // @[MemPrimitives.scala 82:228:@20671.4]
  assign _T_810 = io_wPort_3_en_0 & _T_809; // @[MemPrimitives.scala 83:102:@20672.4]
  assign _T_812 = {_T_804,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20674.4]
  assign _T_814 = {_T_810,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20676.4]
  assign _T_815 = _T_804 ? _T_812 : _T_814; // @[Mux.scala 31:69:@20677.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20684.4]
  assign _T_823 = _T_820 & _T_702; // @[MemPrimitives.scala 82:228:@20686.4]
  assign _T_824 = io_wPort_0_en_0 & _T_823; // @[MemPrimitives.scala 83:102:@20687.4]
  assign _T_826 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20688.4]
  assign _T_829 = _T_826 & _T_708; // @[MemPrimitives.scala 82:228:@20690.4]
  assign _T_830 = io_wPort_2_en_0 & _T_829; // @[MemPrimitives.scala 83:102:@20691.4]
  assign _T_832 = {_T_824,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20693.4]
  assign _T_834 = {_T_830,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20695.4]
  assign _T_835 = _T_824 ? _T_832 : _T_834; // @[Mux.scala 31:69:@20696.4]
  assign _T_840 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20703.4]
  assign _T_843 = _T_840 & _T_722; // @[MemPrimitives.scala 82:228:@20705.4]
  assign _T_844 = io_wPort_1_en_0 & _T_843; // @[MemPrimitives.scala 83:102:@20706.4]
  assign _T_846 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20707.4]
  assign _T_849 = _T_846 & _T_728; // @[MemPrimitives.scala 82:228:@20709.4]
  assign _T_850 = io_wPort_3_en_0 & _T_849; // @[MemPrimitives.scala 83:102:@20710.4]
  assign _T_852 = {_T_844,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20712.4]
  assign _T_854 = {_T_850,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20714.4]
  assign _T_855 = _T_844 ? _T_852 : _T_854; // @[Mux.scala 31:69:@20715.4]
  assign _T_863 = _T_820 & _T_742; // @[MemPrimitives.scala 82:228:@20724.4]
  assign _T_864 = io_wPort_0_en_0 & _T_863; // @[MemPrimitives.scala 83:102:@20725.4]
  assign _T_869 = _T_826 & _T_748; // @[MemPrimitives.scala 82:228:@20728.4]
  assign _T_870 = io_wPort_2_en_0 & _T_869; // @[MemPrimitives.scala 83:102:@20729.4]
  assign _T_872 = {_T_864,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20731.4]
  assign _T_874 = {_T_870,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20733.4]
  assign _T_875 = _T_864 ? _T_872 : _T_874; // @[Mux.scala 31:69:@20734.4]
  assign _T_883 = _T_840 & _T_762; // @[MemPrimitives.scala 82:228:@20743.4]
  assign _T_884 = io_wPort_1_en_0 & _T_883; // @[MemPrimitives.scala 83:102:@20744.4]
  assign _T_889 = _T_846 & _T_768; // @[MemPrimitives.scala 82:228:@20747.4]
  assign _T_890 = io_wPort_3_en_0 & _T_889; // @[MemPrimitives.scala 83:102:@20748.4]
  assign _T_892 = {_T_884,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20750.4]
  assign _T_894 = {_T_890,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20752.4]
  assign _T_895 = _T_884 ? _T_892 : _T_894; // @[Mux.scala 31:69:@20753.4]
  assign _T_903 = _T_820 & _T_782; // @[MemPrimitives.scala 82:228:@20762.4]
  assign _T_904 = io_wPort_0_en_0 & _T_903; // @[MemPrimitives.scala 83:102:@20763.4]
  assign _T_909 = _T_826 & _T_788; // @[MemPrimitives.scala 82:228:@20766.4]
  assign _T_910 = io_wPort_2_en_0 & _T_909; // @[MemPrimitives.scala 83:102:@20767.4]
  assign _T_912 = {_T_904,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20769.4]
  assign _T_914 = {_T_910,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20771.4]
  assign _T_915 = _T_904 ? _T_912 : _T_914; // @[Mux.scala 31:69:@20772.4]
  assign _T_923 = _T_840 & _T_802; // @[MemPrimitives.scala 82:228:@20781.4]
  assign _T_924 = io_wPort_1_en_0 & _T_923; // @[MemPrimitives.scala 83:102:@20782.4]
  assign _T_929 = _T_846 & _T_808; // @[MemPrimitives.scala 82:228:@20785.4]
  assign _T_930 = io_wPort_3_en_0 & _T_929; // @[MemPrimitives.scala 83:102:@20786.4]
  assign _T_932 = {_T_924,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20788.4]
  assign _T_934 = {_T_930,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20790.4]
  assign _T_935 = _T_924 ? _T_932 : _T_934; // @[Mux.scala 31:69:@20791.4]
  assign _T_940 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20798.4]
  assign _T_943 = _T_940 & _T_702; // @[MemPrimitives.scala 82:228:@20800.4]
  assign _T_944 = io_wPort_0_en_0 & _T_943; // @[MemPrimitives.scala 83:102:@20801.4]
  assign _T_946 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20802.4]
  assign _T_949 = _T_946 & _T_708; // @[MemPrimitives.scala 82:228:@20804.4]
  assign _T_950 = io_wPort_2_en_0 & _T_949; // @[MemPrimitives.scala 83:102:@20805.4]
  assign _T_952 = {_T_944,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20807.4]
  assign _T_954 = {_T_950,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20809.4]
  assign _T_955 = _T_944 ? _T_952 : _T_954; // @[Mux.scala 31:69:@20810.4]
  assign _T_960 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20817.4]
  assign _T_963 = _T_960 & _T_722; // @[MemPrimitives.scala 82:228:@20819.4]
  assign _T_964 = io_wPort_1_en_0 & _T_963; // @[MemPrimitives.scala 83:102:@20820.4]
  assign _T_966 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20821.4]
  assign _T_969 = _T_966 & _T_728; // @[MemPrimitives.scala 82:228:@20823.4]
  assign _T_970 = io_wPort_3_en_0 & _T_969; // @[MemPrimitives.scala 83:102:@20824.4]
  assign _T_972 = {_T_964,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20826.4]
  assign _T_974 = {_T_970,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20828.4]
  assign _T_975 = _T_964 ? _T_972 : _T_974; // @[Mux.scala 31:69:@20829.4]
  assign _T_983 = _T_940 & _T_742; // @[MemPrimitives.scala 82:228:@20838.4]
  assign _T_984 = io_wPort_0_en_0 & _T_983; // @[MemPrimitives.scala 83:102:@20839.4]
  assign _T_989 = _T_946 & _T_748; // @[MemPrimitives.scala 82:228:@20842.4]
  assign _T_990 = io_wPort_2_en_0 & _T_989; // @[MemPrimitives.scala 83:102:@20843.4]
  assign _T_992 = {_T_984,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20845.4]
  assign _T_994 = {_T_990,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20847.4]
  assign _T_995 = _T_984 ? _T_992 : _T_994; // @[Mux.scala 31:69:@20848.4]
  assign _T_1003 = _T_960 & _T_762; // @[MemPrimitives.scala 82:228:@20857.4]
  assign _T_1004 = io_wPort_1_en_0 & _T_1003; // @[MemPrimitives.scala 83:102:@20858.4]
  assign _T_1009 = _T_966 & _T_768; // @[MemPrimitives.scala 82:228:@20861.4]
  assign _T_1010 = io_wPort_3_en_0 & _T_1009; // @[MemPrimitives.scala 83:102:@20862.4]
  assign _T_1012 = {_T_1004,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20864.4]
  assign _T_1014 = {_T_1010,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20866.4]
  assign _T_1015 = _T_1004 ? _T_1012 : _T_1014; // @[Mux.scala 31:69:@20867.4]
  assign _T_1023 = _T_940 & _T_782; // @[MemPrimitives.scala 82:228:@20876.4]
  assign _T_1024 = io_wPort_0_en_0 & _T_1023; // @[MemPrimitives.scala 83:102:@20877.4]
  assign _T_1029 = _T_946 & _T_788; // @[MemPrimitives.scala 82:228:@20880.4]
  assign _T_1030 = io_wPort_2_en_0 & _T_1029; // @[MemPrimitives.scala 83:102:@20881.4]
  assign _T_1032 = {_T_1024,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20883.4]
  assign _T_1034 = {_T_1030,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20885.4]
  assign _T_1035 = _T_1024 ? _T_1032 : _T_1034; // @[Mux.scala 31:69:@20886.4]
  assign _T_1043 = _T_960 & _T_802; // @[MemPrimitives.scala 82:228:@20895.4]
  assign _T_1044 = io_wPort_1_en_0 & _T_1043; // @[MemPrimitives.scala 83:102:@20896.4]
  assign _T_1049 = _T_966 & _T_808; // @[MemPrimitives.scala 82:228:@20899.4]
  assign _T_1050 = io_wPort_3_en_0 & _T_1049; // @[MemPrimitives.scala 83:102:@20900.4]
  assign _T_1052 = {_T_1044,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20902.4]
  assign _T_1054 = {_T_1050,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20904.4]
  assign _T_1055 = _T_1044 ? _T_1052 : _T_1054; // @[Mux.scala 31:69:@20905.4]
  assign _T_1060 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20912.4]
  assign _T_1063 = _T_1060 & _T_702; // @[MemPrimitives.scala 82:228:@20914.4]
  assign _T_1064 = io_wPort_0_en_0 & _T_1063; // @[MemPrimitives.scala 83:102:@20915.4]
  assign _T_1066 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20916.4]
  assign _T_1069 = _T_1066 & _T_708; // @[MemPrimitives.scala 82:228:@20918.4]
  assign _T_1070 = io_wPort_2_en_0 & _T_1069; // @[MemPrimitives.scala 83:102:@20919.4]
  assign _T_1072 = {_T_1064,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20921.4]
  assign _T_1074 = {_T_1070,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20923.4]
  assign _T_1075 = _T_1064 ? _T_1072 : _T_1074; // @[Mux.scala 31:69:@20924.4]
  assign _T_1080 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20931.4]
  assign _T_1083 = _T_1080 & _T_722; // @[MemPrimitives.scala 82:228:@20933.4]
  assign _T_1084 = io_wPort_1_en_0 & _T_1083; // @[MemPrimitives.scala 83:102:@20934.4]
  assign _T_1086 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20935.4]
  assign _T_1089 = _T_1086 & _T_728; // @[MemPrimitives.scala 82:228:@20937.4]
  assign _T_1090 = io_wPort_3_en_0 & _T_1089; // @[MemPrimitives.scala 83:102:@20938.4]
  assign _T_1092 = {_T_1084,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20940.4]
  assign _T_1094 = {_T_1090,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20942.4]
  assign _T_1095 = _T_1084 ? _T_1092 : _T_1094; // @[Mux.scala 31:69:@20943.4]
  assign _T_1103 = _T_1060 & _T_742; // @[MemPrimitives.scala 82:228:@20952.4]
  assign _T_1104 = io_wPort_0_en_0 & _T_1103; // @[MemPrimitives.scala 83:102:@20953.4]
  assign _T_1109 = _T_1066 & _T_748; // @[MemPrimitives.scala 82:228:@20956.4]
  assign _T_1110 = io_wPort_2_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@20957.4]
  assign _T_1112 = {_T_1104,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20959.4]
  assign _T_1114 = {_T_1110,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20961.4]
  assign _T_1115 = _T_1104 ? _T_1112 : _T_1114; // @[Mux.scala 31:69:@20962.4]
  assign _T_1123 = _T_1080 & _T_762; // @[MemPrimitives.scala 82:228:@20971.4]
  assign _T_1124 = io_wPort_1_en_0 & _T_1123; // @[MemPrimitives.scala 83:102:@20972.4]
  assign _T_1129 = _T_1086 & _T_768; // @[MemPrimitives.scala 82:228:@20975.4]
  assign _T_1130 = io_wPort_3_en_0 & _T_1129; // @[MemPrimitives.scala 83:102:@20976.4]
  assign _T_1132 = {_T_1124,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20978.4]
  assign _T_1134 = {_T_1130,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20980.4]
  assign _T_1135 = _T_1124 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@20981.4]
  assign _T_1143 = _T_1060 & _T_782; // @[MemPrimitives.scala 82:228:@20990.4]
  assign _T_1144 = io_wPort_0_en_0 & _T_1143; // @[MemPrimitives.scala 83:102:@20991.4]
  assign _T_1149 = _T_1066 & _T_788; // @[MemPrimitives.scala 82:228:@20994.4]
  assign _T_1150 = io_wPort_2_en_0 & _T_1149; // @[MemPrimitives.scala 83:102:@20995.4]
  assign _T_1152 = {_T_1144,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20997.4]
  assign _T_1154 = {_T_1150,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20999.4]
  assign _T_1155 = _T_1144 ? _T_1152 : _T_1154; // @[Mux.scala 31:69:@21000.4]
  assign _T_1163 = _T_1080 & _T_802; // @[MemPrimitives.scala 82:228:@21009.4]
  assign _T_1164 = io_wPort_1_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@21010.4]
  assign _T_1169 = _T_1086 & _T_808; // @[MemPrimitives.scala 82:228:@21013.4]
  assign _T_1170 = io_wPort_3_en_0 & _T_1169; // @[MemPrimitives.scala 83:102:@21014.4]
  assign _T_1172 = {_T_1164,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@21016.4]
  assign _T_1174 = {_T_1170,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@21018.4]
  assign _T_1175 = _T_1164 ? _T_1172 : _T_1174; // @[Mux.scala 31:69:@21019.4]
  assign _T_1180 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21026.4]
  assign _T_1182 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21027.4]
  assign _T_1183 = _T_1180 & _T_1182; // @[MemPrimitives.scala 110:228:@21028.4]
  assign _T_1186 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21030.4]
  assign _T_1188 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21031.4]
  assign _T_1189 = _T_1186 & _T_1188; // @[MemPrimitives.scala 110:228:@21032.4]
  assign _T_1192 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21034.4]
  assign _T_1194 = io_rPort_5_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21035.4]
  assign _T_1195 = _T_1192 & _T_1194; // @[MemPrimitives.scala 110:228:@21036.4]
  assign _T_1198 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21038.4]
  assign _T_1200 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21039.4]
  assign _T_1201 = _T_1198 & _T_1200; // @[MemPrimitives.scala 110:228:@21040.4]
  assign _T_1204 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21042.4]
  assign _T_1206 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21043.4]
  assign _T_1207 = _T_1204 & _T_1206; // @[MemPrimitives.scala 110:228:@21044.4]
  assign _T_1210 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21046.4]
  assign _T_1212 = io_rPort_9_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21047.4]
  assign _T_1213 = _T_1210 & _T_1212; // @[MemPrimitives.scala 110:228:@21048.4]
  assign _T_1216 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21050.4]
  assign _T_1218 = io_rPort_11_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21051.4]
  assign _T_1219 = _T_1216 & _T_1218; // @[MemPrimitives.scala 110:228:@21052.4]
  assign _T_1222 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21054.4]
  assign _T_1224 = io_rPort_14_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21055.4]
  assign _T_1225 = _T_1222 & _T_1224; // @[MemPrimitives.scala 110:228:@21056.4]
  assign _T_1228 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21058.4]
  assign _T_1230 = io_rPort_16_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21059.4]
  assign _T_1231 = _T_1228 & _T_1230; // @[MemPrimitives.scala 110:228:@21060.4]
  assign _T_1233 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@21074.4]
  assign _T_1234 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@21075.4]
  assign _T_1235 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@21076.4]
  assign _T_1236 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@21077.4]
  assign _T_1237 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@21078.4]
  assign _T_1238 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@21079.4]
  assign _T_1239 = StickySelects_io_outs_6; // @[MemPrimitives.scala 126:35:@21080.4]
  assign _T_1240 = StickySelects_io_outs_7; // @[MemPrimitives.scala 126:35:@21081.4]
  assign _T_1241 = StickySelects_io_outs_8; // @[MemPrimitives.scala 126:35:@21082.4]
  assign _T_1243 = {_T_1233,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21084.4]
  assign _T_1245 = {_T_1234,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21086.4]
  assign _T_1247 = {_T_1235,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21088.4]
  assign _T_1249 = {_T_1236,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21090.4]
  assign _T_1251 = {_T_1237,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21092.4]
  assign _T_1253 = {_T_1238,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21094.4]
  assign _T_1255 = {_T_1239,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21096.4]
  assign _T_1257 = {_T_1240,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21098.4]
  assign _T_1259 = {_T_1241,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21100.4]
  assign _T_1260 = _T_1240 ? _T_1257 : _T_1259; // @[Mux.scala 31:69:@21101.4]
  assign _T_1261 = _T_1239 ? _T_1255 : _T_1260; // @[Mux.scala 31:69:@21102.4]
  assign _T_1262 = _T_1238 ? _T_1253 : _T_1261; // @[Mux.scala 31:69:@21103.4]
  assign _T_1263 = _T_1237 ? _T_1251 : _T_1262; // @[Mux.scala 31:69:@21104.4]
  assign _T_1264 = _T_1236 ? _T_1249 : _T_1263; // @[Mux.scala 31:69:@21105.4]
  assign _T_1265 = _T_1235 ? _T_1247 : _T_1264; // @[Mux.scala 31:69:@21106.4]
  assign _T_1266 = _T_1234 ? _T_1245 : _T_1265; // @[Mux.scala 31:69:@21107.4]
  assign _T_1267 = _T_1233 ? _T_1243 : _T_1266; // @[Mux.scala 31:69:@21108.4]
  assign _T_1272 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21115.4]
  assign _T_1274 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21116.4]
  assign _T_1275 = _T_1272 & _T_1274; // @[MemPrimitives.scala 110:228:@21117.4]
  assign _T_1278 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21119.4]
  assign _T_1280 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21120.4]
  assign _T_1281 = _T_1278 & _T_1280; // @[MemPrimitives.scala 110:228:@21121.4]
  assign _T_1284 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21123.4]
  assign _T_1286 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21124.4]
  assign _T_1287 = _T_1284 & _T_1286; // @[MemPrimitives.scala 110:228:@21125.4]
  assign _T_1290 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21127.4]
  assign _T_1292 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21128.4]
  assign _T_1293 = _T_1290 & _T_1292; // @[MemPrimitives.scala 110:228:@21129.4]
  assign _T_1296 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21131.4]
  assign _T_1298 = io_rPort_10_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21132.4]
  assign _T_1299 = _T_1296 & _T_1298; // @[MemPrimitives.scala 110:228:@21133.4]
  assign _T_1302 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21135.4]
  assign _T_1304 = io_rPort_12_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21136.4]
  assign _T_1305 = _T_1302 & _T_1304; // @[MemPrimitives.scala 110:228:@21137.4]
  assign _T_1308 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21139.4]
  assign _T_1310 = io_rPort_13_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21140.4]
  assign _T_1311 = _T_1308 & _T_1310; // @[MemPrimitives.scala 110:228:@21141.4]
  assign _T_1314 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21143.4]
  assign _T_1316 = io_rPort_15_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21144.4]
  assign _T_1317 = _T_1314 & _T_1316; // @[MemPrimitives.scala 110:228:@21145.4]
  assign _T_1320 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21147.4]
  assign _T_1322 = io_rPort_17_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21148.4]
  assign _T_1323 = _T_1320 & _T_1322; // @[MemPrimitives.scala 110:228:@21149.4]
  assign _T_1325 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@21163.4]
  assign _T_1326 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@21164.4]
  assign _T_1327 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@21165.4]
  assign _T_1328 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@21166.4]
  assign _T_1329 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@21167.4]
  assign _T_1330 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@21168.4]
  assign _T_1331 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 126:35:@21169.4]
  assign _T_1332 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 126:35:@21170.4]
  assign _T_1333 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 126:35:@21171.4]
  assign _T_1335 = {_T_1325,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21173.4]
  assign _T_1337 = {_T_1326,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21175.4]
  assign _T_1339 = {_T_1327,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21177.4]
  assign _T_1341 = {_T_1328,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21179.4]
  assign _T_1343 = {_T_1329,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21181.4]
  assign _T_1345 = {_T_1330,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21183.4]
  assign _T_1347 = {_T_1331,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21185.4]
  assign _T_1349 = {_T_1332,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21187.4]
  assign _T_1351 = {_T_1333,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21189.4]
  assign _T_1352 = _T_1332 ? _T_1349 : _T_1351; // @[Mux.scala 31:69:@21190.4]
  assign _T_1353 = _T_1331 ? _T_1347 : _T_1352; // @[Mux.scala 31:69:@21191.4]
  assign _T_1354 = _T_1330 ? _T_1345 : _T_1353; // @[Mux.scala 31:69:@21192.4]
  assign _T_1355 = _T_1329 ? _T_1343 : _T_1354; // @[Mux.scala 31:69:@21193.4]
  assign _T_1356 = _T_1328 ? _T_1341 : _T_1355; // @[Mux.scala 31:69:@21194.4]
  assign _T_1357 = _T_1327 ? _T_1339 : _T_1356; // @[Mux.scala 31:69:@21195.4]
  assign _T_1358 = _T_1326 ? _T_1337 : _T_1357; // @[Mux.scala 31:69:@21196.4]
  assign _T_1359 = _T_1325 ? _T_1335 : _T_1358; // @[Mux.scala 31:69:@21197.4]
  assign _T_1366 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21205.4]
  assign _T_1367 = _T_1180 & _T_1366; // @[MemPrimitives.scala 110:228:@21206.4]
  assign _T_1372 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21209.4]
  assign _T_1373 = _T_1186 & _T_1372; // @[MemPrimitives.scala 110:228:@21210.4]
  assign _T_1378 = io_rPort_5_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21213.4]
  assign _T_1379 = _T_1192 & _T_1378; // @[MemPrimitives.scala 110:228:@21214.4]
  assign _T_1384 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21217.4]
  assign _T_1385 = _T_1198 & _T_1384; // @[MemPrimitives.scala 110:228:@21218.4]
  assign _T_1390 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21221.4]
  assign _T_1391 = _T_1204 & _T_1390; // @[MemPrimitives.scala 110:228:@21222.4]
  assign _T_1396 = io_rPort_9_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21225.4]
  assign _T_1397 = _T_1210 & _T_1396; // @[MemPrimitives.scala 110:228:@21226.4]
  assign _T_1402 = io_rPort_11_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21229.4]
  assign _T_1403 = _T_1216 & _T_1402; // @[MemPrimitives.scala 110:228:@21230.4]
  assign _T_1408 = io_rPort_14_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21233.4]
  assign _T_1409 = _T_1222 & _T_1408; // @[MemPrimitives.scala 110:228:@21234.4]
  assign _T_1414 = io_rPort_16_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21237.4]
  assign _T_1415 = _T_1228 & _T_1414; // @[MemPrimitives.scala 110:228:@21238.4]
  assign _T_1417 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@21252.4]
  assign _T_1418 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@21253.4]
  assign _T_1419 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@21254.4]
  assign _T_1420 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@21255.4]
  assign _T_1421 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@21256.4]
  assign _T_1422 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@21257.4]
  assign _T_1423 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 126:35:@21258.4]
  assign _T_1424 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 126:35:@21259.4]
  assign _T_1425 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 126:35:@21260.4]
  assign _T_1427 = {_T_1417,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21262.4]
  assign _T_1429 = {_T_1418,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21264.4]
  assign _T_1431 = {_T_1419,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21266.4]
  assign _T_1433 = {_T_1420,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21268.4]
  assign _T_1435 = {_T_1421,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21270.4]
  assign _T_1437 = {_T_1422,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21272.4]
  assign _T_1439 = {_T_1423,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21274.4]
  assign _T_1441 = {_T_1424,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21276.4]
  assign _T_1443 = {_T_1425,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21278.4]
  assign _T_1444 = _T_1424 ? _T_1441 : _T_1443; // @[Mux.scala 31:69:@21279.4]
  assign _T_1445 = _T_1423 ? _T_1439 : _T_1444; // @[Mux.scala 31:69:@21280.4]
  assign _T_1446 = _T_1422 ? _T_1437 : _T_1445; // @[Mux.scala 31:69:@21281.4]
  assign _T_1447 = _T_1421 ? _T_1435 : _T_1446; // @[Mux.scala 31:69:@21282.4]
  assign _T_1448 = _T_1420 ? _T_1433 : _T_1447; // @[Mux.scala 31:69:@21283.4]
  assign _T_1449 = _T_1419 ? _T_1431 : _T_1448; // @[Mux.scala 31:69:@21284.4]
  assign _T_1450 = _T_1418 ? _T_1429 : _T_1449; // @[Mux.scala 31:69:@21285.4]
  assign _T_1451 = _T_1417 ? _T_1427 : _T_1450; // @[Mux.scala 31:69:@21286.4]
  assign _T_1458 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21294.4]
  assign _T_1459 = _T_1272 & _T_1458; // @[MemPrimitives.scala 110:228:@21295.4]
  assign _T_1464 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21298.4]
  assign _T_1465 = _T_1278 & _T_1464; // @[MemPrimitives.scala 110:228:@21299.4]
  assign _T_1470 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21302.4]
  assign _T_1471 = _T_1284 & _T_1470; // @[MemPrimitives.scala 110:228:@21303.4]
  assign _T_1476 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21306.4]
  assign _T_1477 = _T_1290 & _T_1476; // @[MemPrimitives.scala 110:228:@21307.4]
  assign _T_1482 = io_rPort_10_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21310.4]
  assign _T_1483 = _T_1296 & _T_1482; // @[MemPrimitives.scala 110:228:@21311.4]
  assign _T_1488 = io_rPort_12_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21314.4]
  assign _T_1489 = _T_1302 & _T_1488; // @[MemPrimitives.scala 110:228:@21315.4]
  assign _T_1494 = io_rPort_13_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21318.4]
  assign _T_1495 = _T_1308 & _T_1494; // @[MemPrimitives.scala 110:228:@21319.4]
  assign _T_1500 = io_rPort_15_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21322.4]
  assign _T_1501 = _T_1314 & _T_1500; // @[MemPrimitives.scala 110:228:@21323.4]
  assign _T_1506 = io_rPort_17_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21326.4]
  assign _T_1507 = _T_1320 & _T_1506; // @[MemPrimitives.scala 110:228:@21327.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@21341.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@21342.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@21343.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@21344.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@21345.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@21346.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 126:35:@21347.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 126:35:@21348.4]
  assign _T_1517 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 126:35:@21349.4]
  assign _T_1519 = {_T_1509,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21351.4]
  assign _T_1521 = {_T_1510,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21353.4]
  assign _T_1523 = {_T_1511,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21355.4]
  assign _T_1525 = {_T_1512,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21357.4]
  assign _T_1527 = {_T_1513,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21359.4]
  assign _T_1529 = {_T_1514,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21361.4]
  assign _T_1531 = {_T_1515,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21363.4]
  assign _T_1533 = {_T_1516,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21365.4]
  assign _T_1535 = {_T_1517,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21367.4]
  assign _T_1536 = _T_1516 ? _T_1533 : _T_1535; // @[Mux.scala 31:69:@21368.4]
  assign _T_1537 = _T_1515 ? _T_1531 : _T_1536; // @[Mux.scala 31:69:@21369.4]
  assign _T_1538 = _T_1514 ? _T_1529 : _T_1537; // @[Mux.scala 31:69:@21370.4]
  assign _T_1539 = _T_1513 ? _T_1527 : _T_1538; // @[Mux.scala 31:69:@21371.4]
  assign _T_1540 = _T_1512 ? _T_1525 : _T_1539; // @[Mux.scala 31:69:@21372.4]
  assign _T_1541 = _T_1511 ? _T_1523 : _T_1540; // @[Mux.scala 31:69:@21373.4]
  assign _T_1542 = _T_1510 ? _T_1521 : _T_1541; // @[Mux.scala 31:69:@21374.4]
  assign _T_1543 = _T_1509 ? _T_1519 : _T_1542; // @[Mux.scala 31:69:@21375.4]
  assign _T_1550 = io_rPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21383.4]
  assign _T_1551 = _T_1180 & _T_1550; // @[MemPrimitives.scala 110:228:@21384.4]
  assign _T_1556 = io_rPort_1_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21387.4]
  assign _T_1557 = _T_1186 & _T_1556; // @[MemPrimitives.scala 110:228:@21388.4]
  assign _T_1562 = io_rPort_5_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21391.4]
  assign _T_1563 = _T_1192 & _T_1562; // @[MemPrimitives.scala 110:228:@21392.4]
  assign _T_1568 = io_rPort_7_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21395.4]
  assign _T_1569 = _T_1198 & _T_1568; // @[MemPrimitives.scala 110:228:@21396.4]
  assign _T_1574 = io_rPort_8_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21399.4]
  assign _T_1575 = _T_1204 & _T_1574; // @[MemPrimitives.scala 110:228:@21400.4]
  assign _T_1580 = io_rPort_9_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21403.4]
  assign _T_1581 = _T_1210 & _T_1580; // @[MemPrimitives.scala 110:228:@21404.4]
  assign _T_1586 = io_rPort_11_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21407.4]
  assign _T_1587 = _T_1216 & _T_1586; // @[MemPrimitives.scala 110:228:@21408.4]
  assign _T_1592 = io_rPort_14_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21411.4]
  assign _T_1593 = _T_1222 & _T_1592; // @[MemPrimitives.scala 110:228:@21412.4]
  assign _T_1598 = io_rPort_16_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21415.4]
  assign _T_1599 = _T_1228 & _T_1598; // @[MemPrimitives.scala 110:228:@21416.4]
  assign _T_1601 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@21430.4]
  assign _T_1602 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@21431.4]
  assign _T_1603 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@21432.4]
  assign _T_1604 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@21433.4]
  assign _T_1605 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@21434.4]
  assign _T_1606 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@21435.4]
  assign _T_1607 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 126:35:@21436.4]
  assign _T_1608 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 126:35:@21437.4]
  assign _T_1609 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 126:35:@21438.4]
  assign _T_1611 = {_T_1601,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21440.4]
  assign _T_1613 = {_T_1602,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21442.4]
  assign _T_1615 = {_T_1603,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21444.4]
  assign _T_1617 = {_T_1604,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21446.4]
  assign _T_1619 = {_T_1605,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21448.4]
  assign _T_1621 = {_T_1606,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21450.4]
  assign _T_1623 = {_T_1607,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21452.4]
  assign _T_1625 = {_T_1608,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21454.4]
  assign _T_1627 = {_T_1609,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21456.4]
  assign _T_1628 = _T_1608 ? _T_1625 : _T_1627; // @[Mux.scala 31:69:@21457.4]
  assign _T_1629 = _T_1607 ? _T_1623 : _T_1628; // @[Mux.scala 31:69:@21458.4]
  assign _T_1630 = _T_1606 ? _T_1621 : _T_1629; // @[Mux.scala 31:69:@21459.4]
  assign _T_1631 = _T_1605 ? _T_1619 : _T_1630; // @[Mux.scala 31:69:@21460.4]
  assign _T_1632 = _T_1604 ? _T_1617 : _T_1631; // @[Mux.scala 31:69:@21461.4]
  assign _T_1633 = _T_1603 ? _T_1615 : _T_1632; // @[Mux.scala 31:69:@21462.4]
  assign _T_1634 = _T_1602 ? _T_1613 : _T_1633; // @[Mux.scala 31:69:@21463.4]
  assign _T_1635 = _T_1601 ? _T_1611 : _T_1634; // @[Mux.scala 31:69:@21464.4]
  assign _T_1642 = io_rPort_2_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21472.4]
  assign _T_1643 = _T_1272 & _T_1642; // @[MemPrimitives.scala 110:228:@21473.4]
  assign _T_1648 = io_rPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21476.4]
  assign _T_1649 = _T_1278 & _T_1648; // @[MemPrimitives.scala 110:228:@21477.4]
  assign _T_1654 = io_rPort_4_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21480.4]
  assign _T_1655 = _T_1284 & _T_1654; // @[MemPrimitives.scala 110:228:@21481.4]
  assign _T_1660 = io_rPort_6_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21484.4]
  assign _T_1661 = _T_1290 & _T_1660; // @[MemPrimitives.scala 110:228:@21485.4]
  assign _T_1666 = io_rPort_10_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21488.4]
  assign _T_1667 = _T_1296 & _T_1666; // @[MemPrimitives.scala 110:228:@21489.4]
  assign _T_1672 = io_rPort_12_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21492.4]
  assign _T_1673 = _T_1302 & _T_1672; // @[MemPrimitives.scala 110:228:@21493.4]
  assign _T_1678 = io_rPort_13_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21496.4]
  assign _T_1679 = _T_1308 & _T_1678; // @[MemPrimitives.scala 110:228:@21497.4]
  assign _T_1684 = io_rPort_15_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21500.4]
  assign _T_1685 = _T_1314 & _T_1684; // @[MemPrimitives.scala 110:228:@21501.4]
  assign _T_1690 = io_rPort_17_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21504.4]
  assign _T_1691 = _T_1320 & _T_1690; // @[MemPrimitives.scala 110:228:@21505.4]
  assign _T_1693 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@21519.4]
  assign _T_1694 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@21520.4]
  assign _T_1695 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@21521.4]
  assign _T_1696 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@21522.4]
  assign _T_1697 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@21523.4]
  assign _T_1698 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@21524.4]
  assign _T_1699 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 126:35:@21525.4]
  assign _T_1700 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 126:35:@21526.4]
  assign _T_1701 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 126:35:@21527.4]
  assign _T_1703 = {_T_1693,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21529.4]
  assign _T_1705 = {_T_1694,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21531.4]
  assign _T_1707 = {_T_1695,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21533.4]
  assign _T_1709 = {_T_1696,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21535.4]
  assign _T_1711 = {_T_1697,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21537.4]
  assign _T_1713 = {_T_1698,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21539.4]
  assign _T_1715 = {_T_1699,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21541.4]
  assign _T_1717 = {_T_1700,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21543.4]
  assign _T_1719 = {_T_1701,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21545.4]
  assign _T_1720 = _T_1700 ? _T_1717 : _T_1719; // @[Mux.scala 31:69:@21546.4]
  assign _T_1721 = _T_1699 ? _T_1715 : _T_1720; // @[Mux.scala 31:69:@21547.4]
  assign _T_1722 = _T_1698 ? _T_1713 : _T_1721; // @[Mux.scala 31:69:@21548.4]
  assign _T_1723 = _T_1697 ? _T_1711 : _T_1722; // @[Mux.scala 31:69:@21549.4]
  assign _T_1724 = _T_1696 ? _T_1709 : _T_1723; // @[Mux.scala 31:69:@21550.4]
  assign _T_1725 = _T_1695 ? _T_1707 : _T_1724; // @[Mux.scala 31:69:@21551.4]
  assign _T_1726 = _T_1694 ? _T_1705 : _T_1725; // @[Mux.scala 31:69:@21552.4]
  assign _T_1727 = _T_1693 ? _T_1703 : _T_1726; // @[Mux.scala 31:69:@21553.4]
  assign _T_1732 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21560.4]
  assign _T_1735 = _T_1732 & _T_1182; // @[MemPrimitives.scala 110:228:@21562.4]
  assign _T_1738 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21564.4]
  assign _T_1741 = _T_1738 & _T_1188; // @[MemPrimitives.scala 110:228:@21566.4]
  assign _T_1744 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21568.4]
  assign _T_1747 = _T_1744 & _T_1194; // @[MemPrimitives.scala 110:228:@21570.4]
  assign _T_1750 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21572.4]
  assign _T_1753 = _T_1750 & _T_1200; // @[MemPrimitives.scala 110:228:@21574.4]
  assign _T_1756 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21576.4]
  assign _T_1759 = _T_1756 & _T_1206; // @[MemPrimitives.scala 110:228:@21578.4]
  assign _T_1762 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21580.4]
  assign _T_1765 = _T_1762 & _T_1212; // @[MemPrimitives.scala 110:228:@21582.4]
  assign _T_1768 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21584.4]
  assign _T_1771 = _T_1768 & _T_1218; // @[MemPrimitives.scala 110:228:@21586.4]
  assign _T_1774 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21588.4]
  assign _T_1777 = _T_1774 & _T_1224; // @[MemPrimitives.scala 110:228:@21590.4]
  assign _T_1780 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21592.4]
  assign _T_1783 = _T_1780 & _T_1230; // @[MemPrimitives.scala 110:228:@21594.4]
  assign _T_1785 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@21608.4]
  assign _T_1786 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@21609.4]
  assign _T_1787 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@21610.4]
  assign _T_1788 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@21611.4]
  assign _T_1789 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@21612.4]
  assign _T_1790 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@21613.4]
  assign _T_1791 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 126:35:@21614.4]
  assign _T_1792 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 126:35:@21615.4]
  assign _T_1793 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 126:35:@21616.4]
  assign _T_1795 = {_T_1785,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21618.4]
  assign _T_1797 = {_T_1786,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21620.4]
  assign _T_1799 = {_T_1787,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21622.4]
  assign _T_1801 = {_T_1788,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21624.4]
  assign _T_1803 = {_T_1789,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21626.4]
  assign _T_1805 = {_T_1790,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21628.4]
  assign _T_1807 = {_T_1791,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21630.4]
  assign _T_1809 = {_T_1792,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21632.4]
  assign _T_1811 = {_T_1793,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21634.4]
  assign _T_1812 = _T_1792 ? _T_1809 : _T_1811; // @[Mux.scala 31:69:@21635.4]
  assign _T_1813 = _T_1791 ? _T_1807 : _T_1812; // @[Mux.scala 31:69:@21636.4]
  assign _T_1814 = _T_1790 ? _T_1805 : _T_1813; // @[Mux.scala 31:69:@21637.4]
  assign _T_1815 = _T_1789 ? _T_1803 : _T_1814; // @[Mux.scala 31:69:@21638.4]
  assign _T_1816 = _T_1788 ? _T_1801 : _T_1815; // @[Mux.scala 31:69:@21639.4]
  assign _T_1817 = _T_1787 ? _T_1799 : _T_1816; // @[Mux.scala 31:69:@21640.4]
  assign _T_1818 = _T_1786 ? _T_1797 : _T_1817; // @[Mux.scala 31:69:@21641.4]
  assign _T_1819 = _T_1785 ? _T_1795 : _T_1818; // @[Mux.scala 31:69:@21642.4]
  assign _T_1824 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21649.4]
  assign _T_1827 = _T_1824 & _T_1274; // @[MemPrimitives.scala 110:228:@21651.4]
  assign _T_1830 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21653.4]
  assign _T_1833 = _T_1830 & _T_1280; // @[MemPrimitives.scala 110:228:@21655.4]
  assign _T_1836 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21657.4]
  assign _T_1839 = _T_1836 & _T_1286; // @[MemPrimitives.scala 110:228:@21659.4]
  assign _T_1842 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21661.4]
  assign _T_1845 = _T_1842 & _T_1292; // @[MemPrimitives.scala 110:228:@21663.4]
  assign _T_1848 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21665.4]
  assign _T_1851 = _T_1848 & _T_1298; // @[MemPrimitives.scala 110:228:@21667.4]
  assign _T_1854 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21669.4]
  assign _T_1857 = _T_1854 & _T_1304; // @[MemPrimitives.scala 110:228:@21671.4]
  assign _T_1860 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21673.4]
  assign _T_1863 = _T_1860 & _T_1310; // @[MemPrimitives.scala 110:228:@21675.4]
  assign _T_1866 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21677.4]
  assign _T_1869 = _T_1866 & _T_1316; // @[MemPrimitives.scala 110:228:@21679.4]
  assign _T_1872 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21681.4]
  assign _T_1875 = _T_1872 & _T_1322; // @[MemPrimitives.scala 110:228:@21683.4]
  assign _T_1877 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@21697.4]
  assign _T_1878 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@21698.4]
  assign _T_1879 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@21699.4]
  assign _T_1880 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@21700.4]
  assign _T_1881 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@21701.4]
  assign _T_1882 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@21702.4]
  assign _T_1883 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 126:35:@21703.4]
  assign _T_1884 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 126:35:@21704.4]
  assign _T_1885 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 126:35:@21705.4]
  assign _T_1887 = {_T_1877,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21707.4]
  assign _T_1889 = {_T_1878,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21709.4]
  assign _T_1891 = {_T_1879,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21711.4]
  assign _T_1893 = {_T_1880,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21713.4]
  assign _T_1895 = {_T_1881,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21715.4]
  assign _T_1897 = {_T_1882,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21717.4]
  assign _T_1899 = {_T_1883,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21719.4]
  assign _T_1901 = {_T_1884,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21721.4]
  assign _T_1903 = {_T_1885,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21723.4]
  assign _T_1904 = _T_1884 ? _T_1901 : _T_1903; // @[Mux.scala 31:69:@21724.4]
  assign _T_1905 = _T_1883 ? _T_1899 : _T_1904; // @[Mux.scala 31:69:@21725.4]
  assign _T_1906 = _T_1882 ? _T_1897 : _T_1905; // @[Mux.scala 31:69:@21726.4]
  assign _T_1907 = _T_1881 ? _T_1895 : _T_1906; // @[Mux.scala 31:69:@21727.4]
  assign _T_1908 = _T_1880 ? _T_1893 : _T_1907; // @[Mux.scala 31:69:@21728.4]
  assign _T_1909 = _T_1879 ? _T_1891 : _T_1908; // @[Mux.scala 31:69:@21729.4]
  assign _T_1910 = _T_1878 ? _T_1889 : _T_1909; // @[Mux.scala 31:69:@21730.4]
  assign _T_1911 = _T_1877 ? _T_1887 : _T_1910; // @[Mux.scala 31:69:@21731.4]
  assign _T_1919 = _T_1732 & _T_1366; // @[MemPrimitives.scala 110:228:@21740.4]
  assign _T_1925 = _T_1738 & _T_1372; // @[MemPrimitives.scala 110:228:@21744.4]
  assign _T_1931 = _T_1744 & _T_1378; // @[MemPrimitives.scala 110:228:@21748.4]
  assign _T_1937 = _T_1750 & _T_1384; // @[MemPrimitives.scala 110:228:@21752.4]
  assign _T_1943 = _T_1756 & _T_1390; // @[MemPrimitives.scala 110:228:@21756.4]
  assign _T_1949 = _T_1762 & _T_1396; // @[MemPrimitives.scala 110:228:@21760.4]
  assign _T_1955 = _T_1768 & _T_1402; // @[MemPrimitives.scala 110:228:@21764.4]
  assign _T_1961 = _T_1774 & _T_1408; // @[MemPrimitives.scala 110:228:@21768.4]
  assign _T_1967 = _T_1780 & _T_1414; // @[MemPrimitives.scala 110:228:@21772.4]
  assign _T_1969 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@21786.4]
  assign _T_1970 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@21787.4]
  assign _T_1971 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@21788.4]
  assign _T_1972 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@21789.4]
  assign _T_1973 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@21790.4]
  assign _T_1974 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@21791.4]
  assign _T_1975 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 126:35:@21792.4]
  assign _T_1976 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 126:35:@21793.4]
  assign _T_1977 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 126:35:@21794.4]
  assign _T_1979 = {_T_1969,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21796.4]
  assign _T_1981 = {_T_1970,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21798.4]
  assign _T_1983 = {_T_1971,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21800.4]
  assign _T_1985 = {_T_1972,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21802.4]
  assign _T_1987 = {_T_1973,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21804.4]
  assign _T_1989 = {_T_1974,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21806.4]
  assign _T_1991 = {_T_1975,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21808.4]
  assign _T_1993 = {_T_1976,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21810.4]
  assign _T_1995 = {_T_1977,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21812.4]
  assign _T_1996 = _T_1976 ? _T_1993 : _T_1995; // @[Mux.scala 31:69:@21813.4]
  assign _T_1997 = _T_1975 ? _T_1991 : _T_1996; // @[Mux.scala 31:69:@21814.4]
  assign _T_1998 = _T_1974 ? _T_1989 : _T_1997; // @[Mux.scala 31:69:@21815.4]
  assign _T_1999 = _T_1973 ? _T_1987 : _T_1998; // @[Mux.scala 31:69:@21816.4]
  assign _T_2000 = _T_1972 ? _T_1985 : _T_1999; // @[Mux.scala 31:69:@21817.4]
  assign _T_2001 = _T_1971 ? _T_1983 : _T_2000; // @[Mux.scala 31:69:@21818.4]
  assign _T_2002 = _T_1970 ? _T_1981 : _T_2001; // @[Mux.scala 31:69:@21819.4]
  assign _T_2003 = _T_1969 ? _T_1979 : _T_2002; // @[Mux.scala 31:69:@21820.4]
  assign _T_2011 = _T_1824 & _T_1458; // @[MemPrimitives.scala 110:228:@21829.4]
  assign _T_2017 = _T_1830 & _T_1464; // @[MemPrimitives.scala 110:228:@21833.4]
  assign _T_2023 = _T_1836 & _T_1470; // @[MemPrimitives.scala 110:228:@21837.4]
  assign _T_2029 = _T_1842 & _T_1476; // @[MemPrimitives.scala 110:228:@21841.4]
  assign _T_2035 = _T_1848 & _T_1482; // @[MemPrimitives.scala 110:228:@21845.4]
  assign _T_2041 = _T_1854 & _T_1488; // @[MemPrimitives.scala 110:228:@21849.4]
  assign _T_2047 = _T_1860 & _T_1494; // @[MemPrimitives.scala 110:228:@21853.4]
  assign _T_2053 = _T_1866 & _T_1500; // @[MemPrimitives.scala 110:228:@21857.4]
  assign _T_2059 = _T_1872 & _T_1506; // @[MemPrimitives.scala 110:228:@21861.4]
  assign _T_2061 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@21875.4]
  assign _T_2062 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@21876.4]
  assign _T_2063 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@21877.4]
  assign _T_2064 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@21878.4]
  assign _T_2065 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@21879.4]
  assign _T_2066 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@21880.4]
  assign _T_2067 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 126:35:@21881.4]
  assign _T_2068 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 126:35:@21882.4]
  assign _T_2069 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 126:35:@21883.4]
  assign _T_2071 = {_T_2061,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21885.4]
  assign _T_2073 = {_T_2062,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21887.4]
  assign _T_2075 = {_T_2063,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21889.4]
  assign _T_2077 = {_T_2064,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21891.4]
  assign _T_2079 = {_T_2065,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21893.4]
  assign _T_2081 = {_T_2066,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21895.4]
  assign _T_2083 = {_T_2067,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21897.4]
  assign _T_2085 = {_T_2068,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21899.4]
  assign _T_2087 = {_T_2069,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21901.4]
  assign _T_2088 = _T_2068 ? _T_2085 : _T_2087; // @[Mux.scala 31:69:@21902.4]
  assign _T_2089 = _T_2067 ? _T_2083 : _T_2088; // @[Mux.scala 31:69:@21903.4]
  assign _T_2090 = _T_2066 ? _T_2081 : _T_2089; // @[Mux.scala 31:69:@21904.4]
  assign _T_2091 = _T_2065 ? _T_2079 : _T_2090; // @[Mux.scala 31:69:@21905.4]
  assign _T_2092 = _T_2064 ? _T_2077 : _T_2091; // @[Mux.scala 31:69:@21906.4]
  assign _T_2093 = _T_2063 ? _T_2075 : _T_2092; // @[Mux.scala 31:69:@21907.4]
  assign _T_2094 = _T_2062 ? _T_2073 : _T_2093; // @[Mux.scala 31:69:@21908.4]
  assign _T_2095 = _T_2061 ? _T_2071 : _T_2094; // @[Mux.scala 31:69:@21909.4]
  assign _T_2103 = _T_1732 & _T_1550; // @[MemPrimitives.scala 110:228:@21918.4]
  assign _T_2109 = _T_1738 & _T_1556; // @[MemPrimitives.scala 110:228:@21922.4]
  assign _T_2115 = _T_1744 & _T_1562; // @[MemPrimitives.scala 110:228:@21926.4]
  assign _T_2121 = _T_1750 & _T_1568; // @[MemPrimitives.scala 110:228:@21930.4]
  assign _T_2127 = _T_1756 & _T_1574; // @[MemPrimitives.scala 110:228:@21934.4]
  assign _T_2133 = _T_1762 & _T_1580; // @[MemPrimitives.scala 110:228:@21938.4]
  assign _T_2139 = _T_1768 & _T_1586; // @[MemPrimitives.scala 110:228:@21942.4]
  assign _T_2145 = _T_1774 & _T_1592; // @[MemPrimitives.scala 110:228:@21946.4]
  assign _T_2151 = _T_1780 & _T_1598; // @[MemPrimitives.scala 110:228:@21950.4]
  assign _T_2153 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@21964.4]
  assign _T_2154 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@21965.4]
  assign _T_2155 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@21966.4]
  assign _T_2156 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@21967.4]
  assign _T_2157 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@21968.4]
  assign _T_2158 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@21969.4]
  assign _T_2159 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 126:35:@21970.4]
  assign _T_2160 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 126:35:@21971.4]
  assign _T_2161 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 126:35:@21972.4]
  assign _T_2163 = {_T_2153,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21974.4]
  assign _T_2165 = {_T_2154,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21976.4]
  assign _T_2167 = {_T_2155,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21978.4]
  assign _T_2169 = {_T_2156,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21980.4]
  assign _T_2171 = {_T_2157,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21982.4]
  assign _T_2173 = {_T_2158,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21984.4]
  assign _T_2175 = {_T_2159,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21986.4]
  assign _T_2177 = {_T_2160,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21988.4]
  assign _T_2179 = {_T_2161,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21990.4]
  assign _T_2180 = _T_2160 ? _T_2177 : _T_2179; // @[Mux.scala 31:69:@21991.4]
  assign _T_2181 = _T_2159 ? _T_2175 : _T_2180; // @[Mux.scala 31:69:@21992.4]
  assign _T_2182 = _T_2158 ? _T_2173 : _T_2181; // @[Mux.scala 31:69:@21993.4]
  assign _T_2183 = _T_2157 ? _T_2171 : _T_2182; // @[Mux.scala 31:69:@21994.4]
  assign _T_2184 = _T_2156 ? _T_2169 : _T_2183; // @[Mux.scala 31:69:@21995.4]
  assign _T_2185 = _T_2155 ? _T_2167 : _T_2184; // @[Mux.scala 31:69:@21996.4]
  assign _T_2186 = _T_2154 ? _T_2165 : _T_2185; // @[Mux.scala 31:69:@21997.4]
  assign _T_2187 = _T_2153 ? _T_2163 : _T_2186; // @[Mux.scala 31:69:@21998.4]
  assign _T_2195 = _T_1824 & _T_1642; // @[MemPrimitives.scala 110:228:@22007.4]
  assign _T_2201 = _T_1830 & _T_1648; // @[MemPrimitives.scala 110:228:@22011.4]
  assign _T_2207 = _T_1836 & _T_1654; // @[MemPrimitives.scala 110:228:@22015.4]
  assign _T_2213 = _T_1842 & _T_1660; // @[MemPrimitives.scala 110:228:@22019.4]
  assign _T_2219 = _T_1848 & _T_1666; // @[MemPrimitives.scala 110:228:@22023.4]
  assign _T_2225 = _T_1854 & _T_1672; // @[MemPrimitives.scala 110:228:@22027.4]
  assign _T_2231 = _T_1860 & _T_1678; // @[MemPrimitives.scala 110:228:@22031.4]
  assign _T_2237 = _T_1866 & _T_1684; // @[MemPrimitives.scala 110:228:@22035.4]
  assign _T_2243 = _T_1872 & _T_1690; // @[MemPrimitives.scala 110:228:@22039.4]
  assign _T_2245 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@22053.4]
  assign _T_2246 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@22054.4]
  assign _T_2247 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@22055.4]
  assign _T_2248 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@22056.4]
  assign _T_2249 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@22057.4]
  assign _T_2250 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@22058.4]
  assign _T_2251 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 126:35:@22059.4]
  assign _T_2252 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 126:35:@22060.4]
  assign _T_2253 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 126:35:@22061.4]
  assign _T_2255 = {_T_2245,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22063.4]
  assign _T_2257 = {_T_2246,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22065.4]
  assign _T_2259 = {_T_2247,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22067.4]
  assign _T_2261 = {_T_2248,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22069.4]
  assign _T_2263 = {_T_2249,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22071.4]
  assign _T_2265 = {_T_2250,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22073.4]
  assign _T_2267 = {_T_2251,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22075.4]
  assign _T_2269 = {_T_2252,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22077.4]
  assign _T_2271 = {_T_2253,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22079.4]
  assign _T_2272 = _T_2252 ? _T_2269 : _T_2271; // @[Mux.scala 31:69:@22080.4]
  assign _T_2273 = _T_2251 ? _T_2267 : _T_2272; // @[Mux.scala 31:69:@22081.4]
  assign _T_2274 = _T_2250 ? _T_2265 : _T_2273; // @[Mux.scala 31:69:@22082.4]
  assign _T_2275 = _T_2249 ? _T_2263 : _T_2274; // @[Mux.scala 31:69:@22083.4]
  assign _T_2276 = _T_2248 ? _T_2261 : _T_2275; // @[Mux.scala 31:69:@22084.4]
  assign _T_2277 = _T_2247 ? _T_2259 : _T_2276; // @[Mux.scala 31:69:@22085.4]
  assign _T_2278 = _T_2246 ? _T_2257 : _T_2277; // @[Mux.scala 31:69:@22086.4]
  assign _T_2279 = _T_2245 ? _T_2255 : _T_2278; // @[Mux.scala 31:69:@22087.4]
  assign _T_2284 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22094.4]
  assign _T_2287 = _T_2284 & _T_1182; // @[MemPrimitives.scala 110:228:@22096.4]
  assign _T_2290 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22098.4]
  assign _T_2293 = _T_2290 & _T_1188; // @[MemPrimitives.scala 110:228:@22100.4]
  assign _T_2296 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22102.4]
  assign _T_2299 = _T_2296 & _T_1194; // @[MemPrimitives.scala 110:228:@22104.4]
  assign _T_2302 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22106.4]
  assign _T_2305 = _T_2302 & _T_1200; // @[MemPrimitives.scala 110:228:@22108.4]
  assign _T_2308 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22110.4]
  assign _T_2311 = _T_2308 & _T_1206; // @[MemPrimitives.scala 110:228:@22112.4]
  assign _T_2314 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22114.4]
  assign _T_2317 = _T_2314 & _T_1212; // @[MemPrimitives.scala 110:228:@22116.4]
  assign _T_2320 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22118.4]
  assign _T_2323 = _T_2320 & _T_1218; // @[MemPrimitives.scala 110:228:@22120.4]
  assign _T_2326 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22122.4]
  assign _T_2329 = _T_2326 & _T_1224; // @[MemPrimitives.scala 110:228:@22124.4]
  assign _T_2332 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22126.4]
  assign _T_2335 = _T_2332 & _T_1230; // @[MemPrimitives.scala 110:228:@22128.4]
  assign _T_2337 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@22142.4]
  assign _T_2338 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@22143.4]
  assign _T_2339 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@22144.4]
  assign _T_2340 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@22145.4]
  assign _T_2341 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@22146.4]
  assign _T_2342 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@22147.4]
  assign _T_2343 = StickySelects_12_io_outs_6; // @[MemPrimitives.scala 126:35:@22148.4]
  assign _T_2344 = StickySelects_12_io_outs_7; // @[MemPrimitives.scala 126:35:@22149.4]
  assign _T_2345 = StickySelects_12_io_outs_8; // @[MemPrimitives.scala 126:35:@22150.4]
  assign _T_2347 = {_T_2337,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22152.4]
  assign _T_2349 = {_T_2338,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22154.4]
  assign _T_2351 = {_T_2339,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22156.4]
  assign _T_2353 = {_T_2340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22158.4]
  assign _T_2355 = {_T_2341,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22160.4]
  assign _T_2357 = {_T_2342,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22162.4]
  assign _T_2359 = {_T_2343,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22164.4]
  assign _T_2361 = {_T_2344,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22166.4]
  assign _T_2363 = {_T_2345,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22168.4]
  assign _T_2364 = _T_2344 ? _T_2361 : _T_2363; // @[Mux.scala 31:69:@22169.4]
  assign _T_2365 = _T_2343 ? _T_2359 : _T_2364; // @[Mux.scala 31:69:@22170.4]
  assign _T_2366 = _T_2342 ? _T_2357 : _T_2365; // @[Mux.scala 31:69:@22171.4]
  assign _T_2367 = _T_2341 ? _T_2355 : _T_2366; // @[Mux.scala 31:69:@22172.4]
  assign _T_2368 = _T_2340 ? _T_2353 : _T_2367; // @[Mux.scala 31:69:@22173.4]
  assign _T_2369 = _T_2339 ? _T_2351 : _T_2368; // @[Mux.scala 31:69:@22174.4]
  assign _T_2370 = _T_2338 ? _T_2349 : _T_2369; // @[Mux.scala 31:69:@22175.4]
  assign _T_2371 = _T_2337 ? _T_2347 : _T_2370; // @[Mux.scala 31:69:@22176.4]
  assign _T_2376 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22183.4]
  assign _T_2379 = _T_2376 & _T_1274; // @[MemPrimitives.scala 110:228:@22185.4]
  assign _T_2382 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22187.4]
  assign _T_2385 = _T_2382 & _T_1280; // @[MemPrimitives.scala 110:228:@22189.4]
  assign _T_2388 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22191.4]
  assign _T_2391 = _T_2388 & _T_1286; // @[MemPrimitives.scala 110:228:@22193.4]
  assign _T_2394 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22195.4]
  assign _T_2397 = _T_2394 & _T_1292; // @[MemPrimitives.scala 110:228:@22197.4]
  assign _T_2400 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22199.4]
  assign _T_2403 = _T_2400 & _T_1298; // @[MemPrimitives.scala 110:228:@22201.4]
  assign _T_2406 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22203.4]
  assign _T_2409 = _T_2406 & _T_1304; // @[MemPrimitives.scala 110:228:@22205.4]
  assign _T_2412 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22207.4]
  assign _T_2415 = _T_2412 & _T_1310; // @[MemPrimitives.scala 110:228:@22209.4]
  assign _T_2418 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22211.4]
  assign _T_2421 = _T_2418 & _T_1316; // @[MemPrimitives.scala 110:228:@22213.4]
  assign _T_2424 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22215.4]
  assign _T_2427 = _T_2424 & _T_1322; // @[MemPrimitives.scala 110:228:@22217.4]
  assign _T_2429 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@22231.4]
  assign _T_2430 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@22232.4]
  assign _T_2431 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@22233.4]
  assign _T_2432 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@22234.4]
  assign _T_2433 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@22235.4]
  assign _T_2434 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@22236.4]
  assign _T_2435 = StickySelects_13_io_outs_6; // @[MemPrimitives.scala 126:35:@22237.4]
  assign _T_2436 = StickySelects_13_io_outs_7; // @[MemPrimitives.scala 126:35:@22238.4]
  assign _T_2437 = StickySelects_13_io_outs_8; // @[MemPrimitives.scala 126:35:@22239.4]
  assign _T_2439 = {_T_2429,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22241.4]
  assign _T_2441 = {_T_2430,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22243.4]
  assign _T_2443 = {_T_2431,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22245.4]
  assign _T_2445 = {_T_2432,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22247.4]
  assign _T_2447 = {_T_2433,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22249.4]
  assign _T_2449 = {_T_2434,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22251.4]
  assign _T_2451 = {_T_2435,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22253.4]
  assign _T_2453 = {_T_2436,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22255.4]
  assign _T_2455 = {_T_2437,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22257.4]
  assign _T_2456 = _T_2436 ? _T_2453 : _T_2455; // @[Mux.scala 31:69:@22258.4]
  assign _T_2457 = _T_2435 ? _T_2451 : _T_2456; // @[Mux.scala 31:69:@22259.4]
  assign _T_2458 = _T_2434 ? _T_2449 : _T_2457; // @[Mux.scala 31:69:@22260.4]
  assign _T_2459 = _T_2433 ? _T_2447 : _T_2458; // @[Mux.scala 31:69:@22261.4]
  assign _T_2460 = _T_2432 ? _T_2445 : _T_2459; // @[Mux.scala 31:69:@22262.4]
  assign _T_2461 = _T_2431 ? _T_2443 : _T_2460; // @[Mux.scala 31:69:@22263.4]
  assign _T_2462 = _T_2430 ? _T_2441 : _T_2461; // @[Mux.scala 31:69:@22264.4]
  assign _T_2463 = _T_2429 ? _T_2439 : _T_2462; // @[Mux.scala 31:69:@22265.4]
  assign _T_2471 = _T_2284 & _T_1366; // @[MemPrimitives.scala 110:228:@22274.4]
  assign _T_2477 = _T_2290 & _T_1372; // @[MemPrimitives.scala 110:228:@22278.4]
  assign _T_2483 = _T_2296 & _T_1378; // @[MemPrimitives.scala 110:228:@22282.4]
  assign _T_2489 = _T_2302 & _T_1384; // @[MemPrimitives.scala 110:228:@22286.4]
  assign _T_2495 = _T_2308 & _T_1390; // @[MemPrimitives.scala 110:228:@22290.4]
  assign _T_2501 = _T_2314 & _T_1396; // @[MemPrimitives.scala 110:228:@22294.4]
  assign _T_2507 = _T_2320 & _T_1402; // @[MemPrimitives.scala 110:228:@22298.4]
  assign _T_2513 = _T_2326 & _T_1408; // @[MemPrimitives.scala 110:228:@22302.4]
  assign _T_2519 = _T_2332 & _T_1414; // @[MemPrimitives.scala 110:228:@22306.4]
  assign _T_2521 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@22320.4]
  assign _T_2522 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@22321.4]
  assign _T_2523 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@22322.4]
  assign _T_2524 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@22323.4]
  assign _T_2525 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@22324.4]
  assign _T_2526 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@22325.4]
  assign _T_2527 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 126:35:@22326.4]
  assign _T_2528 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 126:35:@22327.4]
  assign _T_2529 = StickySelects_14_io_outs_8; // @[MemPrimitives.scala 126:35:@22328.4]
  assign _T_2531 = {_T_2521,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22330.4]
  assign _T_2533 = {_T_2522,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22332.4]
  assign _T_2535 = {_T_2523,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22334.4]
  assign _T_2537 = {_T_2524,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22336.4]
  assign _T_2539 = {_T_2525,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22338.4]
  assign _T_2541 = {_T_2526,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22340.4]
  assign _T_2543 = {_T_2527,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22342.4]
  assign _T_2545 = {_T_2528,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22344.4]
  assign _T_2547 = {_T_2529,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22346.4]
  assign _T_2548 = _T_2528 ? _T_2545 : _T_2547; // @[Mux.scala 31:69:@22347.4]
  assign _T_2549 = _T_2527 ? _T_2543 : _T_2548; // @[Mux.scala 31:69:@22348.4]
  assign _T_2550 = _T_2526 ? _T_2541 : _T_2549; // @[Mux.scala 31:69:@22349.4]
  assign _T_2551 = _T_2525 ? _T_2539 : _T_2550; // @[Mux.scala 31:69:@22350.4]
  assign _T_2552 = _T_2524 ? _T_2537 : _T_2551; // @[Mux.scala 31:69:@22351.4]
  assign _T_2553 = _T_2523 ? _T_2535 : _T_2552; // @[Mux.scala 31:69:@22352.4]
  assign _T_2554 = _T_2522 ? _T_2533 : _T_2553; // @[Mux.scala 31:69:@22353.4]
  assign _T_2555 = _T_2521 ? _T_2531 : _T_2554; // @[Mux.scala 31:69:@22354.4]
  assign _T_2563 = _T_2376 & _T_1458; // @[MemPrimitives.scala 110:228:@22363.4]
  assign _T_2569 = _T_2382 & _T_1464; // @[MemPrimitives.scala 110:228:@22367.4]
  assign _T_2575 = _T_2388 & _T_1470; // @[MemPrimitives.scala 110:228:@22371.4]
  assign _T_2581 = _T_2394 & _T_1476; // @[MemPrimitives.scala 110:228:@22375.4]
  assign _T_2587 = _T_2400 & _T_1482; // @[MemPrimitives.scala 110:228:@22379.4]
  assign _T_2593 = _T_2406 & _T_1488; // @[MemPrimitives.scala 110:228:@22383.4]
  assign _T_2599 = _T_2412 & _T_1494; // @[MemPrimitives.scala 110:228:@22387.4]
  assign _T_2605 = _T_2418 & _T_1500; // @[MemPrimitives.scala 110:228:@22391.4]
  assign _T_2611 = _T_2424 & _T_1506; // @[MemPrimitives.scala 110:228:@22395.4]
  assign _T_2613 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@22409.4]
  assign _T_2614 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@22410.4]
  assign _T_2615 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@22411.4]
  assign _T_2616 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@22412.4]
  assign _T_2617 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@22413.4]
  assign _T_2618 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@22414.4]
  assign _T_2619 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 126:35:@22415.4]
  assign _T_2620 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 126:35:@22416.4]
  assign _T_2621 = StickySelects_15_io_outs_8; // @[MemPrimitives.scala 126:35:@22417.4]
  assign _T_2623 = {_T_2613,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22419.4]
  assign _T_2625 = {_T_2614,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22421.4]
  assign _T_2627 = {_T_2615,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22423.4]
  assign _T_2629 = {_T_2616,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22425.4]
  assign _T_2631 = {_T_2617,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22427.4]
  assign _T_2633 = {_T_2618,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22429.4]
  assign _T_2635 = {_T_2619,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22431.4]
  assign _T_2637 = {_T_2620,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22433.4]
  assign _T_2639 = {_T_2621,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22435.4]
  assign _T_2640 = _T_2620 ? _T_2637 : _T_2639; // @[Mux.scala 31:69:@22436.4]
  assign _T_2641 = _T_2619 ? _T_2635 : _T_2640; // @[Mux.scala 31:69:@22437.4]
  assign _T_2642 = _T_2618 ? _T_2633 : _T_2641; // @[Mux.scala 31:69:@22438.4]
  assign _T_2643 = _T_2617 ? _T_2631 : _T_2642; // @[Mux.scala 31:69:@22439.4]
  assign _T_2644 = _T_2616 ? _T_2629 : _T_2643; // @[Mux.scala 31:69:@22440.4]
  assign _T_2645 = _T_2615 ? _T_2627 : _T_2644; // @[Mux.scala 31:69:@22441.4]
  assign _T_2646 = _T_2614 ? _T_2625 : _T_2645; // @[Mux.scala 31:69:@22442.4]
  assign _T_2647 = _T_2613 ? _T_2623 : _T_2646; // @[Mux.scala 31:69:@22443.4]
  assign _T_2655 = _T_2284 & _T_1550; // @[MemPrimitives.scala 110:228:@22452.4]
  assign _T_2661 = _T_2290 & _T_1556; // @[MemPrimitives.scala 110:228:@22456.4]
  assign _T_2667 = _T_2296 & _T_1562; // @[MemPrimitives.scala 110:228:@22460.4]
  assign _T_2673 = _T_2302 & _T_1568; // @[MemPrimitives.scala 110:228:@22464.4]
  assign _T_2679 = _T_2308 & _T_1574; // @[MemPrimitives.scala 110:228:@22468.4]
  assign _T_2685 = _T_2314 & _T_1580; // @[MemPrimitives.scala 110:228:@22472.4]
  assign _T_2691 = _T_2320 & _T_1586; // @[MemPrimitives.scala 110:228:@22476.4]
  assign _T_2697 = _T_2326 & _T_1592; // @[MemPrimitives.scala 110:228:@22480.4]
  assign _T_2703 = _T_2332 & _T_1598; // @[MemPrimitives.scala 110:228:@22484.4]
  assign _T_2705 = StickySelects_16_io_outs_0; // @[MemPrimitives.scala 126:35:@22498.4]
  assign _T_2706 = StickySelects_16_io_outs_1; // @[MemPrimitives.scala 126:35:@22499.4]
  assign _T_2707 = StickySelects_16_io_outs_2; // @[MemPrimitives.scala 126:35:@22500.4]
  assign _T_2708 = StickySelects_16_io_outs_3; // @[MemPrimitives.scala 126:35:@22501.4]
  assign _T_2709 = StickySelects_16_io_outs_4; // @[MemPrimitives.scala 126:35:@22502.4]
  assign _T_2710 = StickySelects_16_io_outs_5; // @[MemPrimitives.scala 126:35:@22503.4]
  assign _T_2711 = StickySelects_16_io_outs_6; // @[MemPrimitives.scala 126:35:@22504.4]
  assign _T_2712 = StickySelects_16_io_outs_7; // @[MemPrimitives.scala 126:35:@22505.4]
  assign _T_2713 = StickySelects_16_io_outs_8; // @[MemPrimitives.scala 126:35:@22506.4]
  assign _T_2715 = {_T_2705,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22508.4]
  assign _T_2717 = {_T_2706,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22510.4]
  assign _T_2719 = {_T_2707,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22512.4]
  assign _T_2721 = {_T_2708,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22514.4]
  assign _T_2723 = {_T_2709,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22516.4]
  assign _T_2725 = {_T_2710,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22518.4]
  assign _T_2727 = {_T_2711,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22520.4]
  assign _T_2729 = {_T_2712,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22522.4]
  assign _T_2731 = {_T_2713,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22524.4]
  assign _T_2732 = _T_2712 ? _T_2729 : _T_2731; // @[Mux.scala 31:69:@22525.4]
  assign _T_2733 = _T_2711 ? _T_2727 : _T_2732; // @[Mux.scala 31:69:@22526.4]
  assign _T_2734 = _T_2710 ? _T_2725 : _T_2733; // @[Mux.scala 31:69:@22527.4]
  assign _T_2735 = _T_2709 ? _T_2723 : _T_2734; // @[Mux.scala 31:69:@22528.4]
  assign _T_2736 = _T_2708 ? _T_2721 : _T_2735; // @[Mux.scala 31:69:@22529.4]
  assign _T_2737 = _T_2707 ? _T_2719 : _T_2736; // @[Mux.scala 31:69:@22530.4]
  assign _T_2738 = _T_2706 ? _T_2717 : _T_2737; // @[Mux.scala 31:69:@22531.4]
  assign _T_2739 = _T_2705 ? _T_2715 : _T_2738; // @[Mux.scala 31:69:@22532.4]
  assign _T_2747 = _T_2376 & _T_1642; // @[MemPrimitives.scala 110:228:@22541.4]
  assign _T_2753 = _T_2382 & _T_1648; // @[MemPrimitives.scala 110:228:@22545.4]
  assign _T_2759 = _T_2388 & _T_1654; // @[MemPrimitives.scala 110:228:@22549.4]
  assign _T_2765 = _T_2394 & _T_1660; // @[MemPrimitives.scala 110:228:@22553.4]
  assign _T_2771 = _T_2400 & _T_1666; // @[MemPrimitives.scala 110:228:@22557.4]
  assign _T_2777 = _T_2406 & _T_1672; // @[MemPrimitives.scala 110:228:@22561.4]
  assign _T_2783 = _T_2412 & _T_1678; // @[MemPrimitives.scala 110:228:@22565.4]
  assign _T_2789 = _T_2418 & _T_1684; // @[MemPrimitives.scala 110:228:@22569.4]
  assign _T_2795 = _T_2424 & _T_1690; // @[MemPrimitives.scala 110:228:@22573.4]
  assign _T_2797 = StickySelects_17_io_outs_0; // @[MemPrimitives.scala 126:35:@22587.4]
  assign _T_2798 = StickySelects_17_io_outs_1; // @[MemPrimitives.scala 126:35:@22588.4]
  assign _T_2799 = StickySelects_17_io_outs_2; // @[MemPrimitives.scala 126:35:@22589.4]
  assign _T_2800 = StickySelects_17_io_outs_3; // @[MemPrimitives.scala 126:35:@22590.4]
  assign _T_2801 = StickySelects_17_io_outs_4; // @[MemPrimitives.scala 126:35:@22591.4]
  assign _T_2802 = StickySelects_17_io_outs_5; // @[MemPrimitives.scala 126:35:@22592.4]
  assign _T_2803 = StickySelects_17_io_outs_6; // @[MemPrimitives.scala 126:35:@22593.4]
  assign _T_2804 = StickySelects_17_io_outs_7; // @[MemPrimitives.scala 126:35:@22594.4]
  assign _T_2805 = StickySelects_17_io_outs_8; // @[MemPrimitives.scala 126:35:@22595.4]
  assign _T_2807 = {_T_2797,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22597.4]
  assign _T_2809 = {_T_2798,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22599.4]
  assign _T_2811 = {_T_2799,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22601.4]
  assign _T_2813 = {_T_2800,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22603.4]
  assign _T_2815 = {_T_2801,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22605.4]
  assign _T_2817 = {_T_2802,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22607.4]
  assign _T_2819 = {_T_2803,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22609.4]
  assign _T_2821 = {_T_2804,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22611.4]
  assign _T_2823 = {_T_2805,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22613.4]
  assign _T_2824 = _T_2804 ? _T_2821 : _T_2823; // @[Mux.scala 31:69:@22614.4]
  assign _T_2825 = _T_2803 ? _T_2819 : _T_2824; // @[Mux.scala 31:69:@22615.4]
  assign _T_2826 = _T_2802 ? _T_2817 : _T_2825; // @[Mux.scala 31:69:@22616.4]
  assign _T_2827 = _T_2801 ? _T_2815 : _T_2826; // @[Mux.scala 31:69:@22617.4]
  assign _T_2828 = _T_2800 ? _T_2813 : _T_2827; // @[Mux.scala 31:69:@22618.4]
  assign _T_2829 = _T_2799 ? _T_2811 : _T_2828; // @[Mux.scala 31:69:@22619.4]
  assign _T_2830 = _T_2798 ? _T_2809 : _T_2829; // @[Mux.scala 31:69:@22620.4]
  assign _T_2831 = _T_2797 ? _T_2807 : _T_2830; // @[Mux.scala 31:69:@22621.4]
  assign _T_2836 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22628.4]
  assign _T_2839 = _T_2836 & _T_1182; // @[MemPrimitives.scala 110:228:@22630.4]
  assign _T_2842 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22632.4]
  assign _T_2845 = _T_2842 & _T_1188; // @[MemPrimitives.scala 110:228:@22634.4]
  assign _T_2848 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22636.4]
  assign _T_2851 = _T_2848 & _T_1194; // @[MemPrimitives.scala 110:228:@22638.4]
  assign _T_2854 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22640.4]
  assign _T_2857 = _T_2854 & _T_1200; // @[MemPrimitives.scala 110:228:@22642.4]
  assign _T_2860 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22644.4]
  assign _T_2863 = _T_2860 & _T_1206; // @[MemPrimitives.scala 110:228:@22646.4]
  assign _T_2866 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22648.4]
  assign _T_2869 = _T_2866 & _T_1212; // @[MemPrimitives.scala 110:228:@22650.4]
  assign _T_2872 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22652.4]
  assign _T_2875 = _T_2872 & _T_1218; // @[MemPrimitives.scala 110:228:@22654.4]
  assign _T_2878 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22656.4]
  assign _T_2881 = _T_2878 & _T_1224; // @[MemPrimitives.scala 110:228:@22658.4]
  assign _T_2884 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22660.4]
  assign _T_2887 = _T_2884 & _T_1230; // @[MemPrimitives.scala 110:228:@22662.4]
  assign _T_2889 = StickySelects_18_io_outs_0; // @[MemPrimitives.scala 126:35:@22676.4]
  assign _T_2890 = StickySelects_18_io_outs_1; // @[MemPrimitives.scala 126:35:@22677.4]
  assign _T_2891 = StickySelects_18_io_outs_2; // @[MemPrimitives.scala 126:35:@22678.4]
  assign _T_2892 = StickySelects_18_io_outs_3; // @[MemPrimitives.scala 126:35:@22679.4]
  assign _T_2893 = StickySelects_18_io_outs_4; // @[MemPrimitives.scala 126:35:@22680.4]
  assign _T_2894 = StickySelects_18_io_outs_5; // @[MemPrimitives.scala 126:35:@22681.4]
  assign _T_2895 = StickySelects_18_io_outs_6; // @[MemPrimitives.scala 126:35:@22682.4]
  assign _T_2896 = StickySelects_18_io_outs_7; // @[MemPrimitives.scala 126:35:@22683.4]
  assign _T_2897 = StickySelects_18_io_outs_8; // @[MemPrimitives.scala 126:35:@22684.4]
  assign _T_2899 = {_T_2889,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22686.4]
  assign _T_2901 = {_T_2890,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22688.4]
  assign _T_2903 = {_T_2891,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22690.4]
  assign _T_2905 = {_T_2892,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22692.4]
  assign _T_2907 = {_T_2893,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22694.4]
  assign _T_2909 = {_T_2894,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22696.4]
  assign _T_2911 = {_T_2895,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22698.4]
  assign _T_2913 = {_T_2896,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22700.4]
  assign _T_2915 = {_T_2897,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22702.4]
  assign _T_2916 = _T_2896 ? _T_2913 : _T_2915; // @[Mux.scala 31:69:@22703.4]
  assign _T_2917 = _T_2895 ? _T_2911 : _T_2916; // @[Mux.scala 31:69:@22704.4]
  assign _T_2918 = _T_2894 ? _T_2909 : _T_2917; // @[Mux.scala 31:69:@22705.4]
  assign _T_2919 = _T_2893 ? _T_2907 : _T_2918; // @[Mux.scala 31:69:@22706.4]
  assign _T_2920 = _T_2892 ? _T_2905 : _T_2919; // @[Mux.scala 31:69:@22707.4]
  assign _T_2921 = _T_2891 ? _T_2903 : _T_2920; // @[Mux.scala 31:69:@22708.4]
  assign _T_2922 = _T_2890 ? _T_2901 : _T_2921; // @[Mux.scala 31:69:@22709.4]
  assign _T_2923 = _T_2889 ? _T_2899 : _T_2922; // @[Mux.scala 31:69:@22710.4]
  assign _T_2928 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22717.4]
  assign _T_2931 = _T_2928 & _T_1274; // @[MemPrimitives.scala 110:228:@22719.4]
  assign _T_2934 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22721.4]
  assign _T_2937 = _T_2934 & _T_1280; // @[MemPrimitives.scala 110:228:@22723.4]
  assign _T_2940 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22725.4]
  assign _T_2943 = _T_2940 & _T_1286; // @[MemPrimitives.scala 110:228:@22727.4]
  assign _T_2946 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22729.4]
  assign _T_2949 = _T_2946 & _T_1292; // @[MemPrimitives.scala 110:228:@22731.4]
  assign _T_2952 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22733.4]
  assign _T_2955 = _T_2952 & _T_1298; // @[MemPrimitives.scala 110:228:@22735.4]
  assign _T_2958 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22737.4]
  assign _T_2961 = _T_2958 & _T_1304; // @[MemPrimitives.scala 110:228:@22739.4]
  assign _T_2964 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22741.4]
  assign _T_2967 = _T_2964 & _T_1310; // @[MemPrimitives.scala 110:228:@22743.4]
  assign _T_2970 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22745.4]
  assign _T_2973 = _T_2970 & _T_1316; // @[MemPrimitives.scala 110:228:@22747.4]
  assign _T_2976 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22749.4]
  assign _T_2979 = _T_2976 & _T_1322; // @[MemPrimitives.scala 110:228:@22751.4]
  assign _T_2981 = StickySelects_19_io_outs_0; // @[MemPrimitives.scala 126:35:@22765.4]
  assign _T_2982 = StickySelects_19_io_outs_1; // @[MemPrimitives.scala 126:35:@22766.4]
  assign _T_2983 = StickySelects_19_io_outs_2; // @[MemPrimitives.scala 126:35:@22767.4]
  assign _T_2984 = StickySelects_19_io_outs_3; // @[MemPrimitives.scala 126:35:@22768.4]
  assign _T_2985 = StickySelects_19_io_outs_4; // @[MemPrimitives.scala 126:35:@22769.4]
  assign _T_2986 = StickySelects_19_io_outs_5; // @[MemPrimitives.scala 126:35:@22770.4]
  assign _T_2987 = StickySelects_19_io_outs_6; // @[MemPrimitives.scala 126:35:@22771.4]
  assign _T_2988 = StickySelects_19_io_outs_7; // @[MemPrimitives.scala 126:35:@22772.4]
  assign _T_2989 = StickySelects_19_io_outs_8; // @[MemPrimitives.scala 126:35:@22773.4]
  assign _T_2991 = {_T_2981,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22775.4]
  assign _T_2993 = {_T_2982,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22777.4]
  assign _T_2995 = {_T_2983,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22779.4]
  assign _T_2997 = {_T_2984,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22781.4]
  assign _T_2999 = {_T_2985,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22783.4]
  assign _T_3001 = {_T_2986,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22785.4]
  assign _T_3003 = {_T_2987,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22787.4]
  assign _T_3005 = {_T_2988,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22789.4]
  assign _T_3007 = {_T_2989,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22791.4]
  assign _T_3008 = _T_2988 ? _T_3005 : _T_3007; // @[Mux.scala 31:69:@22792.4]
  assign _T_3009 = _T_2987 ? _T_3003 : _T_3008; // @[Mux.scala 31:69:@22793.4]
  assign _T_3010 = _T_2986 ? _T_3001 : _T_3009; // @[Mux.scala 31:69:@22794.4]
  assign _T_3011 = _T_2985 ? _T_2999 : _T_3010; // @[Mux.scala 31:69:@22795.4]
  assign _T_3012 = _T_2984 ? _T_2997 : _T_3011; // @[Mux.scala 31:69:@22796.4]
  assign _T_3013 = _T_2983 ? _T_2995 : _T_3012; // @[Mux.scala 31:69:@22797.4]
  assign _T_3014 = _T_2982 ? _T_2993 : _T_3013; // @[Mux.scala 31:69:@22798.4]
  assign _T_3015 = _T_2981 ? _T_2991 : _T_3014; // @[Mux.scala 31:69:@22799.4]
  assign _T_3023 = _T_2836 & _T_1366; // @[MemPrimitives.scala 110:228:@22808.4]
  assign _T_3029 = _T_2842 & _T_1372; // @[MemPrimitives.scala 110:228:@22812.4]
  assign _T_3035 = _T_2848 & _T_1378; // @[MemPrimitives.scala 110:228:@22816.4]
  assign _T_3041 = _T_2854 & _T_1384; // @[MemPrimitives.scala 110:228:@22820.4]
  assign _T_3047 = _T_2860 & _T_1390; // @[MemPrimitives.scala 110:228:@22824.4]
  assign _T_3053 = _T_2866 & _T_1396; // @[MemPrimitives.scala 110:228:@22828.4]
  assign _T_3059 = _T_2872 & _T_1402; // @[MemPrimitives.scala 110:228:@22832.4]
  assign _T_3065 = _T_2878 & _T_1408; // @[MemPrimitives.scala 110:228:@22836.4]
  assign _T_3071 = _T_2884 & _T_1414; // @[MemPrimitives.scala 110:228:@22840.4]
  assign _T_3073 = StickySelects_20_io_outs_0; // @[MemPrimitives.scala 126:35:@22854.4]
  assign _T_3074 = StickySelects_20_io_outs_1; // @[MemPrimitives.scala 126:35:@22855.4]
  assign _T_3075 = StickySelects_20_io_outs_2; // @[MemPrimitives.scala 126:35:@22856.4]
  assign _T_3076 = StickySelects_20_io_outs_3; // @[MemPrimitives.scala 126:35:@22857.4]
  assign _T_3077 = StickySelects_20_io_outs_4; // @[MemPrimitives.scala 126:35:@22858.4]
  assign _T_3078 = StickySelects_20_io_outs_5; // @[MemPrimitives.scala 126:35:@22859.4]
  assign _T_3079 = StickySelects_20_io_outs_6; // @[MemPrimitives.scala 126:35:@22860.4]
  assign _T_3080 = StickySelects_20_io_outs_7; // @[MemPrimitives.scala 126:35:@22861.4]
  assign _T_3081 = StickySelects_20_io_outs_8; // @[MemPrimitives.scala 126:35:@22862.4]
  assign _T_3083 = {_T_3073,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22864.4]
  assign _T_3085 = {_T_3074,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22866.4]
  assign _T_3087 = {_T_3075,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22868.4]
  assign _T_3089 = {_T_3076,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22870.4]
  assign _T_3091 = {_T_3077,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22872.4]
  assign _T_3093 = {_T_3078,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22874.4]
  assign _T_3095 = {_T_3079,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22876.4]
  assign _T_3097 = {_T_3080,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22878.4]
  assign _T_3099 = {_T_3081,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22880.4]
  assign _T_3100 = _T_3080 ? _T_3097 : _T_3099; // @[Mux.scala 31:69:@22881.4]
  assign _T_3101 = _T_3079 ? _T_3095 : _T_3100; // @[Mux.scala 31:69:@22882.4]
  assign _T_3102 = _T_3078 ? _T_3093 : _T_3101; // @[Mux.scala 31:69:@22883.4]
  assign _T_3103 = _T_3077 ? _T_3091 : _T_3102; // @[Mux.scala 31:69:@22884.4]
  assign _T_3104 = _T_3076 ? _T_3089 : _T_3103; // @[Mux.scala 31:69:@22885.4]
  assign _T_3105 = _T_3075 ? _T_3087 : _T_3104; // @[Mux.scala 31:69:@22886.4]
  assign _T_3106 = _T_3074 ? _T_3085 : _T_3105; // @[Mux.scala 31:69:@22887.4]
  assign _T_3107 = _T_3073 ? _T_3083 : _T_3106; // @[Mux.scala 31:69:@22888.4]
  assign _T_3115 = _T_2928 & _T_1458; // @[MemPrimitives.scala 110:228:@22897.4]
  assign _T_3121 = _T_2934 & _T_1464; // @[MemPrimitives.scala 110:228:@22901.4]
  assign _T_3127 = _T_2940 & _T_1470; // @[MemPrimitives.scala 110:228:@22905.4]
  assign _T_3133 = _T_2946 & _T_1476; // @[MemPrimitives.scala 110:228:@22909.4]
  assign _T_3139 = _T_2952 & _T_1482; // @[MemPrimitives.scala 110:228:@22913.4]
  assign _T_3145 = _T_2958 & _T_1488; // @[MemPrimitives.scala 110:228:@22917.4]
  assign _T_3151 = _T_2964 & _T_1494; // @[MemPrimitives.scala 110:228:@22921.4]
  assign _T_3157 = _T_2970 & _T_1500; // @[MemPrimitives.scala 110:228:@22925.4]
  assign _T_3163 = _T_2976 & _T_1506; // @[MemPrimitives.scala 110:228:@22929.4]
  assign _T_3165 = StickySelects_21_io_outs_0; // @[MemPrimitives.scala 126:35:@22943.4]
  assign _T_3166 = StickySelects_21_io_outs_1; // @[MemPrimitives.scala 126:35:@22944.4]
  assign _T_3167 = StickySelects_21_io_outs_2; // @[MemPrimitives.scala 126:35:@22945.4]
  assign _T_3168 = StickySelects_21_io_outs_3; // @[MemPrimitives.scala 126:35:@22946.4]
  assign _T_3169 = StickySelects_21_io_outs_4; // @[MemPrimitives.scala 126:35:@22947.4]
  assign _T_3170 = StickySelects_21_io_outs_5; // @[MemPrimitives.scala 126:35:@22948.4]
  assign _T_3171 = StickySelects_21_io_outs_6; // @[MemPrimitives.scala 126:35:@22949.4]
  assign _T_3172 = StickySelects_21_io_outs_7; // @[MemPrimitives.scala 126:35:@22950.4]
  assign _T_3173 = StickySelects_21_io_outs_8; // @[MemPrimitives.scala 126:35:@22951.4]
  assign _T_3175 = {_T_3165,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22953.4]
  assign _T_3177 = {_T_3166,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22955.4]
  assign _T_3179 = {_T_3167,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22957.4]
  assign _T_3181 = {_T_3168,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22959.4]
  assign _T_3183 = {_T_3169,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22961.4]
  assign _T_3185 = {_T_3170,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22963.4]
  assign _T_3187 = {_T_3171,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22965.4]
  assign _T_3189 = {_T_3172,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22967.4]
  assign _T_3191 = {_T_3173,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22969.4]
  assign _T_3192 = _T_3172 ? _T_3189 : _T_3191; // @[Mux.scala 31:69:@22970.4]
  assign _T_3193 = _T_3171 ? _T_3187 : _T_3192; // @[Mux.scala 31:69:@22971.4]
  assign _T_3194 = _T_3170 ? _T_3185 : _T_3193; // @[Mux.scala 31:69:@22972.4]
  assign _T_3195 = _T_3169 ? _T_3183 : _T_3194; // @[Mux.scala 31:69:@22973.4]
  assign _T_3196 = _T_3168 ? _T_3181 : _T_3195; // @[Mux.scala 31:69:@22974.4]
  assign _T_3197 = _T_3167 ? _T_3179 : _T_3196; // @[Mux.scala 31:69:@22975.4]
  assign _T_3198 = _T_3166 ? _T_3177 : _T_3197; // @[Mux.scala 31:69:@22976.4]
  assign _T_3199 = _T_3165 ? _T_3175 : _T_3198; // @[Mux.scala 31:69:@22977.4]
  assign _T_3207 = _T_2836 & _T_1550; // @[MemPrimitives.scala 110:228:@22986.4]
  assign _T_3213 = _T_2842 & _T_1556; // @[MemPrimitives.scala 110:228:@22990.4]
  assign _T_3219 = _T_2848 & _T_1562; // @[MemPrimitives.scala 110:228:@22994.4]
  assign _T_3225 = _T_2854 & _T_1568; // @[MemPrimitives.scala 110:228:@22998.4]
  assign _T_3231 = _T_2860 & _T_1574; // @[MemPrimitives.scala 110:228:@23002.4]
  assign _T_3237 = _T_2866 & _T_1580; // @[MemPrimitives.scala 110:228:@23006.4]
  assign _T_3243 = _T_2872 & _T_1586; // @[MemPrimitives.scala 110:228:@23010.4]
  assign _T_3249 = _T_2878 & _T_1592; // @[MemPrimitives.scala 110:228:@23014.4]
  assign _T_3255 = _T_2884 & _T_1598; // @[MemPrimitives.scala 110:228:@23018.4]
  assign _T_3257 = StickySelects_22_io_outs_0; // @[MemPrimitives.scala 126:35:@23032.4]
  assign _T_3258 = StickySelects_22_io_outs_1; // @[MemPrimitives.scala 126:35:@23033.4]
  assign _T_3259 = StickySelects_22_io_outs_2; // @[MemPrimitives.scala 126:35:@23034.4]
  assign _T_3260 = StickySelects_22_io_outs_3; // @[MemPrimitives.scala 126:35:@23035.4]
  assign _T_3261 = StickySelects_22_io_outs_4; // @[MemPrimitives.scala 126:35:@23036.4]
  assign _T_3262 = StickySelects_22_io_outs_5; // @[MemPrimitives.scala 126:35:@23037.4]
  assign _T_3263 = StickySelects_22_io_outs_6; // @[MemPrimitives.scala 126:35:@23038.4]
  assign _T_3264 = StickySelects_22_io_outs_7; // @[MemPrimitives.scala 126:35:@23039.4]
  assign _T_3265 = StickySelects_22_io_outs_8; // @[MemPrimitives.scala 126:35:@23040.4]
  assign _T_3267 = {_T_3257,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@23042.4]
  assign _T_3269 = {_T_3258,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@23044.4]
  assign _T_3271 = {_T_3259,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@23046.4]
  assign _T_3273 = {_T_3260,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@23048.4]
  assign _T_3275 = {_T_3261,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@23050.4]
  assign _T_3277 = {_T_3262,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@23052.4]
  assign _T_3279 = {_T_3263,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@23054.4]
  assign _T_3281 = {_T_3264,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@23056.4]
  assign _T_3283 = {_T_3265,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@23058.4]
  assign _T_3284 = _T_3264 ? _T_3281 : _T_3283; // @[Mux.scala 31:69:@23059.4]
  assign _T_3285 = _T_3263 ? _T_3279 : _T_3284; // @[Mux.scala 31:69:@23060.4]
  assign _T_3286 = _T_3262 ? _T_3277 : _T_3285; // @[Mux.scala 31:69:@23061.4]
  assign _T_3287 = _T_3261 ? _T_3275 : _T_3286; // @[Mux.scala 31:69:@23062.4]
  assign _T_3288 = _T_3260 ? _T_3273 : _T_3287; // @[Mux.scala 31:69:@23063.4]
  assign _T_3289 = _T_3259 ? _T_3271 : _T_3288; // @[Mux.scala 31:69:@23064.4]
  assign _T_3290 = _T_3258 ? _T_3269 : _T_3289; // @[Mux.scala 31:69:@23065.4]
  assign _T_3291 = _T_3257 ? _T_3267 : _T_3290; // @[Mux.scala 31:69:@23066.4]
  assign _T_3299 = _T_2928 & _T_1642; // @[MemPrimitives.scala 110:228:@23075.4]
  assign _T_3305 = _T_2934 & _T_1648; // @[MemPrimitives.scala 110:228:@23079.4]
  assign _T_3311 = _T_2940 & _T_1654; // @[MemPrimitives.scala 110:228:@23083.4]
  assign _T_3317 = _T_2946 & _T_1660; // @[MemPrimitives.scala 110:228:@23087.4]
  assign _T_3323 = _T_2952 & _T_1666; // @[MemPrimitives.scala 110:228:@23091.4]
  assign _T_3329 = _T_2958 & _T_1672; // @[MemPrimitives.scala 110:228:@23095.4]
  assign _T_3335 = _T_2964 & _T_1678; // @[MemPrimitives.scala 110:228:@23099.4]
  assign _T_3341 = _T_2970 & _T_1684; // @[MemPrimitives.scala 110:228:@23103.4]
  assign _T_3347 = _T_2976 & _T_1690; // @[MemPrimitives.scala 110:228:@23107.4]
  assign _T_3349 = StickySelects_23_io_outs_0; // @[MemPrimitives.scala 126:35:@23121.4]
  assign _T_3350 = StickySelects_23_io_outs_1; // @[MemPrimitives.scala 126:35:@23122.4]
  assign _T_3351 = StickySelects_23_io_outs_2; // @[MemPrimitives.scala 126:35:@23123.4]
  assign _T_3352 = StickySelects_23_io_outs_3; // @[MemPrimitives.scala 126:35:@23124.4]
  assign _T_3353 = StickySelects_23_io_outs_4; // @[MemPrimitives.scala 126:35:@23125.4]
  assign _T_3354 = StickySelects_23_io_outs_5; // @[MemPrimitives.scala 126:35:@23126.4]
  assign _T_3355 = StickySelects_23_io_outs_6; // @[MemPrimitives.scala 126:35:@23127.4]
  assign _T_3356 = StickySelects_23_io_outs_7; // @[MemPrimitives.scala 126:35:@23128.4]
  assign _T_3357 = StickySelects_23_io_outs_8; // @[MemPrimitives.scala 126:35:@23129.4]
  assign _T_3359 = {_T_3349,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@23131.4]
  assign _T_3361 = {_T_3350,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@23133.4]
  assign _T_3363 = {_T_3351,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@23135.4]
  assign _T_3365 = {_T_3352,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@23137.4]
  assign _T_3367 = {_T_3353,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@23139.4]
  assign _T_3369 = {_T_3354,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@23141.4]
  assign _T_3371 = {_T_3355,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@23143.4]
  assign _T_3373 = {_T_3356,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@23145.4]
  assign _T_3375 = {_T_3357,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@23147.4]
  assign _T_3376 = _T_3356 ? _T_3373 : _T_3375; // @[Mux.scala 31:69:@23148.4]
  assign _T_3377 = _T_3355 ? _T_3371 : _T_3376; // @[Mux.scala 31:69:@23149.4]
  assign _T_3378 = _T_3354 ? _T_3369 : _T_3377; // @[Mux.scala 31:69:@23150.4]
  assign _T_3379 = _T_3353 ? _T_3367 : _T_3378; // @[Mux.scala 31:69:@23151.4]
  assign _T_3380 = _T_3352 ? _T_3365 : _T_3379; // @[Mux.scala 31:69:@23152.4]
  assign _T_3381 = _T_3351 ? _T_3363 : _T_3380; // @[Mux.scala 31:69:@23153.4]
  assign _T_3382 = _T_3350 ? _T_3361 : _T_3381; // @[Mux.scala 31:69:@23154.4]
  assign _T_3383 = _T_3349 ? _T_3359 : _T_3382; // @[Mux.scala 31:69:@23155.4]
  assign _T_3479 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@23284.4 package.scala 96:25:@23285.4]
  assign _T_3483 = _T_3479 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23294.4]
  assign _T_3476 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@23276.4 package.scala 96:25:@23277.4]
  assign _T_3484 = _T_3476 ? Mem1D_18_io_output : _T_3483; // @[Mux.scala 31:69:@23295.4]
  assign _T_3473 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@23268.4 package.scala 96:25:@23269.4]
  assign _T_3485 = _T_3473 ? Mem1D_16_io_output : _T_3484; // @[Mux.scala 31:69:@23296.4]
  assign _T_3470 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@23260.4 package.scala 96:25:@23261.4]
  assign _T_3486 = _T_3470 ? Mem1D_14_io_output : _T_3485; // @[Mux.scala 31:69:@23297.4]
  assign _T_3467 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@23252.4 package.scala 96:25:@23253.4]
  assign _T_3487 = _T_3467 ? Mem1D_12_io_output : _T_3486; // @[Mux.scala 31:69:@23298.4]
  assign _T_3464 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@23244.4 package.scala 96:25:@23245.4]
  assign _T_3488 = _T_3464 ? Mem1D_10_io_output : _T_3487; // @[Mux.scala 31:69:@23299.4]
  assign _T_3461 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@23236.4 package.scala 96:25:@23237.4]
  assign _T_3489 = _T_3461 ? Mem1D_8_io_output : _T_3488; // @[Mux.scala 31:69:@23300.4]
  assign _T_3458 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@23228.4 package.scala 96:25:@23229.4]
  assign _T_3490 = _T_3458 ? Mem1D_6_io_output : _T_3489; // @[Mux.scala 31:69:@23301.4]
  assign _T_3455 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@23220.4 package.scala 96:25:@23221.4]
  assign _T_3491 = _T_3455 ? Mem1D_4_io_output : _T_3490; // @[Mux.scala 31:69:@23302.4]
  assign _T_3452 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@23212.4 package.scala 96:25:@23213.4]
  assign _T_3492 = _T_3452 ? Mem1D_2_io_output : _T_3491; // @[Mux.scala 31:69:@23303.4]
  assign _T_3449 = RetimeWrapper_io_out; // @[package.scala 96:25:@23204.4 package.scala 96:25:@23205.4]
  assign _T_3586 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@23428.4 package.scala 96:25:@23429.4]
  assign _T_3590 = _T_3586 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23438.4]
  assign _T_3583 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@23420.4 package.scala 96:25:@23421.4]
  assign _T_3591 = _T_3583 ? Mem1D_18_io_output : _T_3590; // @[Mux.scala 31:69:@23439.4]
  assign _T_3580 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@23412.4 package.scala 96:25:@23413.4]
  assign _T_3592 = _T_3580 ? Mem1D_16_io_output : _T_3591; // @[Mux.scala 31:69:@23440.4]
  assign _T_3577 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@23404.4 package.scala 96:25:@23405.4]
  assign _T_3593 = _T_3577 ? Mem1D_14_io_output : _T_3592; // @[Mux.scala 31:69:@23441.4]
  assign _T_3574 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@23396.4 package.scala 96:25:@23397.4]
  assign _T_3594 = _T_3574 ? Mem1D_12_io_output : _T_3593; // @[Mux.scala 31:69:@23442.4]
  assign _T_3571 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@23388.4 package.scala 96:25:@23389.4]
  assign _T_3595 = _T_3571 ? Mem1D_10_io_output : _T_3594; // @[Mux.scala 31:69:@23443.4]
  assign _T_3568 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@23380.4 package.scala 96:25:@23381.4]
  assign _T_3596 = _T_3568 ? Mem1D_8_io_output : _T_3595; // @[Mux.scala 31:69:@23444.4]
  assign _T_3565 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@23372.4 package.scala 96:25:@23373.4]
  assign _T_3597 = _T_3565 ? Mem1D_6_io_output : _T_3596; // @[Mux.scala 31:69:@23445.4]
  assign _T_3562 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@23364.4 package.scala 96:25:@23365.4]
  assign _T_3598 = _T_3562 ? Mem1D_4_io_output : _T_3597; // @[Mux.scala 31:69:@23446.4]
  assign _T_3559 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@23356.4 package.scala 96:25:@23357.4]
  assign _T_3599 = _T_3559 ? Mem1D_2_io_output : _T_3598; // @[Mux.scala 31:69:@23447.4]
  assign _T_3556 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@23348.4 package.scala 96:25:@23349.4]
  assign _T_3693 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@23572.4 package.scala 96:25:@23573.4]
  assign _T_3697 = _T_3693 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23582.4]
  assign _T_3690 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@23564.4 package.scala 96:25:@23565.4]
  assign _T_3698 = _T_3690 ? Mem1D_19_io_output : _T_3697; // @[Mux.scala 31:69:@23583.4]
  assign _T_3687 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@23556.4 package.scala 96:25:@23557.4]
  assign _T_3699 = _T_3687 ? Mem1D_17_io_output : _T_3698; // @[Mux.scala 31:69:@23584.4]
  assign _T_3684 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@23548.4 package.scala 96:25:@23549.4]
  assign _T_3700 = _T_3684 ? Mem1D_15_io_output : _T_3699; // @[Mux.scala 31:69:@23585.4]
  assign _T_3681 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@23540.4 package.scala 96:25:@23541.4]
  assign _T_3701 = _T_3681 ? Mem1D_13_io_output : _T_3700; // @[Mux.scala 31:69:@23586.4]
  assign _T_3678 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@23532.4 package.scala 96:25:@23533.4]
  assign _T_3702 = _T_3678 ? Mem1D_11_io_output : _T_3701; // @[Mux.scala 31:69:@23587.4]
  assign _T_3675 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@23524.4 package.scala 96:25:@23525.4]
  assign _T_3703 = _T_3675 ? Mem1D_9_io_output : _T_3702; // @[Mux.scala 31:69:@23588.4]
  assign _T_3672 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@23516.4 package.scala 96:25:@23517.4]
  assign _T_3704 = _T_3672 ? Mem1D_7_io_output : _T_3703; // @[Mux.scala 31:69:@23589.4]
  assign _T_3669 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@23508.4 package.scala 96:25:@23509.4]
  assign _T_3705 = _T_3669 ? Mem1D_5_io_output : _T_3704; // @[Mux.scala 31:69:@23590.4]
  assign _T_3666 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@23500.4 package.scala 96:25:@23501.4]
  assign _T_3706 = _T_3666 ? Mem1D_3_io_output : _T_3705; // @[Mux.scala 31:69:@23591.4]
  assign _T_3663 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@23492.4 package.scala 96:25:@23493.4]
  assign _T_3800 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@23716.4 package.scala 96:25:@23717.4]
  assign _T_3804 = _T_3800 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23726.4]
  assign _T_3797 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@23708.4 package.scala 96:25:@23709.4]
  assign _T_3805 = _T_3797 ? Mem1D_19_io_output : _T_3804; // @[Mux.scala 31:69:@23727.4]
  assign _T_3794 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@23700.4 package.scala 96:25:@23701.4]
  assign _T_3806 = _T_3794 ? Mem1D_17_io_output : _T_3805; // @[Mux.scala 31:69:@23728.4]
  assign _T_3791 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@23692.4 package.scala 96:25:@23693.4]
  assign _T_3807 = _T_3791 ? Mem1D_15_io_output : _T_3806; // @[Mux.scala 31:69:@23729.4]
  assign _T_3788 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@23684.4 package.scala 96:25:@23685.4]
  assign _T_3808 = _T_3788 ? Mem1D_13_io_output : _T_3807; // @[Mux.scala 31:69:@23730.4]
  assign _T_3785 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@23676.4 package.scala 96:25:@23677.4]
  assign _T_3809 = _T_3785 ? Mem1D_11_io_output : _T_3808; // @[Mux.scala 31:69:@23731.4]
  assign _T_3782 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@23668.4 package.scala 96:25:@23669.4]
  assign _T_3810 = _T_3782 ? Mem1D_9_io_output : _T_3809; // @[Mux.scala 31:69:@23732.4]
  assign _T_3779 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@23660.4 package.scala 96:25:@23661.4]
  assign _T_3811 = _T_3779 ? Mem1D_7_io_output : _T_3810; // @[Mux.scala 31:69:@23733.4]
  assign _T_3776 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@23652.4 package.scala 96:25:@23653.4]
  assign _T_3812 = _T_3776 ? Mem1D_5_io_output : _T_3811; // @[Mux.scala 31:69:@23734.4]
  assign _T_3773 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@23644.4 package.scala 96:25:@23645.4]
  assign _T_3813 = _T_3773 ? Mem1D_3_io_output : _T_3812; // @[Mux.scala 31:69:@23735.4]
  assign _T_3770 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@23636.4 package.scala 96:25:@23637.4]
  assign _T_3907 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@23860.4 package.scala 96:25:@23861.4]
  assign _T_3911 = _T_3907 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23870.4]
  assign _T_3904 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@23852.4 package.scala 96:25:@23853.4]
  assign _T_3912 = _T_3904 ? Mem1D_19_io_output : _T_3911; // @[Mux.scala 31:69:@23871.4]
  assign _T_3901 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@23844.4 package.scala 96:25:@23845.4]
  assign _T_3913 = _T_3901 ? Mem1D_17_io_output : _T_3912; // @[Mux.scala 31:69:@23872.4]
  assign _T_3898 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@23836.4 package.scala 96:25:@23837.4]
  assign _T_3914 = _T_3898 ? Mem1D_15_io_output : _T_3913; // @[Mux.scala 31:69:@23873.4]
  assign _T_3895 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@23828.4 package.scala 96:25:@23829.4]
  assign _T_3915 = _T_3895 ? Mem1D_13_io_output : _T_3914; // @[Mux.scala 31:69:@23874.4]
  assign _T_3892 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@23820.4 package.scala 96:25:@23821.4]
  assign _T_3916 = _T_3892 ? Mem1D_11_io_output : _T_3915; // @[Mux.scala 31:69:@23875.4]
  assign _T_3889 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@23812.4 package.scala 96:25:@23813.4]
  assign _T_3917 = _T_3889 ? Mem1D_9_io_output : _T_3916; // @[Mux.scala 31:69:@23876.4]
  assign _T_3886 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@23804.4 package.scala 96:25:@23805.4]
  assign _T_3918 = _T_3886 ? Mem1D_7_io_output : _T_3917; // @[Mux.scala 31:69:@23877.4]
  assign _T_3883 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@23796.4 package.scala 96:25:@23797.4]
  assign _T_3919 = _T_3883 ? Mem1D_5_io_output : _T_3918; // @[Mux.scala 31:69:@23878.4]
  assign _T_3880 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@23788.4 package.scala 96:25:@23789.4]
  assign _T_3920 = _T_3880 ? Mem1D_3_io_output : _T_3919; // @[Mux.scala 31:69:@23879.4]
  assign _T_3877 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@23780.4 package.scala 96:25:@23781.4]
  assign _T_4014 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@24004.4 package.scala 96:25:@24005.4]
  assign _T_4018 = _T_4014 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24014.4]
  assign _T_4011 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@23996.4 package.scala 96:25:@23997.4]
  assign _T_4019 = _T_4011 ? Mem1D_18_io_output : _T_4018; // @[Mux.scala 31:69:@24015.4]
  assign _T_4008 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@23988.4 package.scala 96:25:@23989.4]
  assign _T_4020 = _T_4008 ? Mem1D_16_io_output : _T_4019; // @[Mux.scala 31:69:@24016.4]
  assign _T_4005 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@23980.4 package.scala 96:25:@23981.4]
  assign _T_4021 = _T_4005 ? Mem1D_14_io_output : _T_4020; // @[Mux.scala 31:69:@24017.4]
  assign _T_4002 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@23972.4 package.scala 96:25:@23973.4]
  assign _T_4022 = _T_4002 ? Mem1D_12_io_output : _T_4021; // @[Mux.scala 31:69:@24018.4]
  assign _T_3999 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@23964.4 package.scala 96:25:@23965.4]
  assign _T_4023 = _T_3999 ? Mem1D_10_io_output : _T_4022; // @[Mux.scala 31:69:@24019.4]
  assign _T_3996 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@23956.4 package.scala 96:25:@23957.4]
  assign _T_4024 = _T_3996 ? Mem1D_8_io_output : _T_4023; // @[Mux.scala 31:69:@24020.4]
  assign _T_3993 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@23948.4 package.scala 96:25:@23949.4]
  assign _T_4025 = _T_3993 ? Mem1D_6_io_output : _T_4024; // @[Mux.scala 31:69:@24021.4]
  assign _T_3990 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@23940.4 package.scala 96:25:@23941.4]
  assign _T_4026 = _T_3990 ? Mem1D_4_io_output : _T_4025; // @[Mux.scala 31:69:@24022.4]
  assign _T_3987 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@23932.4 package.scala 96:25:@23933.4]
  assign _T_4027 = _T_3987 ? Mem1D_2_io_output : _T_4026; // @[Mux.scala 31:69:@24023.4]
  assign _T_3984 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@23924.4 package.scala 96:25:@23925.4]
  assign _T_4121 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@24148.4 package.scala 96:25:@24149.4]
  assign _T_4125 = _T_4121 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24158.4]
  assign _T_4118 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@24140.4 package.scala 96:25:@24141.4]
  assign _T_4126 = _T_4118 ? Mem1D_19_io_output : _T_4125; // @[Mux.scala 31:69:@24159.4]
  assign _T_4115 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@24132.4 package.scala 96:25:@24133.4]
  assign _T_4127 = _T_4115 ? Mem1D_17_io_output : _T_4126; // @[Mux.scala 31:69:@24160.4]
  assign _T_4112 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@24124.4 package.scala 96:25:@24125.4]
  assign _T_4128 = _T_4112 ? Mem1D_15_io_output : _T_4127; // @[Mux.scala 31:69:@24161.4]
  assign _T_4109 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@24116.4 package.scala 96:25:@24117.4]
  assign _T_4129 = _T_4109 ? Mem1D_13_io_output : _T_4128; // @[Mux.scala 31:69:@24162.4]
  assign _T_4106 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@24108.4 package.scala 96:25:@24109.4]
  assign _T_4130 = _T_4106 ? Mem1D_11_io_output : _T_4129; // @[Mux.scala 31:69:@24163.4]
  assign _T_4103 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@24100.4 package.scala 96:25:@24101.4]
  assign _T_4131 = _T_4103 ? Mem1D_9_io_output : _T_4130; // @[Mux.scala 31:69:@24164.4]
  assign _T_4100 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@24092.4 package.scala 96:25:@24093.4]
  assign _T_4132 = _T_4100 ? Mem1D_7_io_output : _T_4131; // @[Mux.scala 31:69:@24165.4]
  assign _T_4097 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@24084.4 package.scala 96:25:@24085.4]
  assign _T_4133 = _T_4097 ? Mem1D_5_io_output : _T_4132; // @[Mux.scala 31:69:@24166.4]
  assign _T_4094 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@24076.4 package.scala 96:25:@24077.4]
  assign _T_4134 = _T_4094 ? Mem1D_3_io_output : _T_4133; // @[Mux.scala 31:69:@24167.4]
  assign _T_4091 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@24068.4 package.scala 96:25:@24069.4]
  assign _T_4228 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@24292.4 package.scala 96:25:@24293.4]
  assign _T_4232 = _T_4228 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24302.4]
  assign _T_4225 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@24284.4 package.scala 96:25:@24285.4]
  assign _T_4233 = _T_4225 ? Mem1D_18_io_output : _T_4232; // @[Mux.scala 31:69:@24303.4]
  assign _T_4222 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@24276.4 package.scala 96:25:@24277.4]
  assign _T_4234 = _T_4222 ? Mem1D_16_io_output : _T_4233; // @[Mux.scala 31:69:@24304.4]
  assign _T_4219 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@24268.4 package.scala 96:25:@24269.4]
  assign _T_4235 = _T_4219 ? Mem1D_14_io_output : _T_4234; // @[Mux.scala 31:69:@24305.4]
  assign _T_4216 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@24260.4 package.scala 96:25:@24261.4]
  assign _T_4236 = _T_4216 ? Mem1D_12_io_output : _T_4235; // @[Mux.scala 31:69:@24306.4]
  assign _T_4213 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@24252.4 package.scala 96:25:@24253.4]
  assign _T_4237 = _T_4213 ? Mem1D_10_io_output : _T_4236; // @[Mux.scala 31:69:@24307.4]
  assign _T_4210 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@24244.4 package.scala 96:25:@24245.4]
  assign _T_4238 = _T_4210 ? Mem1D_8_io_output : _T_4237; // @[Mux.scala 31:69:@24308.4]
  assign _T_4207 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@24236.4 package.scala 96:25:@24237.4]
  assign _T_4239 = _T_4207 ? Mem1D_6_io_output : _T_4238; // @[Mux.scala 31:69:@24309.4]
  assign _T_4204 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@24228.4 package.scala 96:25:@24229.4]
  assign _T_4240 = _T_4204 ? Mem1D_4_io_output : _T_4239; // @[Mux.scala 31:69:@24310.4]
  assign _T_4201 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@24220.4 package.scala 96:25:@24221.4]
  assign _T_4241 = _T_4201 ? Mem1D_2_io_output : _T_4240; // @[Mux.scala 31:69:@24311.4]
  assign _T_4198 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@24212.4 package.scala 96:25:@24213.4]
  assign _T_4335 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@24436.4 package.scala 96:25:@24437.4]
  assign _T_4339 = _T_4335 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24446.4]
  assign _T_4332 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@24428.4 package.scala 96:25:@24429.4]
  assign _T_4340 = _T_4332 ? Mem1D_18_io_output : _T_4339; // @[Mux.scala 31:69:@24447.4]
  assign _T_4329 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@24420.4 package.scala 96:25:@24421.4]
  assign _T_4341 = _T_4329 ? Mem1D_16_io_output : _T_4340; // @[Mux.scala 31:69:@24448.4]
  assign _T_4326 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@24412.4 package.scala 96:25:@24413.4]
  assign _T_4342 = _T_4326 ? Mem1D_14_io_output : _T_4341; // @[Mux.scala 31:69:@24449.4]
  assign _T_4323 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@24404.4 package.scala 96:25:@24405.4]
  assign _T_4343 = _T_4323 ? Mem1D_12_io_output : _T_4342; // @[Mux.scala 31:69:@24450.4]
  assign _T_4320 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@24396.4 package.scala 96:25:@24397.4]
  assign _T_4344 = _T_4320 ? Mem1D_10_io_output : _T_4343; // @[Mux.scala 31:69:@24451.4]
  assign _T_4317 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@24388.4 package.scala 96:25:@24389.4]
  assign _T_4345 = _T_4317 ? Mem1D_8_io_output : _T_4344; // @[Mux.scala 31:69:@24452.4]
  assign _T_4314 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@24380.4 package.scala 96:25:@24381.4]
  assign _T_4346 = _T_4314 ? Mem1D_6_io_output : _T_4345; // @[Mux.scala 31:69:@24453.4]
  assign _T_4311 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@24372.4 package.scala 96:25:@24373.4]
  assign _T_4347 = _T_4311 ? Mem1D_4_io_output : _T_4346; // @[Mux.scala 31:69:@24454.4]
  assign _T_4308 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@24364.4 package.scala 96:25:@24365.4]
  assign _T_4348 = _T_4308 ? Mem1D_2_io_output : _T_4347; // @[Mux.scala 31:69:@24455.4]
  assign _T_4305 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@24356.4 package.scala 96:25:@24357.4]
  assign _T_4442 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@24580.4 package.scala 96:25:@24581.4]
  assign _T_4446 = _T_4442 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24590.4]
  assign _T_4439 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@24572.4 package.scala 96:25:@24573.4]
  assign _T_4447 = _T_4439 ? Mem1D_18_io_output : _T_4446; // @[Mux.scala 31:69:@24591.4]
  assign _T_4436 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@24564.4 package.scala 96:25:@24565.4]
  assign _T_4448 = _T_4436 ? Mem1D_16_io_output : _T_4447; // @[Mux.scala 31:69:@24592.4]
  assign _T_4433 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@24556.4 package.scala 96:25:@24557.4]
  assign _T_4449 = _T_4433 ? Mem1D_14_io_output : _T_4448; // @[Mux.scala 31:69:@24593.4]
  assign _T_4430 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@24548.4 package.scala 96:25:@24549.4]
  assign _T_4450 = _T_4430 ? Mem1D_12_io_output : _T_4449; // @[Mux.scala 31:69:@24594.4]
  assign _T_4427 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@24540.4 package.scala 96:25:@24541.4]
  assign _T_4451 = _T_4427 ? Mem1D_10_io_output : _T_4450; // @[Mux.scala 31:69:@24595.4]
  assign _T_4424 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@24532.4 package.scala 96:25:@24533.4]
  assign _T_4452 = _T_4424 ? Mem1D_8_io_output : _T_4451; // @[Mux.scala 31:69:@24596.4]
  assign _T_4421 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@24524.4 package.scala 96:25:@24525.4]
  assign _T_4453 = _T_4421 ? Mem1D_6_io_output : _T_4452; // @[Mux.scala 31:69:@24597.4]
  assign _T_4418 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@24516.4 package.scala 96:25:@24517.4]
  assign _T_4454 = _T_4418 ? Mem1D_4_io_output : _T_4453; // @[Mux.scala 31:69:@24598.4]
  assign _T_4415 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@24508.4 package.scala 96:25:@24509.4]
  assign _T_4455 = _T_4415 ? Mem1D_2_io_output : _T_4454; // @[Mux.scala 31:69:@24599.4]
  assign _T_4412 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@24500.4 package.scala 96:25:@24501.4]
  assign _T_4549 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@24724.4 package.scala 96:25:@24725.4]
  assign _T_4553 = _T_4549 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24734.4]
  assign _T_4546 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@24716.4 package.scala 96:25:@24717.4]
  assign _T_4554 = _T_4546 ? Mem1D_19_io_output : _T_4553; // @[Mux.scala 31:69:@24735.4]
  assign _T_4543 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@24708.4 package.scala 96:25:@24709.4]
  assign _T_4555 = _T_4543 ? Mem1D_17_io_output : _T_4554; // @[Mux.scala 31:69:@24736.4]
  assign _T_4540 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@24700.4 package.scala 96:25:@24701.4]
  assign _T_4556 = _T_4540 ? Mem1D_15_io_output : _T_4555; // @[Mux.scala 31:69:@24737.4]
  assign _T_4537 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  assign _T_4557 = _T_4537 ? Mem1D_13_io_output : _T_4556; // @[Mux.scala 31:69:@24738.4]
  assign _T_4534 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@24684.4 package.scala 96:25:@24685.4]
  assign _T_4558 = _T_4534 ? Mem1D_11_io_output : _T_4557; // @[Mux.scala 31:69:@24739.4]
  assign _T_4531 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@24676.4 package.scala 96:25:@24677.4]
  assign _T_4559 = _T_4531 ? Mem1D_9_io_output : _T_4558; // @[Mux.scala 31:69:@24740.4]
  assign _T_4528 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@24668.4 package.scala 96:25:@24669.4]
  assign _T_4560 = _T_4528 ? Mem1D_7_io_output : _T_4559; // @[Mux.scala 31:69:@24741.4]
  assign _T_4525 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@24660.4 package.scala 96:25:@24661.4]
  assign _T_4561 = _T_4525 ? Mem1D_5_io_output : _T_4560; // @[Mux.scala 31:69:@24742.4]
  assign _T_4522 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@24652.4 package.scala 96:25:@24653.4]
  assign _T_4562 = _T_4522 ? Mem1D_3_io_output : _T_4561; // @[Mux.scala 31:69:@24743.4]
  assign _T_4519 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@24644.4 package.scala 96:25:@24645.4]
  assign _T_4656 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@24868.4 package.scala 96:25:@24869.4]
  assign _T_4660 = _T_4656 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24878.4]
  assign _T_4653 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@24860.4 package.scala 96:25:@24861.4]
  assign _T_4661 = _T_4653 ? Mem1D_18_io_output : _T_4660; // @[Mux.scala 31:69:@24879.4]
  assign _T_4650 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@24852.4 package.scala 96:25:@24853.4]
  assign _T_4662 = _T_4650 ? Mem1D_16_io_output : _T_4661; // @[Mux.scala 31:69:@24880.4]
  assign _T_4647 = RetimeWrapper_139_io_out; // @[package.scala 96:25:@24844.4 package.scala 96:25:@24845.4]
  assign _T_4663 = _T_4647 ? Mem1D_14_io_output : _T_4662; // @[Mux.scala 31:69:@24881.4]
  assign _T_4644 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@24836.4 package.scala 96:25:@24837.4]
  assign _T_4664 = _T_4644 ? Mem1D_12_io_output : _T_4663; // @[Mux.scala 31:69:@24882.4]
  assign _T_4641 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@24828.4 package.scala 96:25:@24829.4]
  assign _T_4665 = _T_4641 ? Mem1D_10_io_output : _T_4664; // @[Mux.scala 31:69:@24883.4]
  assign _T_4638 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@24820.4 package.scala 96:25:@24821.4]
  assign _T_4666 = _T_4638 ? Mem1D_8_io_output : _T_4665; // @[Mux.scala 31:69:@24884.4]
  assign _T_4635 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  assign _T_4667 = _T_4635 ? Mem1D_6_io_output : _T_4666; // @[Mux.scala 31:69:@24885.4]
  assign _T_4632 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@24804.4 package.scala 96:25:@24805.4]
  assign _T_4668 = _T_4632 ? Mem1D_4_io_output : _T_4667; // @[Mux.scala 31:69:@24886.4]
  assign _T_4629 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@24796.4 package.scala 96:25:@24797.4]
  assign _T_4669 = _T_4629 ? Mem1D_2_io_output : _T_4668; // @[Mux.scala 31:69:@24887.4]
  assign _T_4626 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@24788.4 package.scala 96:25:@24789.4]
  assign _T_4763 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@25012.4 package.scala 96:25:@25013.4]
  assign _T_4767 = _T_4763 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25022.4]
  assign _T_4760 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@25004.4 package.scala 96:25:@25005.4]
  assign _T_4768 = _T_4760 ? Mem1D_19_io_output : _T_4767; // @[Mux.scala 31:69:@25023.4]
  assign _T_4757 = RetimeWrapper_152_io_out; // @[package.scala 96:25:@24996.4 package.scala 96:25:@24997.4]
  assign _T_4769 = _T_4757 ? Mem1D_17_io_output : _T_4768; // @[Mux.scala 31:69:@25024.4]
  assign _T_4754 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@24988.4 package.scala 96:25:@24989.4]
  assign _T_4770 = _T_4754 ? Mem1D_15_io_output : _T_4769; // @[Mux.scala 31:69:@25025.4]
  assign _T_4751 = RetimeWrapper_150_io_out; // @[package.scala 96:25:@24980.4 package.scala 96:25:@24981.4]
  assign _T_4771 = _T_4751 ? Mem1D_13_io_output : _T_4770; // @[Mux.scala 31:69:@25026.4]
  assign _T_4748 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@24972.4 package.scala 96:25:@24973.4]
  assign _T_4772 = _T_4748 ? Mem1D_11_io_output : _T_4771; // @[Mux.scala 31:69:@25027.4]
  assign _T_4745 = RetimeWrapper_148_io_out; // @[package.scala 96:25:@24964.4 package.scala 96:25:@24965.4]
  assign _T_4773 = _T_4745 ? Mem1D_9_io_output : _T_4772; // @[Mux.scala 31:69:@25028.4]
  assign _T_4742 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@24956.4 package.scala 96:25:@24957.4]
  assign _T_4774 = _T_4742 ? Mem1D_7_io_output : _T_4773; // @[Mux.scala 31:69:@25029.4]
  assign _T_4739 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@24948.4 package.scala 96:25:@24949.4]
  assign _T_4775 = _T_4739 ? Mem1D_5_io_output : _T_4774; // @[Mux.scala 31:69:@25030.4]
  assign _T_4736 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@24940.4 package.scala 96:25:@24941.4]
  assign _T_4776 = _T_4736 ? Mem1D_3_io_output : _T_4775; // @[Mux.scala 31:69:@25031.4]
  assign _T_4733 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@24932.4 package.scala 96:25:@24933.4]
  assign _T_4870 = RetimeWrapper_166_io_out; // @[package.scala 96:25:@25156.4 package.scala 96:25:@25157.4]
  assign _T_4874 = _T_4870 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25166.4]
  assign _T_4867 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@25148.4 package.scala 96:25:@25149.4]
  assign _T_4875 = _T_4867 ? Mem1D_19_io_output : _T_4874; // @[Mux.scala 31:69:@25167.4]
  assign _T_4864 = RetimeWrapper_164_io_out; // @[package.scala 96:25:@25140.4 package.scala 96:25:@25141.4]
  assign _T_4876 = _T_4864 ? Mem1D_17_io_output : _T_4875; // @[Mux.scala 31:69:@25168.4]
  assign _T_4861 = RetimeWrapper_163_io_out; // @[package.scala 96:25:@25132.4 package.scala 96:25:@25133.4]
  assign _T_4877 = _T_4861 ? Mem1D_15_io_output : _T_4876; // @[Mux.scala 31:69:@25169.4]
  assign _T_4858 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@25124.4 package.scala 96:25:@25125.4]
  assign _T_4878 = _T_4858 ? Mem1D_13_io_output : _T_4877; // @[Mux.scala 31:69:@25170.4]
  assign _T_4855 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@25116.4 package.scala 96:25:@25117.4]
  assign _T_4879 = _T_4855 ? Mem1D_11_io_output : _T_4878; // @[Mux.scala 31:69:@25171.4]
  assign _T_4852 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@25108.4 package.scala 96:25:@25109.4]
  assign _T_4880 = _T_4852 ? Mem1D_9_io_output : _T_4879; // @[Mux.scala 31:69:@25172.4]
  assign _T_4849 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@25100.4 package.scala 96:25:@25101.4]
  assign _T_4881 = _T_4849 ? Mem1D_7_io_output : _T_4880; // @[Mux.scala 31:69:@25173.4]
  assign _T_4846 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@25092.4 package.scala 96:25:@25093.4]
  assign _T_4882 = _T_4846 ? Mem1D_5_io_output : _T_4881; // @[Mux.scala 31:69:@25174.4]
  assign _T_4843 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@25084.4 package.scala 96:25:@25085.4]
  assign _T_4883 = _T_4843 ? Mem1D_3_io_output : _T_4882; // @[Mux.scala 31:69:@25175.4]
  assign _T_4840 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@25076.4 package.scala 96:25:@25077.4]
  assign _T_4977 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@25300.4 package.scala 96:25:@25301.4]
  assign _T_4981 = _T_4977 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25310.4]
  assign _T_4974 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@25292.4 package.scala 96:25:@25293.4]
  assign _T_4982 = _T_4974 ? Mem1D_18_io_output : _T_4981; // @[Mux.scala 31:69:@25311.4]
  assign _T_4971 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@25284.4 package.scala 96:25:@25285.4]
  assign _T_4983 = _T_4971 ? Mem1D_16_io_output : _T_4982; // @[Mux.scala 31:69:@25312.4]
  assign _T_4968 = RetimeWrapper_175_io_out; // @[package.scala 96:25:@25276.4 package.scala 96:25:@25277.4]
  assign _T_4984 = _T_4968 ? Mem1D_14_io_output : _T_4983; // @[Mux.scala 31:69:@25313.4]
  assign _T_4965 = RetimeWrapper_174_io_out; // @[package.scala 96:25:@25268.4 package.scala 96:25:@25269.4]
  assign _T_4985 = _T_4965 ? Mem1D_12_io_output : _T_4984; // @[Mux.scala 31:69:@25314.4]
  assign _T_4962 = RetimeWrapper_173_io_out; // @[package.scala 96:25:@25260.4 package.scala 96:25:@25261.4]
  assign _T_4986 = _T_4962 ? Mem1D_10_io_output : _T_4985; // @[Mux.scala 31:69:@25315.4]
  assign _T_4959 = RetimeWrapper_172_io_out; // @[package.scala 96:25:@25252.4 package.scala 96:25:@25253.4]
  assign _T_4987 = _T_4959 ? Mem1D_8_io_output : _T_4986; // @[Mux.scala 31:69:@25316.4]
  assign _T_4956 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@25244.4 package.scala 96:25:@25245.4]
  assign _T_4988 = _T_4956 ? Mem1D_6_io_output : _T_4987; // @[Mux.scala 31:69:@25317.4]
  assign _T_4953 = RetimeWrapper_170_io_out; // @[package.scala 96:25:@25236.4 package.scala 96:25:@25237.4]
  assign _T_4989 = _T_4953 ? Mem1D_4_io_output : _T_4988; // @[Mux.scala 31:69:@25318.4]
  assign _T_4950 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@25228.4 package.scala 96:25:@25229.4]
  assign _T_4990 = _T_4950 ? Mem1D_2_io_output : _T_4989; // @[Mux.scala 31:69:@25319.4]
  assign _T_4947 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@25220.4 package.scala 96:25:@25221.4]
  assign _T_5084 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@25444.4 package.scala 96:25:@25445.4]
  assign _T_5088 = _T_5084 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25454.4]
  assign _T_5081 = RetimeWrapper_189_io_out; // @[package.scala 96:25:@25436.4 package.scala 96:25:@25437.4]
  assign _T_5089 = _T_5081 ? Mem1D_19_io_output : _T_5088; // @[Mux.scala 31:69:@25455.4]
  assign _T_5078 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@25428.4 package.scala 96:25:@25429.4]
  assign _T_5090 = _T_5078 ? Mem1D_17_io_output : _T_5089; // @[Mux.scala 31:69:@25456.4]
  assign _T_5075 = RetimeWrapper_187_io_out; // @[package.scala 96:25:@25420.4 package.scala 96:25:@25421.4]
  assign _T_5091 = _T_5075 ? Mem1D_15_io_output : _T_5090; // @[Mux.scala 31:69:@25457.4]
  assign _T_5072 = RetimeWrapper_186_io_out; // @[package.scala 96:25:@25412.4 package.scala 96:25:@25413.4]
  assign _T_5092 = _T_5072 ? Mem1D_13_io_output : _T_5091; // @[Mux.scala 31:69:@25458.4]
  assign _T_5069 = RetimeWrapper_185_io_out; // @[package.scala 96:25:@25404.4 package.scala 96:25:@25405.4]
  assign _T_5093 = _T_5069 ? Mem1D_11_io_output : _T_5092; // @[Mux.scala 31:69:@25459.4]
  assign _T_5066 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@25396.4 package.scala 96:25:@25397.4]
  assign _T_5094 = _T_5066 ? Mem1D_9_io_output : _T_5093; // @[Mux.scala 31:69:@25460.4]
  assign _T_5063 = RetimeWrapper_183_io_out; // @[package.scala 96:25:@25388.4 package.scala 96:25:@25389.4]
  assign _T_5095 = _T_5063 ? Mem1D_7_io_output : _T_5094; // @[Mux.scala 31:69:@25461.4]
  assign _T_5060 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@25380.4 package.scala 96:25:@25381.4]
  assign _T_5096 = _T_5060 ? Mem1D_5_io_output : _T_5095; // @[Mux.scala 31:69:@25462.4]
  assign _T_5057 = RetimeWrapper_181_io_out; // @[package.scala 96:25:@25372.4 package.scala 96:25:@25373.4]
  assign _T_5097 = _T_5057 ? Mem1D_3_io_output : _T_5096; // @[Mux.scala 31:69:@25463.4]
  assign _T_5054 = RetimeWrapper_180_io_out; // @[package.scala 96:25:@25364.4 package.scala 96:25:@25365.4]
  assign _T_5191 = RetimeWrapper_202_io_out; // @[package.scala 96:25:@25588.4 package.scala 96:25:@25589.4]
  assign _T_5195 = _T_5191 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25598.4]
  assign _T_5188 = RetimeWrapper_201_io_out; // @[package.scala 96:25:@25580.4 package.scala 96:25:@25581.4]
  assign _T_5196 = _T_5188 ? Mem1D_18_io_output : _T_5195; // @[Mux.scala 31:69:@25599.4]
  assign _T_5185 = RetimeWrapper_200_io_out; // @[package.scala 96:25:@25572.4 package.scala 96:25:@25573.4]
  assign _T_5197 = _T_5185 ? Mem1D_16_io_output : _T_5196; // @[Mux.scala 31:69:@25600.4]
  assign _T_5182 = RetimeWrapper_199_io_out; // @[package.scala 96:25:@25564.4 package.scala 96:25:@25565.4]
  assign _T_5198 = _T_5182 ? Mem1D_14_io_output : _T_5197; // @[Mux.scala 31:69:@25601.4]
  assign _T_5179 = RetimeWrapper_198_io_out; // @[package.scala 96:25:@25556.4 package.scala 96:25:@25557.4]
  assign _T_5199 = _T_5179 ? Mem1D_12_io_output : _T_5198; // @[Mux.scala 31:69:@25602.4]
  assign _T_5176 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@25548.4 package.scala 96:25:@25549.4]
  assign _T_5200 = _T_5176 ? Mem1D_10_io_output : _T_5199; // @[Mux.scala 31:69:@25603.4]
  assign _T_5173 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@25540.4 package.scala 96:25:@25541.4]
  assign _T_5201 = _T_5173 ? Mem1D_8_io_output : _T_5200; // @[Mux.scala 31:69:@25604.4]
  assign _T_5170 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@25532.4 package.scala 96:25:@25533.4]
  assign _T_5202 = _T_5170 ? Mem1D_6_io_output : _T_5201; // @[Mux.scala 31:69:@25605.4]
  assign _T_5167 = RetimeWrapper_194_io_out; // @[package.scala 96:25:@25524.4 package.scala 96:25:@25525.4]
  assign _T_5203 = _T_5167 ? Mem1D_4_io_output : _T_5202; // @[Mux.scala 31:69:@25606.4]
  assign _T_5164 = RetimeWrapper_193_io_out; // @[package.scala 96:25:@25516.4 package.scala 96:25:@25517.4]
  assign _T_5204 = _T_5164 ? Mem1D_2_io_output : _T_5203; // @[Mux.scala 31:69:@25607.4]
  assign _T_5161 = RetimeWrapper_192_io_out; // @[package.scala 96:25:@25508.4 package.scala 96:25:@25509.4]
  assign _T_5298 = RetimeWrapper_214_io_out; // @[package.scala 96:25:@25732.4 package.scala 96:25:@25733.4]
  assign _T_5302 = _T_5298 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25742.4]
  assign _T_5295 = RetimeWrapper_213_io_out; // @[package.scala 96:25:@25724.4 package.scala 96:25:@25725.4]
  assign _T_5303 = _T_5295 ? Mem1D_19_io_output : _T_5302; // @[Mux.scala 31:69:@25743.4]
  assign _T_5292 = RetimeWrapper_212_io_out; // @[package.scala 96:25:@25716.4 package.scala 96:25:@25717.4]
  assign _T_5304 = _T_5292 ? Mem1D_17_io_output : _T_5303; // @[Mux.scala 31:69:@25744.4]
  assign _T_5289 = RetimeWrapper_211_io_out; // @[package.scala 96:25:@25708.4 package.scala 96:25:@25709.4]
  assign _T_5305 = _T_5289 ? Mem1D_15_io_output : _T_5304; // @[Mux.scala 31:69:@25745.4]
  assign _T_5286 = RetimeWrapper_210_io_out; // @[package.scala 96:25:@25700.4 package.scala 96:25:@25701.4]
  assign _T_5306 = _T_5286 ? Mem1D_13_io_output : _T_5305; // @[Mux.scala 31:69:@25746.4]
  assign _T_5283 = RetimeWrapper_209_io_out; // @[package.scala 96:25:@25692.4 package.scala 96:25:@25693.4]
  assign _T_5307 = _T_5283 ? Mem1D_11_io_output : _T_5306; // @[Mux.scala 31:69:@25747.4]
  assign _T_5280 = RetimeWrapper_208_io_out; // @[package.scala 96:25:@25684.4 package.scala 96:25:@25685.4]
  assign _T_5308 = _T_5280 ? Mem1D_9_io_output : _T_5307; // @[Mux.scala 31:69:@25748.4]
  assign _T_5277 = RetimeWrapper_207_io_out; // @[package.scala 96:25:@25676.4 package.scala 96:25:@25677.4]
  assign _T_5309 = _T_5277 ? Mem1D_7_io_output : _T_5308; // @[Mux.scala 31:69:@25749.4]
  assign _T_5274 = RetimeWrapper_206_io_out; // @[package.scala 96:25:@25668.4 package.scala 96:25:@25669.4]
  assign _T_5310 = _T_5274 ? Mem1D_5_io_output : _T_5309; // @[Mux.scala 31:69:@25750.4]
  assign _T_5271 = RetimeWrapper_205_io_out; // @[package.scala 96:25:@25660.4 package.scala 96:25:@25661.4]
  assign _T_5311 = _T_5271 ? Mem1D_3_io_output : _T_5310; // @[Mux.scala 31:69:@25751.4]
  assign _T_5268 = RetimeWrapper_204_io_out; // @[package.scala 96:25:@25652.4 package.scala 96:25:@25653.4]
  assign io_rPort_17_output_0 = _T_5268 ? Mem1D_1_io_output : _T_5311; // @[MemPrimitives.scala 152:13:@25753.4]
  assign io_rPort_16_output_0 = _T_5161 ? Mem1D_io_output : _T_5204; // @[MemPrimitives.scala 152:13:@25609.4]
  assign io_rPort_15_output_0 = _T_5054 ? Mem1D_1_io_output : _T_5097; // @[MemPrimitives.scala 152:13:@25465.4]
  assign io_rPort_14_output_0 = _T_4947 ? Mem1D_io_output : _T_4990; // @[MemPrimitives.scala 152:13:@25321.4]
  assign io_rPort_13_output_0 = _T_4840 ? Mem1D_1_io_output : _T_4883; // @[MemPrimitives.scala 152:13:@25177.4]
  assign io_rPort_12_output_0 = _T_4733 ? Mem1D_1_io_output : _T_4776; // @[MemPrimitives.scala 152:13:@25033.4]
  assign io_rPort_11_output_0 = _T_4626 ? Mem1D_io_output : _T_4669; // @[MemPrimitives.scala 152:13:@24889.4]
  assign io_rPort_10_output_0 = _T_4519 ? Mem1D_1_io_output : _T_4562; // @[MemPrimitives.scala 152:13:@24745.4]
  assign io_rPort_9_output_0 = _T_4412 ? Mem1D_io_output : _T_4455; // @[MemPrimitives.scala 152:13:@24601.4]
  assign io_rPort_8_output_0 = _T_4305 ? Mem1D_io_output : _T_4348; // @[MemPrimitives.scala 152:13:@24457.4]
  assign io_rPort_7_output_0 = _T_4198 ? Mem1D_io_output : _T_4241; // @[MemPrimitives.scala 152:13:@24313.4]
  assign io_rPort_6_output_0 = _T_4091 ? Mem1D_1_io_output : _T_4134; // @[MemPrimitives.scala 152:13:@24169.4]
  assign io_rPort_5_output_0 = _T_3984 ? Mem1D_io_output : _T_4027; // @[MemPrimitives.scala 152:13:@24025.4]
  assign io_rPort_4_output_0 = _T_3877 ? Mem1D_1_io_output : _T_3920; // @[MemPrimitives.scala 152:13:@23881.4]
  assign io_rPort_3_output_0 = _T_3770 ? Mem1D_1_io_output : _T_3813; // @[MemPrimitives.scala 152:13:@23737.4]
  assign io_rPort_2_output_0 = _T_3663 ? Mem1D_1_io_output : _T_3706; // @[MemPrimitives.scala 152:13:@23593.4]
  assign io_rPort_1_output_0 = _T_3556 ? Mem1D_io_output : _T_3599; // @[MemPrimitives.scala 152:13:@23449.4]
  assign io_rPort_0_output_0 = _T_3449 ? Mem1D_io_output : _T_3492; // @[MemPrimitives.scala 152:13:@23305.4]
  assign Mem1D_clock = clock; // @[:@20187.4]
  assign Mem1D_reset = reset; // @[:@20188.4]
  assign Mem1D_io_r_ofs_0 = _T_1267[8:0]; // @[MemPrimitives.scala 131:28:@21112.4]
  assign Mem1D_io_r_backpressure = _T_1267[9]; // @[MemPrimitives.scala 132:32:@21113.4]
  assign Mem1D_io_w_ofs_0 = _T_715[8:0]; // @[MemPrimitives.scala 94:28:@20586.4]
  assign Mem1D_io_w_data_0 = _T_715[40:9]; // @[MemPrimitives.scala 95:29:@20587.4]
  assign Mem1D_io_w_en_0 = _T_715[41]; // @[MemPrimitives.scala 96:27:@20588.4]
  assign Mem1D_1_clock = clock; // @[:@20203.4]
  assign Mem1D_1_reset = reset; // @[:@20204.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@21201.4]
  assign Mem1D_1_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@21202.4]
  assign Mem1D_1_io_w_ofs_0 = _T_735[8:0]; // @[MemPrimitives.scala 94:28:@20605.4]
  assign Mem1D_1_io_w_data_0 = _T_735[40:9]; // @[MemPrimitives.scala 95:29:@20606.4]
  assign Mem1D_1_io_w_en_0 = _T_735[41]; // @[MemPrimitives.scala 96:27:@20607.4]
  assign Mem1D_2_clock = clock; // @[:@20219.4]
  assign Mem1D_2_reset = reset; // @[:@20220.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1451[8:0]; // @[MemPrimitives.scala 131:28:@21290.4]
  assign Mem1D_2_io_r_backpressure = _T_1451[9]; // @[MemPrimitives.scala 132:32:@21291.4]
  assign Mem1D_2_io_w_ofs_0 = _T_755[8:0]; // @[MemPrimitives.scala 94:28:@20624.4]
  assign Mem1D_2_io_w_data_0 = _T_755[40:9]; // @[MemPrimitives.scala 95:29:@20625.4]
  assign Mem1D_2_io_w_en_0 = _T_755[41]; // @[MemPrimitives.scala 96:27:@20626.4]
  assign Mem1D_3_clock = clock; // @[:@20235.4]
  assign Mem1D_3_reset = reset; // @[:@20236.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1543[8:0]; // @[MemPrimitives.scala 131:28:@21379.4]
  assign Mem1D_3_io_r_backpressure = _T_1543[9]; // @[MemPrimitives.scala 132:32:@21380.4]
  assign Mem1D_3_io_w_ofs_0 = _T_775[8:0]; // @[MemPrimitives.scala 94:28:@20643.4]
  assign Mem1D_3_io_w_data_0 = _T_775[40:9]; // @[MemPrimitives.scala 95:29:@20644.4]
  assign Mem1D_3_io_w_en_0 = _T_775[41]; // @[MemPrimitives.scala 96:27:@20645.4]
  assign Mem1D_4_clock = clock; // @[:@20251.4]
  assign Mem1D_4_reset = reset; // @[:@20252.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1635[8:0]; // @[MemPrimitives.scala 131:28:@21468.4]
  assign Mem1D_4_io_r_backpressure = _T_1635[9]; // @[MemPrimitives.scala 132:32:@21469.4]
  assign Mem1D_4_io_w_ofs_0 = _T_795[8:0]; // @[MemPrimitives.scala 94:28:@20662.4]
  assign Mem1D_4_io_w_data_0 = _T_795[40:9]; // @[MemPrimitives.scala 95:29:@20663.4]
  assign Mem1D_4_io_w_en_0 = _T_795[41]; // @[MemPrimitives.scala 96:27:@20664.4]
  assign Mem1D_5_clock = clock; // @[:@20267.4]
  assign Mem1D_5_reset = reset; // @[:@20268.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1727[8:0]; // @[MemPrimitives.scala 131:28:@21557.4]
  assign Mem1D_5_io_r_backpressure = _T_1727[9]; // @[MemPrimitives.scala 132:32:@21558.4]
  assign Mem1D_5_io_w_ofs_0 = _T_815[8:0]; // @[MemPrimitives.scala 94:28:@20681.4]
  assign Mem1D_5_io_w_data_0 = _T_815[40:9]; // @[MemPrimitives.scala 95:29:@20682.4]
  assign Mem1D_5_io_w_en_0 = _T_815[41]; // @[MemPrimitives.scala 96:27:@20683.4]
  assign Mem1D_6_clock = clock; // @[:@20283.4]
  assign Mem1D_6_reset = reset; // @[:@20284.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1819[8:0]; // @[MemPrimitives.scala 131:28:@21646.4]
  assign Mem1D_6_io_r_backpressure = _T_1819[9]; // @[MemPrimitives.scala 132:32:@21647.4]
  assign Mem1D_6_io_w_ofs_0 = _T_835[8:0]; // @[MemPrimitives.scala 94:28:@20700.4]
  assign Mem1D_6_io_w_data_0 = _T_835[40:9]; // @[MemPrimitives.scala 95:29:@20701.4]
  assign Mem1D_6_io_w_en_0 = _T_835[41]; // @[MemPrimitives.scala 96:27:@20702.4]
  assign Mem1D_7_clock = clock; // @[:@20299.4]
  assign Mem1D_7_reset = reset; // @[:@20300.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1911[8:0]; // @[MemPrimitives.scala 131:28:@21735.4]
  assign Mem1D_7_io_r_backpressure = _T_1911[9]; // @[MemPrimitives.scala 132:32:@21736.4]
  assign Mem1D_7_io_w_ofs_0 = _T_855[8:0]; // @[MemPrimitives.scala 94:28:@20719.4]
  assign Mem1D_7_io_w_data_0 = _T_855[40:9]; // @[MemPrimitives.scala 95:29:@20720.4]
  assign Mem1D_7_io_w_en_0 = _T_855[41]; // @[MemPrimitives.scala 96:27:@20721.4]
  assign Mem1D_8_clock = clock; // @[:@20315.4]
  assign Mem1D_8_reset = reset; // @[:@20316.4]
  assign Mem1D_8_io_r_ofs_0 = _T_2003[8:0]; // @[MemPrimitives.scala 131:28:@21824.4]
  assign Mem1D_8_io_r_backpressure = _T_2003[9]; // @[MemPrimitives.scala 132:32:@21825.4]
  assign Mem1D_8_io_w_ofs_0 = _T_875[8:0]; // @[MemPrimitives.scala 94:28:@20738.4]
  assign Mem1D_8_io_w_data_0 = _T_875[40:9]; // @[MemPrimitives.scala 95:29:@20739.4]
  assign Mem1D_8_io_w_en_0 = _T_875[41]; // @[MemPrimitives.scala 96:27:@20740.4]
  assign Mem1D_9_clock = clock; // @[:@20331.4]
  assign Mem1D_9_reset = reset; // @[:@20332.4]
  assign Mem1D_9_io_r_ofs_0 = _T_2095[8:0]; // @[MemPrimitives.scala 131:28:@21913.4]
  assign Mem1D_9_io_r_backpressure = _T_2095[9]; // @[MemPrimitives.scala 132:32:@21914.4]
  assign Mem1D_9_io_w_ofs_0 = _T_895[8:0]; // @[MemPrimitives.scala 94:28:@20757.4]
  assign Mem1D_9_io_w_data_0 = _T_895[40:9]; // @[MemPrimitives.scala 95:29:@20758.4]
  assign Mem1D_9_io_w_en_0 = _T_895[41]; // @[MemPrimitives.scala 96:27:@20759.4]
  assign Mem1D_10_clock = clock; // @[:@20347.4]
  assign Mem1D_10_reset = reset; // @[:@20348.4]
  assign Mem1D_10_io_r_ofs_0 = _T_2187[8:0]; // @[MemPrimitives.scala 131:28:@22002.4]
  assign Mem1D_10_io_r_backpressure = _T_2187[9]; // @[MemPrimitives.scala 132:32:@22003.4]
  assign Mem1D_10_io_w_ofs_0 = _T_915[8:0]; // @[MemPrimitives.scala 94:28:@20776.4]
  assign Mem1D_10_io_w_data_0 = _T_915[40:9]; // @[MemPrimitives.scala 95:29:@20777.4]
  assign Mem1D_10_io_w_en_0 = _T_915[41]; // @[MemPrimitives.scala 96:27:@20778.4]
  assign Mem1D_11_clock = clock; // @[:@20363.4]
  assign Mem1D_11_reset = reset; // @[:@20364.4]
  assign Mem1D_11_io_r_ofs_0 = _T_2279[8:0]; // @[MemPrimitives.scala 131:28:@22091.4]
  assign Mem1D_11_io_r_backpressure = _T_2279[9]; // @[MemPrimitives.scala 132:32:@22092.4]
  assign Mem1D_11_io_w_ofs_0 = _T_935[8:0]; // @[MemPrimitives.scala 94:28:@20795.4]
  assign Mem1D_11_io_w_data_0 = _T_935[40:9]; // @[MemPrimitives.scala 95:29:@20796.4]
  assign Mem1D_11_io_w_en_0 = _T_935[41]; // @[MemPrimitives.scala 96:27:@20797.4]
  assign Mem1D_12_clock = clock; // @[:@20379.4]
  assign Mem1D_12_reset = reset; // @[:@20380.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2371[8:0]; // @[MemPrimitives.scala 131:28:@22180.4]
  assign Mem1D_12_io_r_backpressure = _T_2371[9]; // @[MemPrimitives.scala 132:32:@22181.4]
  assign Mem1D_12_io_w_ofs_0 = _T_955[8:0]; // @[MemPrimitives.scala 94:28:@20814.4]
  assign Mem1D_12_io_w_data_0 = _T_955[40:9]; // @[MemPrimitives.scala 95:29:@20815.4]
  assign Mem1D_12_io_w_en_0 = _T_955[41]; // @[MemPrimitives.scala 96:27:@20816.4]
  assign Mem1D_13_clock = clock; // @[:@20395.4]
  assign Mem1D_13_reset = reset; // @[:@20396.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2463[8:0]; // @[MemPrimitives.scala 131:28:@22269.4]
  assign Mem1D_13_io_r_backpressure = _T_2463[9]; // @[MemPrimitives.scala 132:32:@22270.4]
  assign Mem1D_13_io_w_ofs_0 = _T_975[8:0]; // @[MemPrimitives.scala 94:28:@20833.4]
  assign Mem1D_13_io_w_data_0 = _T_975[40:9]; // @[MemPrimitives.scala 95:29:@20834.4]
  assign Mem1D_13_io_w_en_0 = _T_975[41]; // @[MemPrimitives.scala 96:27:@20835.4]
  assign Mem1D_14_clock = clock; // @[:@20411.4]
  assign Mem1D_14_reset = reset; // @[:@20412.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2555[8:0]; // @[MemPrimitives.scala 131:28:@22358.4]
  assign Mem1D_14_io_r_backpressure = _T_2555[9]; // @[MemPrimitives.scala 132:32:@22359.4]
  assign Mem1D_14_io_w_ofs_0 = _T_995[8:0]; // @[MemPrimitives.scala 94:28:@20852.4]
  assign Mem1D_14_io_w_data_0 = _T_995[40:9]; // @[MemPrimitives.scala 95:29:@20853.4]
  assign Mem1D_14_io_w_en_0 = _T_995[41]; // @[MemPrimitives.scala 96:27:@20854.4]
  assign Mem1D_15_clock = clock; // @[:@20427.4]
  assign Mem1D_15_reset = reset; // @[:@20428.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2647[8:0]; // @[MemPrimitives.scala 131:28:@22447.4]
  assign Mem1D_15_io_r_backpressure = _T_2647[9]; // @[MemPrimitives.scala 132:32:@22448.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1015[8:0]; // @[MemPrimitives.scala 94:28:@20871.4]
  assign Mem1D_15_io_w_data_0 = _T_1015[40:9]; // @[MemPrimitives.scala 95:29:@20872.4]
  assign Mem1D_15_io_w_en_0 = _T_1015[41]; // @[MemPrimitives.scala 96:27:@20873.4]
  assign Mem1D_16_clock = clock; // @[:@20443.4]
  assign Mem1D_16_reset = reset; // @[:@20444.4]
  assign Mem1D_16_io_r_ofs_0 = _T_2739[8:0]; // @[MemPrimitives.scala 131:28:@22536.4]
  assign Mem1D_16_io_r_backpressure = _T_2739[9]; // @[MemPrimitives.scala 132:32:@22537.4]
  assign Mem1D_16_io_w_ofs_0 = _T_1035[8:0]; // @[MemPrimitives.scala 94:28:@20890.4]
  assign Mem1D_16_io_w_data_0 = _T_1035[40:9]; // @[MemPrimitives.scala 95:29:@20891.4]
  assign Mem1D_16_io_w_en_0 = _T_1035[41]; // @[MemPrimitives.scala 96:27:@20892.4]
  assign Mem1D_17_clock = clock; // @[:@20459.4]
  assign Mem1D_17_reset = reset; // @[:@20460.4]
  assign Mem1D_17_io_r_ofs_0 = _T_2831[8:0]; // @[MemPrimitives.scala 131:28:@22625.4]
  assign Mem1D_17_io_r_backpressure = _T_2831[9]; // @[MemPrimitives.scala 132:32:@22626.4]
  assign Mem1D_17_io_w_ofs_0 = _T_1055[8:0]; // @[MemPrimitives.scala 94:28:@20909.4]
  assign Mem1D_17_io_w_data_0 = _T_1055[40:9]; // @[MemPrimitives.scala 95:29:@20910.4]
  assign Mem1D_17_io_w_en_0 = _T_1055[41]; // @[MemPrimitives.scala 96:27:@20911.4]
  assign Mem1D_18_clock = clock; // @[:@20475.4]
  assign Mem1D_18_reset = reset; // @[:@20476.4]
  assign Mem1D_18_io_r_ofs_0 = _T_2923[8:0]; // @[MemPrimitives.scala 131:28:@22714.4]
  assign Mem1D_18_io_r_backpressure = _T_2923[9]; // @[MemPrimitives.scala 132:32:@22715.4]
  assign Mem1D_18_io_w_ofs_0 = _T_1075[8:0]; // @[MemPrimitives.scala 94:28:@20928.4]
  assign Mem1D_18_io_w_data_0 = _T_1075[40:9]; // @[MemPrimitives.scala 95:29:@20929.4]
  assign Mem1D_18_io_w_en_0 = _T_1075[41]; // @[MemPrimitives.scala 96:27:@20930.4]
  assign Mem1D_19_clock = clock; // @[:@20491.4]
  assign Mem1D_19_reset = reset; // @[:@20492.4]
  assign Mem1D_19_io_r_ofs_0 = _T_3015[8:0]; // @[MemPrimitives.scala 131:28:@22803.4]
  assign Mem1D_19_io_r_backpressure = _T_3015[9]; // @[MemPrimitives.scala 132:32:@22804.4]
  assign Mem1D_19_io_w_ofs_0 = _T_1095[8:0]; // @[MemPrimitives.scala 94:28:@20947.4]
  assign Mem1D_19_io_w_data_0 = _T_1095[40:9]; // @[MemPrimitives.scala 95:29:@20948.4]
  assign Mem1D_19_io_w_en_0 = _T_1095[41]; // @[MemPrimitives.scala 96:27:@20949.4]
  assign Mem1D_20_clock = clock; // @[:@20507.4]
  assign Mem1D_20_reset = reset; // @[:@20508.4]
  assign Mem1D_20_io_r_ofs_0 = _T_3107[8:0]; // @[MemPrimitives.scala 131:28:@22892.4]
  assign Mem1D_20_io_r_backpressure = _T_3107[9]; // @[MemPrimitives.scala 132:32:@22893.4]
  assign Mem1D_20_io_w_ofs_0 = _T_1115[8:0]; // @[MemPrimitives.scala 94:28:@20966.4]
  assign Mem1D_20_io_w_data_0 = _T_1115[40:9]; // @[MemPrimitives.scala 95:29:@20967.4]
  assign Mem1D_20_io_w_en_0 = _T_1115[41]; // @[MemPrimitives.scala 96:27:@20968.4]
  assign Mem1D_21_clock = clock; // @[:@20523.4]
  assign Mem1D_21_reset = reset; // @[:@20524.4]
  assign Mem1D_21_io_r_ofs_0 = _T_3199[8:0]; // @[MemPrimitives.scala 131:28:@22981.4]
  assign Mem1D_21_io_r_backpressure = _T_3199[9]; // @[MemPrimitives.scala 132:32:@22982.4]
  assign Mem1D_21_io_w_ofs_0 = _T_1135[8:0]; // @[MemPrimitives.scala 94:28:@20985.4]
  assign Mem1D_21_io_w_data_0 = _T_1135[40:9]; // @[MemPrimitives.scala 95:29:@20986.4]
  assign Mem1D_21_io_w_en_0 = _T_1135[41]; // @[MemPrimitives.scala 96:27:@20987.4]
  assign Mem1D_22_clock = clock; // @[:@20539.4]
  assign Mem1D_22_reset = reset; // @[:@20540.4]
  assign Mem1D_22_io_r_ofs_0 = _T_3291[8:0]; // @[MemPrimitives.scala 131:28:@23070.4]
  assign Mem1D_22_io_r_backpressure = _T_3291[9]; // @[MemPrimitives.scala 132:32:@23071.4]
  assign Mem1D_22_io_w_ofs_0 = _T_1155[8:0]; // @[MemPrimitives.scala 94:28:@21004.4]
  assign Mem1D_22_io_w_data_0 = _T_1155[40:9]; // @[MemPrimitives.scala 95:29:@21005.4]
  assign Mem1D_22_io_w_en_0 = _T_1155[41]; // @[MemPrimitives.scala 96:27:@21006.4]
  assign Mem1D_23_clock = clock; // @[:@20555.4]
  assign Mem1D_23_reset = reset; // @[:@20556.4]
  assign Mem1D_23_io_r_ofs_0 = _T_3383[8:0]; // @[MemPrimitives.scala 131:28:@23159.4]
  assign Mem1D_23_io_r_backpressure = _T_3383[9]; // @[MemPrimitives.scala 132:32:@23160.4]
  assign Mem1D_23_io_w_ofs_0 = _T_1175[8:0]; // @[MemPrimitives.scala 94:28:@21023.4]
  assign Mem1D_23_io_w_data_0 = _T_1175[40:9]; // @[MemPrimitives.scala 95:29:@21024.4]
  assign Mem1D_23_io_w_en_0 = _T_1175[41]; // @[MemPrimitives.scala 96:27:@21025.4]
  assign StickySelects_clock = clock; // @[:@21063.4]
  assign StickySelects_reset = reset; // @[:@21064.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_1183; // @[MemPrimitives.scala 125:64:@21065.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_1189; // @[MemPrimitives.scala 125:64:@21066.4]
  assign StickySelects_io_ins_2 = io_rPort_5_en_0 & _T_1195; // @[MemPrimitives.scala 125:64:@21067.4]
  assign StickySelects_io_ins_3 = io_rPort_7_en_0 & _T_1201; // @[MemPrimitives.scala 125:64:@21068.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_1207; // @[MemPrimitives.scala 125:64:@21069.4]
  assign StickySelects_io_ins_5 = io_rPort_9_en_0 & _T_1213; // @[MemPrimitives.scala 125:64:@21070.4]
  assign StickySelects_io_ins_6 = io_rPort_11_en_0 & _T_1219; // @[MemPrimitives.scala 125:64:@21071.4]
  assign StickySelects_io_ins_7 = io_rPort_14_en_0 & _T_1225; // @[MemPrimitives.scala 125:64:@21072.4]
  assign StickySelects_io_ins_8 = io_rPort_16_en_0 & _T_1231; // @[MemPrimitives.scala 125:64:@21073.4]
  assign StickySelects_1_clock = clock; // @[:@21152.4]
  assign StickySelects_1_reset = reset; // @[:@21153.4]
  assign StickySelects_1_io_ins_0 = io_rPort_2_en_0 & _T_1275; // @[MemPrimitives.scala 125:64:@21154.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_1281; // @[MemPrimitives.scala 125:64:@21155.4]
  assign StickySelects_1_io_ins_2 = io_rPort_4_en_0 & _T_1287; // @[MemPrimitives.scala 125:64:@21156.4]
  assign StickySelects_1_io_ins_3 = io_rPort_6_en_0 & _T_1293; // @[MemPrimitives.scala 125:64:@21157.4]
  assign StickySelects_1_io_ins_4 = io_rPort_10_en_0 & _T_1299; // @[MemPrimitives.scala 125:64:@21158.4]
  assign StickySelects_1_io_ins_5 = io_rPort_12_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@21159.4]
  assign StickySelects_1_io_ins_6 = io_rPort_13_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@21160.4]
  assign StickySelects_1_io_ins_7 = io_rPort_15_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@21161.4]
  assign StickySelects_1_io_ins_8 = io_rPort_17_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@21162.4]
  assign StickySelects_2_clock = clock; // @[:@21241.4]
  assign StickySelects_2_reset = reset; // @[:@21242.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@21243.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@21244.4]
  assign StickySelects_2_io_ins_2 = io_rPort_5_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@21245.4]
  assign StickySelects_2_io_ins_3 = io_rPort_7_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@21246.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@21247.4]
  assign StickySelects_2_io_ins_5 = io_rPort_9_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@21248.4]
  assign StickySelects_2_io_ins_6 = io_rPort_11_en_0 & _T_1403; // @[MemPrimitives.scala 125:64:@21249.4]
  assign StickySelects_2_io_ins_7 = io_rPort_14_en_0 & _T_1409; // @[MemPrimitives.scala 125:64:@21250.4]
  assign StickySelects_2_io_ins_8 = io_rPort_16_en_0 & _T_1415; // @[MemPrimitives.scala 125:64:@21251.4]
  assign StickySelects_3_clock = clock; // @[:@21330.4]
  assign StickySelects_3_reset = reset; // @[:@21331.4]
  assign StickySelects_3_io_ins_0 = io_rPort_2_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@21332.4]
  assign StickySelects_3_io_ins_1 = io_rPort_3_en_0 & _T_1465; // @[MemPrimitives.scala 125:64:@21333.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_1471; // @[MemPrimitives.scala 125:64:@21334.4]
  assign StickySelects_3_io_ins_3 = io_rPort_6_en_0 & _T_1477; // @[MemPrimitives.scala 125:64:@21335.4]
  assign StickySelects_3_io_ins_4 = io_rPort_10_en_0 & _T_1483; // @[MemPrimitives.scala 125:64:@21336.4]
  assign StickySelects_3_io_ins_5 = io_rPort_12_en_0 & _T_1489; // @[MemPrimitives.scala 125:64:@21337.4]
  assign StickySelects_3_io_ins_6 = io_rPort_13_en_0 & _T_1495; // @[MemPrimitives.scala 125:64:@21338.4]
  assign StickySelects_3_io_ins_7 = io_rPort_15_en_0 & _T_1501; // @[MemPrimitives.scala 125:64:@21339.4]
  assign StickySelects_3_io_ins_8 = io_rPort_17_en_0 & _T_1507; // @[MemPrimitives.scala 125:64:@21340.4]
  assign StickySelects_4_clock = clock; // @[:@21419.4]
  assign StickySelects_4_reset = reset; // @[:@21420.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_1551; // @[MemPrimitives.scala 125:64:@21421.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_1557; // @[MemPrimitives.scala 125:64:@21422.4]
  assign StickySelects_4_io_ins_2 = io_rPort_5_en_0 & _T_1563; // @[MemPrimitives.scala 125:64:@21423.4]
  assign StickySelects_4_io_ins_3 = io_rPort_7_en_0 & _T_1569; // @[MemPrimitives.scala 125:64:@21424.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_1575; // @[MemPrimitives.scala 125:64:@21425.4]
  assign StickySelects_4_io_ins_5 = io_rPort_9_en_0 & _T_1581; // @[MemPrimitives.scala 125:64:@21426.4]
  assign StickySelects_4_io_ins_6 = io_rPort_11_en_0 & _T_1587; // @[MemPrimitives.scala 125:64:@21427.4]
  assign StickySelects_4_io_ins_7 = io_rPort_14_en_0 & _T_1593; // @[MemPrimitives.scala 125:64:@21428.4]
  assign StickySelects_4_io_ins_8 = io_rPort_16_en_0 & _T_1599; // @[MemPrimitives.scala 125:64:@21429.4]
  assign StickySelects_5_clock = clock; // @[:@21508.4]
  assign StickySelects_5_reset = reset; // @[:@21509.4]
  assign StickySelects_5_io_ins_0 = io_rPort_2_en_0 & _T_1643; // @[MemPrimitives.scala 125:64:@21510.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_1649; // @[MemPrimitives.scala 125:64:@21511.4]
  assign StickySelects_5_io_ins_2 = io_rPort_4_en_0 & _T_1655; // @[MemPrimitives.scala 125:64:@21512.4]
  assign StickySelects_5_io_ins_3 = io_rPort_6_en_0 & _T_1661; // @[MemPrimitives.scala 125:64:@21513.4]
  assign StickySelects_5_io_ins_4 = io_rPort_10_en_0 & _T_1667; // @[MemPrimitives.scala 125:64:@21514.4]
  assign StickySelects_5_io_ins_5 = io_rPort_12_en_0 & _T_1673; // @[MemPrimitives.scala 125:64:@21515.4]
  assign StickySelects_5_io_ins_6 = io_rPort_13_en_0 & _T_1679; // @[MemPrimitives.scala 125:64:@21516.4]
  assign StickySelects_5_io_ins_7 = io_rPort_15_en_0 & _T_1685; // @[MemPrimitives.scala 125:64:@21517.4]
  assign StickySelects_5_io_ins_8 = io_rPort_17_en_0 & _T_1691; // @[MemPrimitives.scala 125:64:@21518.4]
  assign StickySelects_6_clock = clock; // @[:@21597.4]
  assign StickySelects_6_reset = reset; // @[:@21598.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1735; // @[MemPrimitives.scala 125:64:@21599.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1741; // @[MemPrimitives.scala 125:64:@21600.4]
  assign StickySelects_6_io_ins_2 = io_rPort_5_en_0 & _T_1747; // @[MemPrimitives.scala 125:64:@21601.4]
  assign StickySelects_6_io_ins_3 = io_rPort_7_en_0 & _T_1753; // @[MemPrimitives.scala 125:64:@21602.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1759; // @[MemPrimitives.scala 125:64:@21603.4]
  assign StickySelects_6_io_ins_5 = io_rPort_9_en_0 & _T_1765; // @[MemPrimitives.scala 125:64:@21604.4]
  assign StickySelects_6_io_ins_6 = io_rPort_11_en_0 & _T_1771; // @[MemPrimitives.scala 125:64:@21605.4]
  assign StickySelects_6_io_ins_7 = io_rPort_14_en_0 & _T_1777; // @[MemPrimitives.scala 125:64:@21606.4]
  assign StickySelects_6_io_ins_8 = io_rPort_16_en_0 & _T_1783; // @[MemPrimitives.scala 125:64:@21607.4]
  assign StickySelects_7_clock = clock; // @[:@21686.4]
  assign StickySelects_7_reset = reset; // @[:@21687.4]
  assign StickySelects_7_io_ins_0 = io_rPort_2_en_0 & _T_1827; // @[MemPrimitives.scala 125:64:@21688.4]
  assign StickySelects_7_io_ins_1 = io_rPort_3_en_0 & _T_1833; // @[MemPrimitives.scala 125:64:@21689.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_1839; // @[MemPrimitives.scala 125:64:@21690.4]
  assign StickySelects_7_io_ins_3 = io_rPort_6_en_0 & _T_1845; // @[MemPrimitives.scala 125:64:@21691.4]
  assign StickySelects_7_io_ins_4 = io_rPort_10_en_0 & _T_1851; // @[MemPrimitives.scala 125:64:@21692.4]
  assign StickySelects_7_io_ins_5 = io_rPort_12_en_0 & _T_1857; // @[MemPrimitives.scala 125:64:@21693.4]
  assign StickySelects_7_io_ins_6 = io_rPort_13_en_0 & _T_1863; // @[MemPrimitives.scala 125:64:@21694.4]
  assign StickySelects_7_io_ins_7 = io_rPort_15_en_0 & _T_1869; // @[MemPrimitives.scala 125:64:@21695.4]
  assign StickySelects_7_io_ins_8 = io_rPort_17_en_0 & _T_1875; // @[MemPrimitives.scala 125:64:@21696.4]
  assign StickySelects_8_clock = clock; // @[:@21775.4]
  assign StickySelects_8_reset = reset; // @[:@21776.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1919; // @[MemPrimitives.scala 125:64:@21777.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1925; // @[MemPrimitives.scala 125:64:@21778.4]
  assign StickySelects_8_io_ins_2 = io_rPort_5_en_0 & _T_1931; // @[MemPrimitives.scala 125:64:@21779.4]
  assign StickySelects_8_io_ins_3 = io_rPort_7_en_0 & _T_1937; // @[MemPrimitives.scala 125:64:@21780.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1943; // @[MemPrimitives.scala 125:64:@21781.4]
  assign StickySelects_8_io_ins_5 = io_rPort_9_en_0 & _T_1949; // @[MemPrimitives.scala 125:64:@21782.4]
  assign StickySelects_8_io_ins_6 = io_rPort_11_en_0 & _T_1955; // @[MemPrimitives.scala 125:64:@21783.4]
  assign StickySelects_8_io_ins_7 = io_rPort_14_en_0 & _T_1961; // @[MemPrimitives.scala 125:64:@21784.4]
  assign StickySelects_8_io_ins_8 = io_rPort_16_en_0 & _T_1967; // @[MemPrimitives.scala 125:64:@21785.4]
  assign StickySelects_9_clock = clock; // @[:@21864.4]
  assign StickySelects_9_reset = reset; // @[:@21865.4]
  assign StickySelects_9_io_ins_0 = io_rPort_2_en_0 & _T_2011; // @[MemPrimitives.scala 125:64:@21866.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_2017; // @[MemPrimitives.scala 125:64:@21867.4]
  assign StickySelects_9_io_ins_2 = io_rPort_4_en_0 & _T_2023; // @[MemPrimitives.scala 125:64:@21868.4]
  assign StickySelects_9_io_ins_3 = io_rPort_6_en_0 & _T_2029; // @[MemPrimitives.scala 125:64:@21869.4]
  assign StickySelects_9_io_ins_4 = io_rPort_10_en_0 & _T_2035; // @[MemPrimitives.scala 125:64:@21870.4]
  assign StickySelects_9_io_ins_5 = io_rPort_12_en_0 & _T_2041; // @[MemPrimitives.scala 125:64:@21871.4]
  assign StickySelects_9_io_ins_6 = io_rPort_13_en_0 & _T_2047; // @[MemPrimitives.scala 125:64:@21872.4]
  assign StickySelects_9_io_ins_7 = io_rPort_15_en_0 & _T_2053; // @[MemPrimitives.scala 125:64:@21873.4]
  assign StickySelects_9_io_ins_8 = io_rPort_17_en_0 & _T_2059; // @[MemPrimitives.scala 125:64:@21874.4]
  assign StickySelects_10_clock = clock; // @[:@21953.4]
  assign StickySelects_10_reset = reset; // @[:@21954.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_2103; // @[MemPrimitives.scala 125:64:@21955.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_2109; // @[MemPrimitives.scala 125:64:@21956.4]
  assign StickySelects_10_io_ins_2 = io_rPort_5_en_0 & _T_2115; // @[MemPrimitives.scala 125:64:@21957.4]
  assign StickySelects_10_io_ins_3 = io_rPort_7_en_0 & _T_2121; // @[MemPrimitives.scala 125:64:@21958.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_2127; // @[MemPrimitives.scala 125:64:@21959.4]
  assign StickySelects_10_io_ins_5 = io_rPort_9_en_0 & _T_2133; // @[MemPrimitives.scala 125:64:@21960.4]
  assign StickySelects_10_io_ins_6 = io_rPort_11_en_0 & _T_2139; // @[MemPrimitives.scala 125:64:@21961.4]
  assign StickySelects_10_io_ins_7 = io_rPort_14_en_0 & _T_2145; // @[MemPrimitives.scala 125:64:@21962.4]
  assign StickySelects_10_io_ins_8 = io_rPort_16_en_0 & _T_2151; // @[MemPrimitives.scala 125:64:@21963.4]
  assign StickySelects_11_clock = clock; // @[:@22042.4]
  assign StickySelects_11_reset = reset; // @[:@22043.4]
  assign StickySelects_11_io_ins_0 = io_rPort_2_en_0 & _T_2195; // @[MemPrimitives.scala 125:64:@22044.4]
  assign StickySelects_11_io_ins_1 = io_rPort_3_en_0 & _T_2201; // @[MemPrimitives.scala 125:64:@22045.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_2207; // @[MemPrimitives.scala 125:64:@22046.4]
  assign StickySelects_11_io_ins_3 = io_rPort_6_en_0 & _T_2213; // @[MemPrimitives.scala 125:64:@22047.4]
  assign StickySelects_11_io_ins_4 = io_rPort_10_en_0 & _T_2219; // @[MemPrimitives.scala 125:64:@22048.4]
  assign StickySelects_11_io_ins_5 = io_rPort_12_en_0 & _T_2225; // @[MemPrimitives.scala 125:64:@22049.4]
  assign StickySelects_11_io_ins_6 = io_rPort_13_en_0 & _T_2231; // @[MemPrimitives.scala 125:64:@22050.4]
  assign StickySelects_11_io_ins_7 = io_rPort_15_en_0 & _T_2237; // @[MemPrimitives.scala 125:64:@22051.4]
  assign StickySelects_11_io_ins_8 = io_rPort_17_en_0 & _T_2243; // @[MemPrimitives.scala 125:64:@22052.4]
  assign StickySelects_12_clock = clock; // @[:@22131.4]
  assign StickySelects_12_reset = reset; // @[:@22132.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_2287; // @[MemPrimitives.scala 125:64:@22133.4]
  assign StickySelects_12_io_ins_1 = io_rPort_1_en_0 & _T_2293; // @[MemPrimitives.scala 125:64:@22134.4]
  assign StickySelects_12_io_ins_2 = io_rPort_5_en_0 & _T_2299; // @[MemPrimitives.scala 125:64:@22135.4]
  assign StickySelects_12_io_ins_3 = io_rPort_7_en_0 & _T_2305; // @[MemPrimitives.scala 125:64:@22136.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_2311; // @[MemPrimitives.scala 125:64:@22137.4]
  assign StickySelects_12_io_ins_5 = io_rPort_9_en_0 & _T_2317; // @[MemPrimitives.scala 125:64:@22138.4]
  assign StickySelects_12_io_ins_6 = io_rPort_11_en_0 & _T_2323; // @[MemPrimitives.scala 125:64:@22139.4]
  assign StickySelects_12_io_ins_7 = io_rPort_14_en_0 & _T_2329; // @[MemPrimitives.scala 125:64:@22140.4]
  assign StickySelects_12_io_ins_8 = io_rPort_16_en_0 & _T_2335; // @[MemPrimitives.scala 125:64:@22141.4]
  assign StickySelects_13_clock = clock; // @[:@22220.4]
  assign StickySelects_13_reset = reset; // @[:@22221.4]
  assign StickySelects_13_io_ins_0 = io_rPort_2_en_0 & _T_2379; // @[MemPrimitives.scala 125:64:@22222.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_2385; // @[MemPrimitives.scala 125:64:@22223.4]
  assign StickySelects_13_io_ins_2 = io_rPort_4_en_0 & _T_2391; // @[MemPrimitives.scala 125:64:@22224.4]
  assign StickySelects_13_io_ins_3 = io_rPort_6_en_0 & _T_2397; // @[MemPrimitives.scala 125:64:@22225.4]
  assign StickySelects_13_io_ins_4 = io_rPort_10_en_0 & _T_2403; // @[MemPrimitives.scala 125:64:@22226.4]
  assign StickySelects_13_io_ins_5 = io_rPort_12_en_0 & _T_2409; // @[MemPrimitives.scala 125:64:@22227.4]
  assign StickySelects_13_io_ins_6 = io_rPort_13_en_0 & _T_2415; // @[MemPrimitives.scala 125:64:@22228.4]
  assign StickySelects_13_io_ins_7 = io_rPort_15_en_0 & _T_2421; // @[MemPrimitives.scala 125:64:@22229.4]
  assign StickySelects_13_io_ins_8 = io_rPort_17_en_0 & _T_2427; // @[MemPrimitives.scala 125:64:@22230.4]
  assign StickySelects_14_clock = clock; // @[:@22309.4]
  assign StickySelects_14_reset = reset; // @[:@22310.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_2471; // @[MemPrimitives.scala 125:64:@22311.4]
  assign StickySelects_14_io_ins_1 = io_rPort_1_en_0 & _T_2477; // @[MemPrimitives.scala 125:64:@22312.4]
  assign StickySelects_14_io_ins_2 = io_rPort_5_en_0 & _T_2483; // @[MemPrimitives.scala 125:64:@22313.4]
  assign StickySelects_14_io_ins_3 = io_rPort_7_en_0 & _T_2489; // @[MemPrimitives.scala 125:64:@22314.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_2495; // @[MemPrimitives.scala 125:64:@22315.4]
  assign StickySelects_14_io_ins_5 = io_rPort_9_en_0 & _T_2501; // @[MemPrimitives.scala 125:64:@22316.4]
  assign StickySelects_14_io_ins_6 = io_rPort_11_en_0 & _T_2507; // @[MemPrimitives.scala 125:64:@22317.4]
  assign StickySelects_14_io_ins_7 = io_rPort_14_en_0 & _T_2513; // @[MemPrimitives.scala 125:64:@22318.4]
  assign StickySelects_14_io_ins_8 = io_rPort_16_en_0 & _T_2519; // @[MemPrimitives.scala 125:64:@22319.4]
  assign StickySelects_15_clock = clock; // @[:@22398.4]
  assign StickySelects_15_reset = reset; // @[:@22399.4]
  assign StickySelects_15_io_ins_0 = io_rPort_2_en_0 & _T_2563; // @[MemPrimitives.scala 125:64:@22400.4]
  assign StickySelects_15_io_ins_1 = io_rPort_3_en_0 & _T_2569; // @[MemPrimitives.scala 125:64:@22401.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_2575; // @[MemPrimitives.scala 125:64:@22402.4]
  assign StickySelects_15_io_ins_3 = io_rPort_6_en_0 & _T_2581; // @[MemPrimitives.scala 125:64:@22403.4]
  assign StickySelects_15_io_ins_4 = io_rPort_10_en_0 & _T_2587; // @[MemPrimitives.scala 125:64:@22404.4]
  assign StickySelects_15_io_ins_5 = io_rPort_12_en_0 & _T_2593; // @[MemPrimitives.scala 125:64:@22405.4]
  assign StickySelects_15_io_ins_6 = io_rPort_13_en_0 & _T_2599; // @[MemPrimitives.scala 125:64:@22406.4]
  assign StickySelects_15_io_ins_7 = io_rPort_15_en_0 & _T_2605; // @[MemPrimitives.scala 125:64:@22407.4]
  assign StickySelects_15_io_ins_8 = io_rPort_17_en_0 & _T_2611; // @[MemPrimitives.scala 125:64:@22408.4]
  assign StickySelects_16_clock = clock; // @[:@22487.4]
  assign StickySelects_16_reset = reset; // @[:@22488.4]
  assign StickySelects_16_io_ins_0 = io_rPort_0_en_0 & _T_2655; // @[MemPrimitives.scala 125:64:@22489.4]
  assign StickySelects_16_io_ins_1 = io_rPort_1_en_0 & _T_2661; // @[MemPrimitives.scala 125:64:@22490.4]
  assign StickySelects_16_io_ins_2 = io_rPort_5_en_0 & _T_2667; // @[MemPrimitives.scala 125:64:@22491.4]
  assign StickySelects_16_io_ins_3 = io_rPort_7_en_0 & _T_2673; // @[MemPrimitives.scala 125:64:@22492.4]
  assign StickySelects_16_io_ins_4 = io_rPort_8_en_0 & _T_2679; // @[MemPrimitives.scala 125:64:@22493.4]
  assign StickySelects_16_io_ins_5 = io_rPort_9_en_0 & _T_2685; // @[MemPrimitives.scala 125:64:@22494.4]
  assign StickySelects_16_io_ins_6 = io_rPort_11_en_0 & _T_2691; // @[MemPrimitives.scala 125:64:@22495.4]
  assign StickySelects_16_io_ins_7 = io_rPort_14_en_0 & _T_2697; // @[MemPrimitives.scala 125:64:@22496.4]
  assign StickySelects_16_io_ins_8 = io_rPort_16_en_0 & _T_2703; // @[MemPrimitives.scala 125:64:@22497.4]
  assign StickySelects_17_clock = clock; // @[:@22576.4]
  assign StickySelects_17_reset = reset; // @[:@22577.4]
  assign StickySelects_17_io_ins_0 = io_rPort_2_en_0 & _T_2747; // @[MemPrimitives.scala 125:64:@22578.4]
  assign StickySelects_17_io_ins_1 = io_rPort_3_en_0 & _T_2753; // @[MemPrimitives.scala 125:64:@22579.4]
  assign StickySelects_17_io_ins_2 = io_rPort_4_en_0 & _T_2759; // @[MemPrimitives.scala 125:64:@22580.4]
  assign StickySelects_17_io_ins_3 = io_rPort_6_en_0 & _T_2765; // @[MemPrimitives.scala 125:64:@22581.4]
  assign StickySelects_17_io_ins_4 = io_rPort_10_en_0 & _T_2771; // @[MemPrimitives.scala 125:64:@22582.4]
  assign StickySelects_17_io_ins_5 = io_rPort_12_en_0 & _T_2777; // @[MemPrimitives.scala 125:64:@22583.4]
  assign StickySelects_17_io_ins_6 = io_rPort_13_en_0 & _T_2783; // @[MemPrimitives.scala 125:64:@22584.4]
  assign StickySelects_17_io_ins_7 = io_rPort_15_en_0 & _T_2789; // @[MemPrimitives.scala 125:64:@22585.4]
  assign StickySelects_17_io_ins_8 = io_rPort_17_en_0 & _T_2795; // @[MemPrimitives.scala 125:64:@22586.4]
  assign StickySelects_18_clock = clock; // @[:@22665.4]
  assign StickySelects_18_reset = reset; // @[:@22666.4]
  assign StickySelects_18_io_ins_0 = io_rPort_0_en_0 & _T_2839; // @[MemPrimitives.scala 125:64:@22667.4]
  assign StickySelects_18_io_ins_1 = io_rPort_1_en_0 & _T_2845; // @[MemPrimitives.scala 125:64:@22668.4]
  assign StickySelects_18_io_ins_2 = io_rPort_5_en_0 & _T_2851; // @[MemPrimitives.scala 125:64:@22669.4]
  assign StickySelects_18_io_ins_3 = io_rPort_7_en_0 & _T_2857; // @[MemPrimitives.scala 125:64:@22670.4]
  assign StickySelects_18_io_ins_4 = io_rPort_8_en_0 & _T_2863; // @[MemPrimitives.scala 125:64:@22671.4]
  assign StickySelects_18_io_ins_5 = io_rPort_9_en_0 & _T_2869; // @[MemPrimitives.scala 125:64:@22672.4]
  assign StickySelects_18_io_ins_6 = io_rPort_11_en_0 & _T_2875; // @[MemPrimitives.scala 125:64:@22673.4]
  assign StickySelects_18_io_ins_7 = io_rPort_14_en_0 & _T_2881; // @[MemPrimitives.scala 125:64:@22674.4]
  assign StickySelects_18_io_ins_8 = io_rPort_16_en_0 & _T_2887; // @[MemPrimitives.scala 125:64:@22675.4]
  assign StickySelects_19_clock = clock; // @[:@22754.4]
  assign StickySelects_19_reset = reset; // @[:@22755.4]
  assign StickySelects_19_io_ins_0 = io_rPort_2_en_0 & _T_2931; // @[MemPrimitives.scala 125:64:@22756.4]
  assign StickySelects_19_io_ins_1 = io_rPort_3_en_0 & _T_2937; // @[MemPrimitives.scala 125:64:@22757.4]
  assign StickySelects_19_io_ins_2 = io_rPort_4_en_0 & _T_2943; // @[MemPrimitives.scala 125:64:@22758.4]
  assign StickySelects_19_io_ins_3 = io_rPort_6_en_0 & _T_2949; // @[MemPrimitives.scala 125:64:@22759.4]
  assign StickySelects_19_io_ins_4 = io_rPort_10_en_0 & _T_2955; // @[MemPrimitives.scala 125:64:@22760.4]
  assign StickySelects_19_io_ins_5 = io_rPort_12_en_0 & _T_2961; // @[MemPrimitives.scala 125:64:@22761.4]
  assign StickySelects_19_io_ins_6 = io_rPort_13_en_0 & _T_2967; // @[MemPrimitives.scala 125:64:@22762.4]
  assign StickySelects_19_io_ins_7 = io_rPort_15_en_0 & _T_2973; // @[MemPrimitives.scala 125:64:@22763.4]
  assign StickySelects_19_io_ins_8 = io_rPort_17_en_0 & _T_2979; // @[MemPrimitives.scala 125:64:@22764.4]
  assign StickySelects_20_clock = clock; // @[:@22843.4]
  assign StickySelects_20_reset = reset; // @[:@22844.4]
  assign StickySelects_20_io_ins_0 = io_rPort_0_en_0 & _T_3023; // @[MemPrimitives.scala 125:64:@22845.4]
  assign StickySelects_20_io_ins_1 = io_rPort_1_en_0 & _T_3029; // @[MemPrimitives.scala 125:64:@22846.4]
  assign StickySelects_20_io_ins_2 = io_rPort_5_en_0 & _T_3035; // @[MemPrimitives.scala 125:64:@22847.4]
  assign StickySelects_20_io_ins_3 = io_rPort_7_en_0 & _T_3041; // @[MemPrimitives.scala 125:64:@22848.4]
  assign StickySelects_20_io_ins_4 = io_rPort_8_en_0 & _T_3047; // @[MemPrimitives.scala 125:64:@22849.4]
  assign StickySelects_20_io_ins_5 = io_rPort_9_en_0 & _T_3053; // @[MemPrimitives.scala 125:64:@22850.4]
  assign StickySelects_20_io_ins_6 = io_rPort_11_en_0 & _T_3059; // @[MemPrimitives.scala 125:64:@22851.4]
  assign StickySelects_20_io_ins_7 = io_rPort_14_en_0 & _T_3065; // @[MemPrimitives.scala 125:64:@22852.4]
  assign StickySelects_20_io_ins_8 = io_rPort_16_en_0 & _T_3071; // @[MemPrimitives.scala 125:64:@22853.4]
  assign StickySelects_21_clock = clock; // @[:@22932.4]
  assign StickySelects_21_reset = reset; // @[:@22933.4]
  assign StickySelects_21_io_ins_0 = io_rPort_2_en_0 & _T_3115; // @[MemPrimitives.scala 125:64:@22934.4]
  assign StickySelects_21_io_ins_1 = io_rPort_3_en_0 & _T_3121; // @[MemPrimitives.scala 125:64:@22935.4]
  assign StickySelects_21_io_ins_2 = io_rPort_4_en_0 & _T_3127; // @[MemPrimitives.scala 125:64:@22936.4]
  assign StickySelects_21_io_ins_3 = io_rPort_6_en_0 & _T_3133; // @[MemPrimitives.scala 125:64:@22937.4]
  assign StickySelects_21_io_ins_4 = io_rPort_10_en_0 & _T_3139; // @[MemPrimitives.scala 125:64:@22938.4]
  assign StickySelects_21_io_ins_5 = io_rPort_12_en_0 & _T_3145; // @[MemPrimitives.scala 125:64:@22939.4]
  assign StickySelects_21_io_ins_6 = io_rPort_13_en_0 & _T_3151; // @[MemPrimitives.scala 125:64:@22940.4]
  assign StickySelects_21_io_ins_7 = io_rPort_15_en_0 & _T_3157; // @[MemPrimitives.scala 125:64:@22941.4]
  assign StickySelects_21_io_ins_8 = io_rPort_17_en_0 & _T_3163; // @[MemPrimitives.scala 125:64:@22942.4]
  assign StickySelects_22_clock = clock; // @[:@23021.4]
  assign StickySelects_22_reset = reset; // @[:@23022.4]
  assign StickySelects_22_io_ins_0 = io_rPort_0_en_0 & _T_3207; // @[MemPrimitives.scala 125:64:@23023.4]
  assign StickySelects_22_io_ins_1 = io_rPort_1_en_0 & _T_3213; // @[MemPrimitives.scala 125:64:@23024.4]
  assign StickySelects_22_io_ins_2 = io_rPort_5_en_0 & _T_3219; // @[MemPrimitives.scala 125:64:@23025.4]
  assign StickySelects_22_io_ins_3 = io_rPort_7_en_0 & _T_3225; // @[MemPrimitives.scala 125:64:@23026.4]
  assign StickySelects_22_io_ins_4 = io_rPort_8_en_0 & _T_3231; // @[MemPrimitives.scala 125:64:@23027.4]
  assign StickySelects_22_io_ins_5 = io_rPort_9_en_0 & _T_3237; // @[MemPrimitives.scala 125:64:@23028.4]
  assign StickySelects_22_io_ins_6 = io_rPort_11_en_0 & _T_3243; // @[MemPrimitives.scala 125:64:@23029.4]
  assign StickySelects_22_io_ins_7 = io_rPort_14_en_0 & _T_3249; // @[MemPrimitives.scala 125:64:@23030.4]
  assign StickySelects_22_io_ins_8 = io_rPort_16_en_0 & _T_3255; // @[MemPrimitives.scala 125:64:@23031.4]
  assign StickySelects_23_clock = clock; // @[:@23110.4]
  assign StickySelects_23_reset = reset; // @[:@23111.4]
  assign StickySelects_23_io_ins_0 = io_rPort_2_en_0 & _T_3299; // @[MemPrimitives.scala 125:64:@23112.4]
  assign StickySelects_23_io_ins_1 = io_rPort_3_en_0 & _T_3305; // @[MemPrimitives.scala 125:64:@23113.4]
  assign StickySelects_23_io_ins_2 = io_rPort_4_en_0 & _T_3311; // @[MemPrimitives.scala 125:64:@23114.4]
  assign StickySelects_23_io_ins_3 = io_rPort_6_en_0 & _T_3317; // @[MemPrimitives.scala 125:64:@23115.4]
  assign StickySelects_23_io_ins_4 = io_rPort_10_en_0 & _T_3323; // @[MemPrimitives.scala 125:64:@23116.4]
  assign StickySelects_23_io_ins_5 = io_rPort_12_en_0 & _T_3329; // @[MemPrimitives.scala 125:64:@23117.4]
  assign StickySelects_23_io_ins_6 = io_rPort_13_en_0 & _T_3335; // @[MemPrimitives.scala 125:64:@23118.4]
  assign StickySelects_23_io_ins_7 = io_rPort_15_en_0 & _T_3341; // @[MemPrimitives.scala 125:64:@23119.4]
  assign StickySelects_23_io_ins_8 = io_rPort_17_en_0 & _T_3347; // @[MemPrimitives.scala 125:64:@23120.4]
  assign RetimeWrapper_clock = clock; // @[:@23200.4]
  assign RetimeWrapper_reset = reset; // @[:@23201.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23203.4]
  assign RetimeWrapper_io_in = _T_1183 & io_rPort_0_en_0; // @[package.scala 94:16:@23202.4]
  assign RetimeWrapper_1_clock = clock; // @[:@23208.4]
  assign RetimeWrapper_1_reset = reset; // @[:@23209.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23211.4]
  assign RetimeWrapper_1_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@23210.4]
  assign RetimeWrapper_2_clock = clock; // @[:@23216.4]
  assign RetimeWrapper_2_reset = reset; // @[:@23217.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23219.4]
  assign RetimeWrapper_2_io_in = _T_1551 & io_rPort_0_en_0; // @[package.scala 94:16:@23218.4]
  assign RetimeWrapper_3_clock = clock; // @[:@23224.4]
  assign RetimeWrapper_3_reset = reset; // @[:@23225.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23227.4]
  assign RetimeWrapper_3_io_in = _T_1735 & io_rPort_0_en_0; // @[package.scala 94:16:@23226.4]
  assign RetimeWrapper_4_clock = clock; // @[:@23232.4]
  assign RetimeWrapper_4_reset = reset; // @[:@23233.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23235.4]
  assign RetimeWrapper_4_io_in = _T_1919 & io_rPort_0_en_0; // @[package.scala 94:16:@23234.4]
  assign RetimeWrapper_5_clock = clock; // @[:@23240.4]
  assign RetimeWrapper_5_reset = reset; // @[:@23241.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23243.4]
  assign RetimeWrapper_5_io_in = _T_2103 & io_rPort_0_en_0; // @[package.scala 94:16:@23242.4]
  assign RetimeWrapper_6_clock = clock; // @[:@23248.4]
  assign RetimeWrapper_6_reset = reset; // @[:@23249.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23251.4]
  assign RetimeWrapper_6_io_in = _T_2287 & io_rPort_0_en_0; // @[package.scala 94:16:@23250.4]
  assign RetimeWrapper_7_clock = clock; // @[:@23256.4]
  assign RetimeWrapper_7_reset = reset; // @[:@23257.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23259.4]
  assign RetimeWrapper_7_io_in = _T_2471 & io_rPort_0_en_0; // @[package.scala 94:16:@23258.4]
  assign RetimeWrapper_8_clock = clock; // @[:@23264.4]
  assign RetimeWrapper_8_reset = reset; // @[:@23265.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23267.4]
  assign RetimeWrapper_8_io_in = _T_2655 & io_rPort_0_en_0; // @[package.scala 94:16:@23266.4]
  assign RetimeWrapper_9_clock = clock; // @[:@23272.4]
  assign RetimeWrapper_9_reset = reset; // @[:@23273.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23275.4]
  assign RetimeWrapper_9_io_in = _T_2839 & io_rPort_0_en_0; // @[package.scala 94:16:@23274.4]
  assign RetimeWrapper_10_clock = clock; // @[:@23280.4]
  assign RetimeWrapper_10_reset = reset; // @[:@23281.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23283.4]
  assign RetimeWrapper_10_io_in = _T_3023 & io_rPort_0_en_0; // @[package.scala 94:16:@23282.4]
  assign RetimeWrapper_11_clock = clock; // @[:@23288.4]
  assign RetimeWrapper_11_reset = reset; // @[:@23289.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23291.4]
  assign RetimeWrapper_11_io_in = _T_3207 & io_rPort_0_en_0; // @[package.scala 94:16:@23290.4]
  assign RetimeWrapper_12_clock = clock; // @[:@23344.4]
  assign RetimeWrapper_12_reset = reset; // @[:@23345.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23347.4]
  assign RetimeWrapper_12_io_in = _T_1189 & io_rPort_1_en_0; // @[package.scala 94:16:@23346.4]
  assign RetimeWrapper_13_clock = clock; // @[:@23352.4]
  assign RetimeWrapper_13_reset = reset; // @[:@23353.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23355.4]
  assign RetimeWrapper_13_io_in = _T_1373 & io_rPort_1_en_0; // @[package.scala 94:16:@23354.4]
  assign RetimeWrapper_14_clock = clock; // @[:@23360.4]
  assign RetimeWrapper_14_reset = reset; // @[:@23361.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23363.4]
  assign RetimeWrapper_14_io_in = _T_1557 & io_rPort_1_en_0; // @[package.scala 94:16:@23362.4]
  assign RetimeWrapper_15_clock = clock; // @[:@23368.4]
  assign RetimeWrapper_15_reset = reset; // @[:@23369.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23371.4]
  assign RetimeWrapper_15_io_in = _T_1741 & io_rPort_1_en_0; // @[package.scala 94:16:@23370.4]
  assign RetimeWrapper_16_clock = clock; // @[:@23376.4]
  assign RetimeWrapper_16_reset = reset; // @[:@23377.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23379.4]
  assign RetimeWrapper_16_io_in = _T_1925 & io_rPort_1_en_0; // @[package.scala 94:16:@23378.4]
  assign RetimeWrapper_17_clock = clock; // @[:@23384.4]
  assign RetimeWrapper_17_reset = reset; // @[:@23385.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23387.4]
  assign RetimeWrapper_17_io_in = _T_2109 & io_rPort_1_en_0; // @[package.scala 94:16:@23386.4]
  assign RetimeWrapper_18_clock = clock; // @[:@23392.4]
  assign RetimeWrapper_18_reset = reset; // @[:@23393.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23395.4]
  assign RetimeWrapper_18_io_in = _T_2293 & io_rPort_1_en_0; // @[package.scala 94:16:@23394.4]
  assign RetimeWrapper_19_clock = clock; // @[:@23400.4]
  assign RetimeWrapper_19_reset = reset; // @[:@23401.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23403.4]
  assign RetimeWrapper_19_io_in = _T_2477 & io_rPort_1_en_0; // @[package.scala 94:16:@23402.4]
  assign RetimeWrapper_20_clock = clock; // @[:@23408.4]
  assign RetimeWrapper_20_reset = reset; // @[:@23409.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23411.4]
  assign RetimeWrapper_20_io_in = _T_2661 & io_rPort_1_en_0; // @[package.scala 94:16:@23410.4]
  assign RetimeWrapper_21_clock = clock; // @[:@23416.4]
  assign RetimeWrapper_21_reset = reset; // @[:@23417.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23419.4]
  assign RetimeWrapper_21_io_in = _T_2845 & io_rPort_1_en_0; // @[package.scala 94:16:@23418.4]
  assign RetimeWrapper_22_clock = clock; // @[:@23424.4]
  assign RetimeWrapper_22_reset = reset; // @[:@23425.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23427.4]
  assign RetimeWrapper_22_io_in = _T_3029 & io_rPort_1_en_0; // @[package.scala 94:16:@23426.4]
  assign RetimeWrapper_23_clock = clock; // @[:@23432.4]
  assign RetimeWrapper_23_reset = reset; // @[:@23433.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23435.4]
  assign RetimeWrapper_23_io_in = _T_3213 & io_rPort_1_en_0; // @[package.scala 94:16:@23434.4]
  assign RetimeWrapper_24_clock = clock; // @[:@23488.4]
  assign RetimeWrapper_24_reset = reset; // @[:@23489.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23491.4]
  assign RetimeWrapper_24_io_in = _T_1275 & io_rPort_2_en_0; // @[package.scala 94:16:@23490.4]
  assign RetimeWrapper_25_clock = clock; // @[:@23496.4]
  assign RetimeWrapper_25_reset = reset; // @[:@23497.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23499.4]
  assign RetimeWrapper_25_io_in = _T_1459 & io_rPort_2_en_0; // @[package.scala 94:16:@23498.4]
  assign RetimeWrapper_26_clock = clock; // @[:@23504.4]
  assign RetimeWrapper_26_reset = reset; // @[:@23505.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23507.4]
  assign RetimeWrapper_26_io_in = _T_1643 & io_rPort_2_en_0; // @[package.scala 94:16:@23506.4]
  assign RetimeWrapper_27_clock = clock; // @[:@23512.4]
  assign RetimeWrapper_27_reset = reset; // @[:@23513.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23515.4]
  assign RetimeWrapper_27_io_in = _T_1827 & io_rPort_2_en_0; // @[package.scala 94:16:@23514.4]
  assign RetimeWrapper_28_clock = clock; // @[:@23520.4]
  assign RetimeWrapper_28_reset = reset; // @[:@23521.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23523.4]
  assign RetimeWrapper_28_io_in = _T_2011 & io_rPort_2_en_0; // @[package.scala 94:16:@23522.4]
  assign RetimeWrapper_29_clock = clock; // @[:@23528.4]
  assign RetimeWrapper_29_reset = reset; // @[:@23529.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23531.4]
  assign RetimeWrapper_29_io_in = _T_2195 & io_rPort_2_en_0; // @[package.scala 94:16:@23530.4]
  assign RetimeWrapper_30_clock = clock; // @[:@23536.4]
  assign RetimeWrapper_30_reset = reset; // @[:@23537.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23539.4]
  assign RetimeWrapper_30_io_in = _T_2379 & io_rPort_2_en_0; // @[package.scala 94:16:@23538.4]
  assign RetimeWrapper_31_clock = clock; // @[:@23544.4]
  assign RetimeWrapper_31_reset = reset; // @[:@23545.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23547.4]
  assign RetimeWrapper_31_io_in = _T_2563 & io_rPort_2_en_0; // @[package.scala 94:16:@23546.4]
  assign RetimeWrapper_32_clock = clock; // @[:@23552.4]
  assign RetimeWrapper_32_reset = reset; // @[:@23553.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23555.4]
  assign RetimeWrapper_32_io_in = _T_2747 & io_rPort_2_en_0; // @[package.scala 94:16:@23554.4]
  assign RetimeWrapper_33_clock = clock; // @[:@23560.4]
  assign RetimeWrapper_33_reset = reset; // @[:@23561.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23563.4]
  assign RetimeWrapper_33_io_in = _T_2931 & io_rPort_2_en_0; // @[package.scala 94:16:@23562.4]
  assign RetimeWrapper_34_clock = clock; // @[:@23568.4]
  assign RetimeWrapper_34_reset = reset; // @[:@23569.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23571.4]
  assign RetimeWrapper_34_io_in = _T_3115 & io_rPort_2_en_0; // @[package.scala 94:16:@23570.4]
  assign RetimeWrapper_35_clock = clock; // @[:@23576.4]
  assign RetimeWrapper_35_reset = reset; // @[:@23577.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23579.4]
  assign RetimeWrapper_35_io_in = _T_3299 & io_rPort_2_en_0; // @[package.scala 94:16:@23578.4]
  assign RetimeWrapper_36_clock = clock; // @[:@23632.4]
  assign RetimeWrapper_36_reset = reset; // @[:@23633.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23635.4]
  assign RetimeWrapper_36_io_in = _T_1281 & io_rPort_3_en_0; // @[package.scala 94:16:@23634.4]
  assign RetimeWrapper_37_clock = clock; // @[:@23640.4]
  assign RetimeWrapper_37_reset = reset; // @[:@23641.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23643.4]
  assign RetimeWrapper_37_io_in = _T_1465 & io_rPort_3_en_0; // @[package.scala 94:16:@23642.4]
  assign RetimeWrapper_38_clock = clock; // @[:@23648.4]
  assign RetimeWrapper_38_reset = reset; // @[:@23649.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23651.4]
  assign RetimeWrapper_38_io_in = _T_1649 & io_rPort_3_en_0; // @[package.scala 94:16:@23650.4]
  assign RetimeWrapper_39_clock = clock; // @[:@23656.4]
  assign RetimeWrapper_39_reset = reset; // @[:@23657.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23659.4]
  assign RetimeWrapper_39_io_in = _T_1833 & io_rPort_3_en_0; // @[package.scala 94:16:@23658.4]
  assign RetimeWrapper_40_clock = clock; // @[:@23664.4]
  assign RetimeWrapper_40_reset = reset; // @[:@23665.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23667.4]
  assign RetimeWrapper_40_io_in = _T_2017 & io_rPort_3_en_0; // @[package.scala 94:16:@23666.4]
  assign RetimeWrapper_41_clock = clock; // @[:@23672.4]
  assign RetimeWrapper_41_reset = reset; // @[:@23673.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23675.4]
  assign RetimeWrapper_41_io_in = _T_2201 & io_rPort_3_en_0; // @[package.scala 94:16:@23674.4]
  assign RetimeWrapper_42_clock = clock; // @[:@23680.4]
  assign RetimeWrapper_42_reset = reset; // @[:@23681.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23683.4]
  assign RetimeWrapper_42_io_in = _T_2385 & io_rPort_3_en_0; // @[package.scala 94:16:@23682.4]
  assign RetimeWrapper_43_clock = clock; // @[:@23688.4]
  assign RetimeWrapper_43_reset = reset; // @[:@23689.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23691.4]
  assign RetimeWrapper_43_io_in = _T_2569 & io_rPort_3_en_0; // @[package.scala 94:16:@23690.4]
  assign RetimeWrapper_44_clock = clock; // @[:@23696.4]
  assign RetimeWrapper_44_reset = reset; // @[:@23697.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23699.4]
  assign RetimeWrapper_44_io_in = _T_2753 & io_rPort_3_en_0; // @[package.scala 94:16:@23698.4]
  assign RetimeWrapper_45_clock = clock; // @[:@23704.4]
  assign RetimeWrapper_45_reset = reset; // @[:@23705.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23707.4]
  assign RetimeWrapper_45_io_in = _T_2937 & io_rPort_3_en_0; // @[package.scala 94:16:@23706.4]
  assign RetimeWrapper_46_clock = clock; // @[:@23712.4]
  assign RetimeWrapper_46_reset = reset; // @[:@23713.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23715.4]
  assign RetimeWrapper_46_io_in = _T_3121 & io_rPort_3_en_0; // @[package.scala 94:16:@23714.4]
  assign RetimeWrapper_47_clock = clock; // @[:@23720.4]
  assign RetimeWrapper_47_reset = reset; // @[:@23721.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23723.4]
  assign RetimeWrapper_47_io_in = _T_3305 & io_rPort_3_en_0; // @[package.scala 94:16:@23722.4]
  assign RetimeWrapper_48_clock = clock; // @[:@23776.4]
  assign RetimeWrapper_48_reset = reset; // @[:@23777.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23779.4]
  assign RetimeWrapper_48_io_in = _T_1287 & io_rPort_4_en_0; // @[package.scala 94:16:@23778.4]
  assign RetimeWrapper_49_clock = clock; // @[:@23784.4]
  assign RetimeWrapper_49_reset = reset; // @[:@23785.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23787.4]
  assign RetimeWrapper_49_io_in = _T_1471 & io_rPort_4_en_0; // @[package.scala 94:16:@23786.4]
  assign RetimeWrapper_50_clock = clock; // @[:@23792.4]
  assign RetimeWrapper_50_reset = reset; // @[:@23793.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23795.4]
  assign RetimeWrapper_50_io_in = _T_1655 & io_rPort_4_en_0; // @[package.scala 94:16:@23794.4]
  assign RetimeWrapper_51_clock = clock; // @[:@23800.4]
  assign RetimeWrapper_51_reset = reset; // @[:@23801.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23803.4]
  assign RetimeWrapper_51_io_in = _T_1839 & io_rPort_4_en_0; // @[package.scala 94:16:@23802.4]
  assign RetimeWrapper_52_clock = clock; // @[:@23808.4]
  assign RetimeWrapper_52_reset = reset; // @[:@23809.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23811.4]
  assign RetimeWrapper_52_io_in = _T_2023 & io_rPort_4_en_0; // @[package.scala 94:16:@23810.4]
  assign RetimeWrapper_53_clock = clock; // @[:@23816.4]
  assign RetimeWrapper_53_reset = reset; // @[:@23817.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23819.4]
  assign RetimeWrapper_53_io_in = _T_2207 & io_rPort_4_en_0; // @[package.scala 94:16:@23818.4]
  assign RetimeWrapper_54_clock = clock; // @[:@23824.4]
  assign RetimeWrapper_54_reset = reset; // @[:@23825.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23827.4]
  assign RetimeWrapper_54_io_in = _T_2391 & io_rPort_4_en_0; // @[package.scala 94:16:@23826.4]
  assign RetimeWrapper_55_clock = clock; // @[:@23832.4]
  assign RetimeWrapper_55_reset = reset; // @[:@23833.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23835.4]
  assign RetimeWrapper_55_io_in = _T_2575 & io_rPort_4_en_0; // @[package.scala 94:16:@23834.4]
  assign RetimeWrapper_56_clock = clock; // @[:@23840.4]
  assign RetimeWrapper_56_reset = reset; // @[:@23841.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23843.4]
  assign RetimeWrapper_56_io_in = _T_2759 & io_rPort_4_en_0; // @[package.scala 94:16:@23842.4]
  assign RetimeWrapper_57_clock = clock; // @[:@23848.4]
  assign RetimeWrapper_57_reset = reset; // @[:@23849.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23851.4]
  assign RetimeWrapper_57_io_in = _T_2943 & io_rPort_4_en_0; // @[package.scala 94:16:@23850.4]
  assign RetimeWrapper_58_clock = clock; // @[:@23856.4]
  assign RetimeWrapper_58_reset = reset; // @[:@23857.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23859.4]
  assign RetimeWrapper_58_io_in = _T_3127 & io_rPort_4_en_0; // @[package.scala 94:16:@23858.4]
  assign RetimeWrapper_59_clock = clock; // @[:@23864.4]
  assign RetimeWrapper_59_reset = reset; // @[:@23865.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23867.4]
  assign RetimeWrapper_59_io_in = _T_3311 & io_rPort_4_en_0; // @[package.scala 94:16:@23866.4]
  assign RetimeWrapper_60_clock = clock; // @[:@23920.4]
  assign RetimeWrapper_60_reset = reset; // @[:@23921.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23923.4]
  assign RetimeWrapper_60_io_in = _T_1195 & io_rPort_5_en_0; // @[package.scala 94:16:@23922.4]
  assign RetimeWrapper_61_clock = clock; // @[:@23928.4]
  assign RetimeWrapper_61_reset = reset; // @[:@23929.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23931.4]
  assign RetimeWrapper_61_io_in = _T_1379 & io_rPort_5_en_0; // @[package.scala 94:16:@23930.4]
  assign RetimeWrapper_62_clock = clock; // @[:@23936.4]
  assign RetimeWrapper_62_reset = reset; // @[:@23937.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23939.4]
  assign RetimeWrapper_62_io_in = _T_1563 & io_rPort_5_en_0; // @[package.scala 94:16:@23938.4]
  assign RetimeWrapper_63_clock = clock; // @[:@23944.4]
  assign RetimeWrapper_63_reset = reset; // @[:@23945.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23947.4]
  assign RetimeWrapper_63_io_in = _T_1747 & io_rPort_5_en_0; // @[package.scala 94:16:@23946.4]
  assign RetimeWrapper_64_clock = clock; // @[:@23952.4]
  assign RetimeWrapper_64_reset = reset; // @[:@23953.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23955.4]
  assign RetimeWrapper_64_io_in = _T_1931 & io_rPort_5_en_0; // @[package.scala 94:16:@23954.4]
  assign RetimeWrapper_65_clock = clock; // @[:@23960.4]
  assign RetimeWrapper_65_reset = reset; // @[:@23961.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23963.4]
  assign RetimeWrapper_65_io_in = _T_2115 & io_rPort_5_en_0; // @[package.scala 94:16:@23962.4]
  assign RetimeWrapper_66_clock = clock; // @[:@23968.4]
  assign RetimeWrapper_66_reset = reset; // @[:@23969.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23971.4]
  assign RetimeWrapper_66_io_in = _T_2299 & io_rPort_5_en_0; // @[package.scala 94:16:@23970.4]
  assign RetimeWrapper_67_clock = clock; // @[:@23976.4]
  assign RetimeWrapper_67_reset = reset; // @[:@23977.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23979.4]
  assign RetimeWrapper_67_io_in = _T_2483 & io_rPort_5_en_0; // @[package.scala 94:16:@23978.4]
  assign RetimeWrapper_68_clock = clock; // @[:@23984.4]
  assign RetimeWrapper_68_reset = reset; // @[:@23985.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23987.4]
  assign RetimeWrapper_68_io_in = _T_2667 & io_rPort_5_en_0; // @[package.scala 94:16:@23986.4]
  assign RetimeWrapper_69_clock = clock; // @[:@23992.4]
  assign RetimeWrapper_69_reset = reset; // @[:@23993.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23995.4]
  assign RetimeWrapper_69_io_in = _T_2851 & io_rPort_5_en_0; // @[package.scala 94:16:@23994.4]
  assign RetimeWrapper_70_clock = clock; // @[:@24000.4]
  assign RetimeWrapper_70_reset = reset; // @[:@24001.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@24003.4]
  assign RetimeWrapper_70_io_in = _T_3035 & io_rPort_5_en_0; // @[package.scala 94:16:@24002.4]
  assign RetimeWrapper_71_clock = clock; // @[:@24008.4]
  assign RetimeWrapper_71_reset = reset; // @[:@24009.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@24011.4]
  assign RetimeWrapper_71_io_in = _T_3219 & io_rPort_5_en_0; // @[package.scala 94:16:@24010.4]
  assign RetimeWrapper_72_clock = clock; // @[:@24064.4]
  assign RetimeWrapper_72_reset = reset; // @[:@24065.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24067.4]
  assign RetimeWrapper_72_io_in = _T_1293 & io_rPort_6_en_0; // @[package.scala 94:16:@24066.4]
  assign RetimeWrapper_73_clock = clock; // @[:@24072.4]
  assign RetimeWrapper_73_reset = reset; // @[:@24073.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24075.4]
  assign RetimeWrapper_73_io_in = _T_1477 & io_rPort_6_en_0; // @[package.scala 94:16:@24074.4]
  assign RetimeWrapper_74_clock = clock; // @[:@24080.4]
  assign RetimeWrapper_74_reset = reset; // @[:@24081.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24083.4]
  assign RetimeWrapper_74_io_in = _T_1661 & io_rPort_6_en_0; // @[package.scala 94:16:@24082.4]
  assign RetimeWrapper_75_clock = clock; // @[:@24088.4]
  assign RetimeWrapper_75_reset = reset; // @[:@24089.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24091.4]
  assign RetimeWrapper_75_io_in = _T_1845 & io_rPort_6_en_0; // @[package.scala 94:16:@24090.4]
  assign RetimeWrapper_76_clock = clock; // @[:@24096.4]
  assign RetimeWrapper_76_reset = reset; // @[:@24097.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24099.4]
  assign RetimeWrapper_76_io_in = _T_2029 & io_rPort_6_en_0; // @[package.scala 94:16:@24098.4]
  assign RetimeWrapper_77_clock = clock; // @[:@24104.4]
  assign RetimeWrapper_77_reset = reset; // @[:@24105.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24107.4]
  assign RetimeWrapper_77_io_in = _T_2213 & io_rPort_6_en_0; // @[package.scala 94:16:@24106.4]
  assign RetimeWrapper_78_clock = clock; // @[:@24112.4]
  assign RetimeWrapper_78_reset = reset; // @[:@24113.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24115.4]
  assign RetimeWrapper_78_io_in = _T_2397 & io_rPort_6_en_0; // @[package.scala 94:16:@24114.4]
  assign RetimeWrapper_79_clock = clock; // @[:@24120.4]
  assign RetimeWrapper_79_reset = reset; // @[:@24121.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24123.4]
  assign RetimeWrapper_79_io_in = _T_2581 & io_rPort_6_en_0; // @[package.scala 94:16:@24122.4]
  assign RetimeWrapper_80_clock = clock; // @[:@24128.4]
  assign RetimeWrapper_80_reset = reset; // @[:@24129.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24131.4]
  assign RetimeWrapper_80_io_in = _T_2765 & io_rPort_6_en_0; // @[package.scala 94:16:@24130.4]
  assign RetimeWrapper_81_clock = clock; // @[:@24136.4]
  assign RetimeWrapper_81_reset = reset; // @[:@24137.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24139.4]
  assign RetimeWrapper_81_io_in = _T_2949 & io_rPort_6_en_0; // @[package.scala 94:16:@24138.4]
  assign RetimeWrapper_82_clock = clock; // @[:@24144.4]
  assign RetimeWrapper_82_reset = reset; // @[:@24145.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24147.4]
  assign RetimeWrapper_82_io_in = _T_3133 & io_rPort_6_en_0; // @[package.scala 94:16:@24146.4]
  assign RetimeWrapper_83_clock = clock; // @[:@24152.4]
  assign RetimeWrapper_83_reset = reset; // @[:@24153.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24155.4]
  assign RetimeWrapper_83_io_in = _T_3317 & io_rPort_6_en_0; // @[package.scala 94:16:@24154.4]
  assign RetimeWrapper_84_clock = clock; // @[:@24208.4]
  assign RetimeWrapper_84_reset = reset; // @[:@24209.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24211.4]
  assign RetimeWrapper_84_io_in = _T_1201 & io_rPort_7_en_0; // @[package.scala 94:16:@24210.4]
  assign RetimeWrapper_85_clock = clock; // @[:@24216.4]
  assign RetimeWrapper_85_reset = reset; // @[:@24217.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24219.4]
  assign RetimeWrapper_85_io_in = _T_1385 & io_rPort_7_en_0; // @[package.scala 94:16:@24218.4]
  assign RetimeWrapper_86_clock = clock; // @[:@24224.4]
  assign RetimeWrapper_86_reset = reset; // @[:@24225.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24227.4]
  assign RetimeWrapper_86_io_in = _T_1569 & io_rPort_7_en_0; // @[package.scala 94:16:@24226.4]
  assign RetimeWrapper_87_clock = clock; // @[:@24232.4]
  assign RetimeWrapper_87_reset = reset; // @[:@24233.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24235.4]
  assign RetimeWrapper_87_io_in = _T_1753 & io_rPort_7_en_0; // @[package.scala 94:16:@24234.4]
  assign RetimeWrapper_88_clock = clock; // @[:@24240.4]
  assign RetimeWrapper_88_reset = reset; // @[:@24241.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24243.4]
  assign RetimeWrapper_88_io_in = _T_1937 & io_rPort_7_en_0; // @[package.scala 94:16:@24242.4]
  assign RetimeWrapper_89_clock = clock; // @[:@24248.4]
  assign RetimeWrapper_89_reset = reset; // @[:@24249.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24251.4]
  assign RetimeWrapper_89_io_in = _T_2121 & io_rPort_7_en_0; // @[package.scala 94:16:@24250.4]
  assign RetimeWrapper_90_clock = clock; // @[:@24256.4]
  assign RetimeWrapper_90_reset = reset; // @[:@24257.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24259.4]
  assign RetimeWrapper_90_io_in = _T_2305 & io_rPort_7_en_0; // @[package.scala 94:16:@24258.4]
  assign RetimeWrapper_91_clock = clock; // @[:@24264.4]
  assign RetimeWrapper_91_reset = reset; // @[:@24265.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24267.4]
  assign RetimeWrapper_91_io_in = _T_2489 & io_rPort_7_en_0; // @[package.scala 94:16:@24266.4]
  assign RetimeWrapper_92_clock = clock; // @[:@24272.4]
  assign RetimeWrapper_92_reset = reset; // @[:@24273.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24275.4]
  assign RetimeWrapper_92_io_in = _T_2673 & io_rPort_7_en_0; // @[package.scala 94:16:@24274.4]
  assign RetimeWrapper_93_clock = clock; // @[:@24280.4]
  assign RetimeWrapper_93_reset = reset; // @[:@24281.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24283.4]
  assign RetimeWrapper_93_io_in = _T_2857 & io_rPort_7_en_0; // @[package.scala 94:16:@24282.4]
  assign RetimeWrapper_94_clock = clock; // @[:@24288.4]
  assign RetimeWrapper_94_reset = reset; // @[:@24289.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24291.4]
  assign RetimeWrapper_94_io_in = _T_3041 & io_rPort_7_en_0; // @[package.scala 94:16:@24290.4]
  assign RetimeWrapper_95_clock = clock; // @[:@24296.4]
  assign RetimeWrapper_95_reset = reset; // @[:@24297.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24299.4]
  assign RetimeWrapper_95_io_in = _T_3225 & io_rPort_7_en_0; // @[package.scala 94:16:@24298.4]
  assign RetimeWrapper_96_clock = clock; // @[:@24352.4]
  assign RetimeWrapper_96_reset = reset; // @[:@24353.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24355.4]
  assign RetimeWrapper_96_io_in = _T_1207 & io_rPort_8_en_0; // @[package.scala 94:16:@24354.4]
  assign RetimeWrapper_97_clock = clock; // @[:@24360.4]
  assign RetimeWrapper_97_reset = reset; // @[:@24361.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24363.4]
  assign RetimeWrapper_97_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@24362.4]
  assign RetimeWrapper_98_clock = clock; // @[:@24368.4]
  assign RetimeWrapper_98_reset = reset; // @[:@24369.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24371.4]
  assign RetimeWrapper_98_io_in = _T_1575 & io_rPort_8_en_0; // @[package.scala 94:16:@24370.4]
  assign RetimeWrapper_99_clock = clock; // @[:@24376.4]
  assign RetimeWrapper_99_reset = reset; // @[:@24377.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24379.4]
  assign RetimeWrapper_99_io_in = _T_1759 & io_rPort_8_en_0; // @[package.scala 94:16:@24378.4]
  assign RetimeWrapper_100_clock = clock; // @[:@24384.4]
  assign RetimeWrapper_100_reset = reset; // @[:@24385.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24387.4]
  assign RetimeWrapper_100_io_in = _T_1943 & io_rPort_8_en_0; // @[package.scala 94:16:@24386.4]
  assign RetimeWrapper_101_clock = clock; // @[:@24392.4]
  assign RetimeWrapper_101_reset = reset; // @[:@24393.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24395.4]
  assign RetimeWrapper_101_io_in = _T_2127 & io_rPort_8_en_0; // @[package.scala 94:16:@24394.4]
  assign RetimeWrapper_102_clock = clock; // @[:@24400.4]
  assign RetimeWrapper_102_reset = reset; // @[:@24401.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24403.4]
  assign RetimeWrapper_102_io_in = _T_2311 & io_rPort_8_en_0; // @[package.scala 94:16:@24402.4]
  assign RetimeWrapper_103_clock = clock; // @[:@24408.4]
  assign RetimeWrapper_103_reset = reset; // @[:@24409.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24411.4]
  assign RetimeWrapper_103_io_in = _T_2495 & io_rPort_8_en_0; // @[package.scala 94:16:@24410.4]
  assign RetimeWrapper_104_clock = clock; // @[:@24416.4]
  assign RetimeWrapper_104_reset = reset; // @[:@24417.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24419.4]
  assign RetimeWrapper_104_io_in = _T_2679 & io_rPort_8_en_0; // @[package.scala 94:16:@24418.4]
  assign RetimeWrapper_105_clock = clock; // @[:@24424.4]
  assign RetimeWrapper_105_reset = reset; // @[:@24425.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24427.4]
  assign RetimeWrapper_105_io_in = _T_2863 & io_rPort_8_en_0; // @[package.scala 94:16:@24426.4]
  assign RetimeWrapper_106_clock = clock; // @[:@24432.4]
  assign RetimeWrapper_106_reset = reset; // @[:@24433.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24435.4]
  assign RetimeWrapper_106_io_in = _T_3047 & io_rPort_8_en_0; // @[package.scala 94:16:@24434.4]
  assign RetimeWrapper_107_clock = clock; // @[:@24440.4]
  assign RetimeWrapper_107_reset = reset; // @[:@24441.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24443.4]
  assign RetimeWrapper_107_io_in = _T_3231 & io_rPort_8_en_0; // @[package.scala 94:16:@24442.4]
  assign RetimeWrapper_108_clock = clock; // @[:@24496.4]
  assign RetimeWrapper_108_reset = reset; // @[:@24497.4]
  assign RetimeWrapper_108_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24499.4]
  assign RetimeWrapper_108_io_in = _T_1213 & io_rPort_9_en_0; // @[package.scala 94:16:@24498.4]
  assign RetimeWrapper_109_clock = clock; // @[:@24504.4]
  assign RetimeWrapper_109_reset = reset; // @[:@24505.4]
  assign RetimeWrapper_109_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24507.4]
  assign RetimeWrapper_109_io_in = _T_1397 & io_rPort_9_en_0; // @[package.scala 94:16:@24506.4]
  assign RetimeWrapper_110_clock = clock; // @[:@24512.4]
  assign RetimeWrapper_110_reset = reset; // @[:@24513.4]
  assign RetimeWrapper_110_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24515.4]
  assign RetimeWrapper_110_io_in = _T_1581 & io_rPort_9_en_0; // @[package.scala 94:16:@24514.4]
  assign RetimeWrapper_111_clock = clock; // @[:@24520.4]
  assign RetimeWrapper_111_reset = reset; // @[:@24521.4]
  assign RetimeWrapper_111_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24523.4]
  assign RetimeWrapper_111_io_in = _T_1765 & io_rPort_9_en_0; // @[package.scala 94:16:@24522.4]
  assign RetimeWrapper_112_clock = clock; // @[:@24528.4]
  assign RetimeWrapper_112_reset = reset; // @[:@24529.4]
  assign RetimeWrapper_112_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24531.4]
  assign RetimeWrapper_112_io_in = _T_1949 & io_rPort_9_en_0; // @[package.scala 94:16:@24530.4]
  assign RetimeWrapper_113_clock = clock; // @[:@24536.4]
  assign RetimeWrapper_113_reset = reset; // @[:@24537.4]
  assign RetimeWrapper_113_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24539.4]
  assign RetimeWrapper_113_io_in = _T_2133 & io_rPort_9_en_0; // @[package.scala 94:16:@24538.4]
  assign RetimeWrapper_114_clock = clock; // @[:@24544.4]
  assign RetimeWrapper_114_reset = reset; // @[:@24545.4]
  assign RetimeWrapper_114_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24547.4]
  assign RetimeWrapper_114_io_in = _T_2317 & io_rPort_9_en_0; // @[package.scala 94:16:@24546.4]
  assign RetimeWrapper_115_clock = clock; // @[:@24552.4]
  assign RetimeWrapper_115_reset = reset; // @[:@24553.4]
  assign RetimeWrapper_115_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24555.4]
  assign RetimeWrapper_115_io_in = _T_2501 & io_rPort_9_en_0; // @[package.scala 94:16:@24554.4]
  assign RetimeWrapper_116_clock = clock; // @[:@24560.4]
  assign RetimeWrapper_116_reset = reset; // @[:@24561.4]
  assign RetimeWrapper_116_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24563.4]
  assign RetimeWrapper_116_io_in = _T_2685 & io_rPort_9_en_0; // @[package.scala 94:16:@24562.4]
  assign RetimeWrapper_117_clock = clock; // @[:@24568.4]
  assign RetimeWrapper_117_reset = reset; // @[:@24569.4]
  assign RetimeWrapper_117_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24571.4]
  assign RetimeWrapper_117_io_in = _T_2869 & io_rPort_9_en_0; // @[package.scala 94:16:@24570.4]
  assign RetimeWrapper_118_clock = clock; // @[:@24576.4]
  assign RetimeWrapper_118_reset = reset; // @[:@24577.4]
  assign RetimeWrapper_118_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24579.4]
  assign RetimeWrapper_118_io_in = _T_3053 & io_rPort_9_en_0; // @[package.scala 94:16:@24578.4]
  assign RetimeWrapper_119_clock = clock; // @[:@24584.4]
  assign RetimeWrapper_119_reset = reset; // @[:@24585.4]
  assign RetimeWrapper_119_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24587.4]
  assign RetimeWrapper_119_io_in = _T_3237 & io_rPort_9_en_0; // @[package.scala 94:16:@24586.4]
  assign RetimeWrapper_120_clock = clock; // @[:@24640.4]
  assign RetimeWrapper_120_reset = reset; // @[:@24641.4]
  assign RetimeWrapper_120_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24643.4]
  assign RetimeWrapper_120_io_in = _T_1299 & io_rPort_10_en_0; // @[package.scala 94:16:@24642.4]
  assign RetimeWrapper_121_clock = clock; // @[:@24648.4]
  assign RetimeWrapper_121_reset = reset; // @[:@24649.4]
  assign RetimeWrapper_121_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24651.4]
  assign RetimeWrapper_121_io_in = _T_1483 & io_rPort_10_en_0; // @[package.scala 94:16:@24650.4]
  assign RetimeWrapper_122_clock = clock; // @[:@24656.4]
  assign RetimeWrapper_122_reset = reset; // @[:@24657.4]
  assign RetimeWrapper_122_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24659.4]
  assign RetimeWrapper_122_io_in = _T_1667 & io_rPort_10_en_0; // @[package.scala 94:16:@24658.4]
  assign RetimeWrapper_123_clock = clock; // @[:@24664.4]
  assign RetimeWrapper_123_reset = reset; // @[:@24665.4]
  assign RetimeWrapper_123_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24667.4]
  assign RetimeWrapper_123_io_in = _T_1851 & io_rPort_10_en_0; // @[package.scala 94:16:@24666.4]
  assign RetimeWrapper_124_clock = clock; // @[:@24672.4]
  assign RetimeWrapper_124_reset = reset; // @[:@24673.4]
  assign RetimeWrapper_124_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24675.4]
  assign RetimeWrapper_124_io_in = _T_2035 & io_rPort_10_en_0; // @[package.scala 94:16:@24674.4]
  assign RetimeWrapper_125_clock = clock; // @[:@24680.4]
  assign RetimeWrapper_125_reset = reset; // @[:@24681.4]
  assign RetimeWrapper_125_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24683.4]
  assign RetimeWrapper_125_io_in = _T_2219 & io_rPort_10_en_0; // @[package.scala 94:16:@24682.4]
  assign RetimeWrapper_126_clock = clock; // @[:@24688.4]
  assign RetimeWrapper_126_reset = reset; // @[:@24689.4]
  assign RetimeWrapper_126_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24691.4]
  assign RetimeWrapper_126_io_in = _T_2403 & io_rPort_10_en_0; // @[package.scala 94:16:@24690.4]
  assign RetimeWrapper_127_clock = clock; // @[:@24696.4]
  assign RetimeWrapper_127_reset = reset; // @[:@24697.4]
  assign RetimeWrapper_127_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24699.4]
  assign RetimeWrapper_127_io_in = _T_2587 & io_rPort_10_en_0; // @[package.scala 94:16:@24698.4]
  assign RetimeWrapper_128_clock = clock; // @[:@24704.4]
  assign RetimeWrapper_128_reset = reset; // @[:@24705.4]
  assign RetimeWrapper_128_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24707.4]
  assign RetimeWrapper_128_io_in = _T_2771 & io_rPort_10_en_0; // @[package.scala 94:16:@24706.4]
  assign RetimeWrapper_129_clock = clock; // @[:@24712.4]
  assign RetimeWrapper_129_reset = reset; // @[:@24713.4]
  assign RetimeWrapper_129_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24715.4]
  assign RetimeWrapper_129_io_in = _T_2955 & io_rPort_10_en_0; // @[package.scala 94:16:@24714.4]
  assign RetimeWrapper_130_clock = clock; // @[:@24720.4]
  assign RetimeWrapper_130_reset = reset; // @[:@24721.4]
  assign RetimeWrapper_130_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24723.4]
  assign RetimeWrapper_130_io_in = _T_3139 & io_rPort_10_en_0; // @[package.scala 94:16:@24722.4]
  assign RetimeWrapper_131_clock = clock; // @[:@24728.4]
  assign RetimeWrapper_131_reset = reset; // @[:@24729.4]
  assign RetimeWrapper_131_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24731.4]
  assign RetimeWrapper_131_io_in = _T_3323 & io_rPort_10_en_0; // @[package.scala 94:16:@24730.4]
  assign RetimeWrapper_132_clock = clock; // @[:@24784.4]
  assign RetimeWrapper_132_reset = reset; // @[:@24785.4]
  assign RetimeWrapper_132_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24787.4]
  assign RetimeWrapper_132_io_in = _T_1219 & io_rPort_11_en_0; // @[package.scala 94:16:@24786.4]
  assign RetimeWrapper_133_clock = clock; // @[:@24792.4]
  assign RetimeWrapper_133_reset = reset; // @[:@24793.4]
  assign RetimeWrapper_133_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24795.4]
  assign RetimeWrapper_133_io_in = _T_1403 & io_rPort_11_en_0; // @[package.scala 94:16:@24794.4]
  assign RetimeWrapper_134_clock = clock; // @[:@24800.4]
  assign RetimeWrapper_134_reset = reset; // @[:@24801.4]
  assign RetimeWrapper_134_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24803.4]
  assign RetimeWrapper_134_io_in = _T_1587 & io_rPort_11_en_0; // @[package.scala 94:16:@24802.4]
  assign RetimeWrapper_135_clock = clock; // @[:@24808.4]
  assign RetimeWrapper_135_reset = reset; // @[:@24809.4]
  assign RetimeWrapper_135_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24811.4]
  assign RetimeWrapper_135_io_in = _T_1771 & io_rPort_11_en_0; // @[package.scala 94:16:@24810.4]
  assign RetimeWrapper_136_clock = clock; // @[:@24816.4]
  assign RetimeWrapper_136_reset = reset; // @[:@24817.4]
  assign RetimeWrapper_136_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24819.4]
  assign RetimeWrapper_136_io_in = _T_1955 & io_rPort_11_en_0; // @[package.scala 94:16:@24818.4]
  assign RetimeWrapper_137_clock = clock; // @[:@24824.4]
  assign RetimeWrapper_137_reset = reset; // @[:@24825.4]
  assign RetimeWrapper_137_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24827.4]
  assign RetimeWrapper_137_io_in = _T_2139 & io_rPort_11_en_0; // @[package.scala 94:16:@24826.4]
  assign RetimeWrapper_138_clock = clock; // @[:@24832.4]
  assign RetimeWrapper_138_reset = reset; // @[:@24833.4]
  assign RetimeWrapper_138_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24835.4]
  assign RetimeWrapper_138_io_in = _T_2323 & io_rPort_11_en_0; // @[package.scala 94:16:@24834.4]
  assign RetimeWrapper_139_clock = clock; // @[:@24840.4]
  assign RetimeWrapper_139_reset = reset; // @[:@24841.4]
  assign RetimeWrapper_139_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24843.4]
  assign RetimeWrapper_139_io_in = _T_2507 & io_rPort_11_en_0; // @[package.scala 94:16:@24842.4]
  assign RetimeWrapper_140_clock = clock; // @[:@24848.4]
  assign RetimeWrapper_140_reset = reset; // @[:@24849.4]
  assign RetimeWrapper_140_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24851.4]
  assign RetimeWrapper_140_io_in = _T_2691 & io_rPort_11_en_0; // @[package.scala 94:16:@24850.4]
  assign RetimeWrapper_141_clock = clock; // @[:@24856.4]
  assign RetimeWrapper_141_reset = reset; // @[:@24857.4]
  assign RetimeWrapper_141_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24859.4]
  assign RetimeWrapper_141_io_in = _T_2875 & io_rPort_11_en_0; // @[package.scala 94:16:@24858.4]
  assign RetimeWrapper_142_clock = clock; // @[:@24864.4]
  assign RetimeWrapper_142_reset = reset; // @[:@24865.4]
  assign RetimeWrapper_142_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24867.4]
  assign RetimeWrapper_142_io_in = _T_3059 & io_rPort_11_en_0; // @[package.scala 94:16:@24866.4]
  assign RetimeWrapper_143_clock = clock; // @[:@24872.4]
  assign RetimeWrapper_143_reset = reset; // @[:@24873.4]
  assign RetimeWrapper_143_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24875.4]
  assign RetimeWrapper_143_io_in = _T_3243 & io_rPort_11_en_0; // @[package.scala 94:16:@24874.4]
  assign RetimeWrapper_144_clock = clock; // @[:@24928.4]
  assign RetimeWrapper_144_reset = reset; // @[:@24929.4]
  assign RetimeWrapper_144_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24931.4]
  assign RetimeWrapper_144_io_in = _T_1305 & io_rPort_12_en_0; // @[package.scala 94:16:@24930.4]
  assign RetimeWrapper_145_clock = clock; // @[:@24936.4]
  assign RetimeWrapper_145_reset = reset; // @[:@24937.4]
  assign RetimeWrapper_145_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24939.4]
  assign RetimeWrapper_145_io_in = _T_1489 & io_rPort_12_en_0; // @[package.scala 94:16:@24938.4]
  assign RetimeWrapper_146_clock = clock; // @[:@24944.4]
  assign RetimeWrapper_146_reset = reset; // @[:@24945.4]
  assign RetimeWrapper_146_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24947.4]
  assign RetimeWrapper_146_io_in = _T_1673 & io_rPort_12_en_0; // @[package.scala 94:16:@24946.4]
  assign RetimeWrapper_147_clock = clock; // @[:@24952.4]
  assign RetimeWrapper_147_reset = reset; // @[:@24953.4]
  assign RetimeWrapper_147_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24955.4]
  assign RetimeWrapper_147_io_in = _T_1857 & io_rPort_12_en_0; // @[package.scala 94:16:@24954.4]
  assign RetimeWrapper_148_clock = clock; // @[:@24960.4]
  assign RetimeWrapper_148_reset = reset; // @[:@24961.4]
  assign RetimeWrapper_148_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24963.4]
  assign RetimeWrapper_148_io_in = _T_2041 & io_rPort_12_en_0; // @[package.scala 94:16:@24962.4]
  assign RetimeWrapper_149_clock = clock; // @[:@24968.4]
  assign RetimeWrapper_149_reset = reset; // @[:@24969.4]
  assign RetimeWrapper_149_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24971.4]
  assign RetimeWrapper_149_io_in = _T_2225 & io_rPort_12_en_0; // @[package.scala 94:16:@24970.4]
  assign RetimeWrapper_150_clock = clock; // @[:@24976.4]
  assign RetimeWrapper_150_reset = reset; // @[:@24977.4]
  assign RetimeWrapper_150_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24979.4]
  assign RetimeWrapper_150_io_in = _T_2409 & io_rPort_12_en_0; // @[package.scala 94:16:@24978.4]
  assign RetimeWrapper_151_clock = clock; // @[:@24984.4]
  assign RetimeWrapper_151_reset = reset; // @[:@24985.4]
  assign RetimeWrapper_151_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24987.4]
  assign RetimeWrapper_151_io_in = _T_2593 & io_rPort_12_en_0; // @[package.scala 94:16:@24986.4]
  assign RetimeWrapper_152_clock = clock; // @[:@24992.4]
  assign RetimeWrapper_152_reset = reset; // @[:@24993.4]
  assign RetimeWrapper_152_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24995.4]
  assign RetimeWrapper_152_io_in = _T_2777 & io_rPort_12_en_0; // @[package.scala 94:16:@24994.4]
  assign RetimeWrapper_153_clock = clock; // @[:@25000.4]
  assign RetimeWrapper_153_reset = reset; // @[:@25001.4]
  assign RetimeWrapper_153_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@25003.4]
  assign RetimeWrapper_153_io_in = _T_2961 & io_rPort_12_en_0; // @[package.scala 94:16:@25002.4]
  assign RetimeWrapper_154_clock = clock; // @[:@25008.4]
  assign RetimeWrapper_154_reset = reset; // @[:@25009.4]
  assign RetimeWrapper_154_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@25011.4]
  assign RetimeWrapper_154_io_in = _T_3145 & io_rPort_12_en_0; // @[package.scala 94:16:@25010.4]
  assign RetimeWrapper_155_clock = clock; // @[:@25016.4]
  assign RetimeWrapper_155_reset = reset; // @[:@25017.4]
  assign RetimeWrapper_155_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@25019.4]
  assign RetimeWrapper_155_io_in = _T_3329 & io_rPort_12_en_0; // @[package.scala 94:16:@25018.4]
  assign RetimeWrapper_156_clock = clock; // @[:@25072.4]
  assign RetimeWrapper_156_reset = reset; // @[:@25073.4]
  assign RetimeWrapper_156_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25075.4]
  assign RetimeWrapper_156_io_in = _T_1311 & io_rPort_13_en_0; // @[package.scala 94:16:@25074.4]
  assign RetimeWrapper_157_clock = clock; // @[:@25080.4]
  assign RetimeWrapper_157_reset = reset; // @[:@25081.4]
  assign RetimeWrapper_157_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25083.4]
  assign RetimeWrapper_157_io_in = _T_1495 & io_rPort_13_en_0; // @[package.scala 94:16:@25082.4]
  assign RetimeWrapper_158_clock = clock; // @[:@25088.4]
  assign RetimeWrapper_158_reset = reset; // @[:@25089.4]
  assign RetimeWrapper_158_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25091.4]
  assign RetimeWrapper_158_io_in = _T_1679 & io_rPort_13_en_0; // @[package.scala 94:16:@25090.4]
  assign RetimeWrapper_159_clock = clock; // @[:@25096.4]
  assign RetimeWrapper_159_reset = reset; // @[:@25097.4]
  assign RetimeWrapper_159_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25099.4]
  assign RetimeWrapper_159_io_in = _T_1863 & io_rPort_13_en_0; // @[package.scala 94:16:@25098.4]
  assign RetimeWrapper_160_clock = clock; // @[:@25104.4]
  assign RetimeWrapper_160_reset = reset; // @[:@25105.4]
  assign RetimeWrapper_160_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25107.4]
  assign RetimeWrapper_160_io_in = _T_2047 & io_rPort_13_en_0; // @[package.scala 94:16:@25106.4]
  assign RetimeWrapper_161_clock = clock; // @[:@25112.4]
  assign RetimeWrapper_161_reset = reset; // @[:@25113.4]
  assign RetimeWrapper_161_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25115.4]
  assign RetimeWrapper_161_io_in = _T_2231 & io_rPort_13_en_0; // @[package.scala 94:16:@25114.4]
  assign RetimeWrapper_162_clock = clock; // @[:@25120.4]
  assign RetimeWrapper_162_reset = reset; // @[:@25121.4]
  assign RetimeWrapper_162_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25123.4]
  assign RetimeWrapper_162_io_in = _T_2415 & io_rPort_13_en_0; // @[package.scala 94:16:@25122.4]
  assign RetimeWrapper_163_clock = clock; // @[:@25128.4]
  assign RetimeWrapper_163_reset = reset; // @[:@25129.4]
  assign RetimeWrapper_163_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25131.4]
  assign RetimeWrapper_163_io_in = _T_2599 & io_rPort_13_en_0; // @[package.scala 94:16:@25130.4]
  assign RetimeWrapper_164_clock = clock; // @[:@25136.4]
  assign RetimeWrapper_164_reset = reset; // @[:@25137.4]
  assign RetimeWrapper_164_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25139.4]
  assign RetimeWrapper_164_io_in = _T_2783 & io_rPort_13_en_0; // @[package.scala 94:16:@25138.4]
  assign RetimeWrapper_165_clock = clock; // @[:@25144.4]
  assign RetimeWrapper_165_reset = reset; // @[:@25145.4]
  assign RetimeWrapper_165_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25147.4]
  assign RetimeWrapper_165_io_in = _T_2967 & io_rPort_13_en_0; // @[package.scala 94:16:@25146.4]
  assign RetimeWrapper_166_clock = clock; // @[:@25152.4]
  assign RetimeWrapper_166_reset = reset; // @[:@25153.4]
  assign RetimeWrapper_166_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25155.4]
  assign RetimeWrapper_166_io_in = _T_3151 & io_rPort_13_en_0; // @[package.scala 94:16:@25154.4]
  assign RetimeWrapper_167_clock = clock; // @[:@25160.4]
  assign RetimeWrapper_167_reset = reset; // @[:@25161.4]
  assign RetimeWrapper_167_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25163.4]
  assign RetimeWrapper_167_io_in = _T_3335 & io_rPort_13_en_0; // @[package.scala 94:16:@25162.4]
  assign RetimeWrapper_168_clock = clock; // @[:@25216.4]
  assign RetimeWrapper_168_reset = reset; // @[:@25217.4]
  assign RetimeWrapper_168_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25219.4]
  assign RetimeWrapper_168_io_in = _T_1225 & io_rPort_14_en_0; // @[package.scala 94:16:@25218.4]
  assign RetimeWrapper_169_clock = clock; // @[:@25224.4]
  assign RetimeWrapper_169_reset = reset; // @[:@25225.4]
  assign RetimeWrapper_169_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25227.4]
  assign RetimeWrapper_169_io_in = _T_1409 & io_rPort_14_en_0; // @[package.scala 94:16:@25226.4]
  assign RetimeWrapper_170_clock = clock; // @[:@25232.4]
  assign RetimeWrapper_170_reset = reset; // @[:@25233.4]
  assign RetimeWrapper_170_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25235.4]
  assign RetimeWrapper_170_io_in = _T_1593 & io_rPort_14_en_0; // @[package.scala 94:16:@25234.4]
  assign RetimeWrapper_171_clock = clock; // @[:@25240.4]
  assign RetimeWrapper_171_reset = reset; // @[:@25241.4]
  assign RetimeWrapper_171_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25243.4]
  assign RetimeWrapper_171_io_in = _T_1777 & io_rPort_14_en_0; // @[package.scala 94:16:@25242.4]
  assign RetimeWrapper_172_clock = clock; // @[:@25248.4]
  assign RetimeWrapper_172_reset = reset; // @[:@25249.4]
  assign RetimeWrapper_172_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25251.4]
  assign RetimeWrapper_172_io_in = _T_1961 & io_rPort_14_en_0; // @[package.scala 94:16:@25250.4]
  assign RetimeWrapper_173_clock = clock; // @[:@25256.4]
  assign RetimeWrapper_173_reset = reset; // @[:@25257.4]
  assign RetimeWrapper_173_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25259.4]
  assign RetimeWrapper_173_io_in = _T_2145 & io_rPort_14_en_0; // @[package.scala 94:16:@25258.4]
  assign RetimeWrapper_174_clock = clock; // @[:@25264.4]
  assign RetimeWrapper_174_reset = reset; // @[:@25265.4]
  assign RetimeWrapper_174_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25267.4]
  assign RetimeWrapper_174_io_in = _T_2329 & io_rPort_14_en_0; // @[package.scala 94:16:@25266.4]
  assign RetimeWrapper_175_clock = clock; // @[:@25272.4]
  assign RetimeWrapper_175_reset = reset; // @[:@25273.4]
  assign RetimeWrapper_175_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25275.4]
  assign RetimeWrapper_175_io_in = _T_2513 & io_rPort_14_en_0; // @[package.scala 94:16:@25274.4]
  assign RetimeWrapper_176_clock = clock; // @[:@25280.4]
  assign RetimeWrapper_176_reset = reset; // @[:@25281.4]
  assign RetimeWrapper_176_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25283.4]
  assign RetimeWrapper_176_io_in = _T_2697 & io_rPort_14_en_0; // @[package.scala 94:16:@25282.4]
  assign RetimeWrapper_177_clock = clock; // @[:@25288.4]
  assign RetimeWrapper_177_reset = reset; // @[:@25289.4]
  assign RetimeWrapper_177_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25291.4]
  assign RetimeWrapper_177_io_in = _T_2881 & io_rPort_14_en_0; // @[package.scala 94:16:@25290.4]
  assign RetimeWrapper_178_clock = clock; // @[:@25296.4]
  assign RetimeWrapper_178_reset = reset; // @[:@25297.4]
  assign RetimeWrapper_178_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25299.4]
  assign RetimeWrapper_178_io_in = _T_3065 & io_rPort_14_en_0; // @[package.scala 94:16:@25298.4]
  assign RetimeWrapper_179_clock = clock; // @[:@25304.4]
  assign RetimeWrapper_179_reset = reset; // @[:@25305.4]
  assign RetimeWrapper_179_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25307.4]
  assign RetimeWrapper_179_io_in = _T_3249 & io_rPort_14_en_0; // @[package.scala 94:16:@25306.4]
  assign RetimeWrapper_180_clock = clock; // @[:@25360.4]
  assign RetimeWrapper_180_reset = reset; // @[:@25361.4]
  assign RetimeWrapper_180_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25363.4]
  assign RetimeWrapper_180_io_in = _T_1317 & io_rPort_15_en_0; // @[package.scala 94:16:@25362.4]
  assign RetimeWrapper_181_clock = clock; // @[:@25368.4]
  assign RetimeWrapper_181_reset = reset; // @[:@25369.4]
  assign RetimeWrapper_181_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25371.4]
  assign RetimeWrapper_181_io_in = _T_1501 & io_rPort_15_en_0; // @[package.scala 94:16:@25370.4]
  assign RetimeWrapper_182_clock = clock; // @[:@25376.4]
  assign RetimeWrapper_182_reset = reset; // @[:@25377.4]
  assign RetimeWrapper_182_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25379.4]
  assign RetimeWrapper_182_io_in = _T_1685 & io_rPort_15_en_0; // @[package.scala 94:16:@25378.4]
  assign RetimeWrapper_183_clock = clock; // @[:@25384.4]
  assign RetimeWrapper_183_reset = reset; // @[:@25385.4]
  assign RetimeWrapper_183_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25387.4]
  assign RetimeWrapper_183_io_in = _T_1869 & io_rPort_15_en_0; // @[package.scala 94:16:@25386.4]
  assign RetimeWrapper_184_clock = clock; // @[:@25392.4]
  assign RetimeWrapper_184_reset = reset; // @[:@25393.4]
  assign RetimeWrapper_184_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25395.4]
  assign RetimeWrapper_184_io_in = _T_2053 & io_rPort_15_en_0; // @[package.scala 94:16:@25394.4]
  assign RetimeWrapper_185_clock = clock; // @[:@25400.4]
  assign RetimeWrapper_185_reset = reset; // @[:@25401.4]
  assign RetimeWrapper_185_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25403.4]
  assign RetimeWrapper_185_io_in = _T_2237 & io_rPort_15_en_0; // @[package.scala 94:16:@25402.4]
  assign RetimeWrapper_186_clock = clock; // @[:@25408.4]
  assign RetimeWrapper_186_reset = reset; // @[:@25409.4]
  assign RetimeWrapper_186_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25411.4]
  assign RetimeWrapper_186_io_in = _T_2421 & io_rPort_15_en_0; // @[package.scala 94:16:@25410.4]
  assign RetimeWrapper_187_clock = clock; // @[:@25416.4]
  assign RetimeWrapper_187_reset = reset; // @[:@25417.4]
  assign RetimeWrapper_187_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25419.4]
  assign RetimeWrapper_187_io_in = _T_2605 & io_rPort_15_en_0; // @[package.scala 94:16:@25418.4]
  assign RetimeWrapper_188_clock = clock; // @[:@25424.4]
  assign RetimeWrapper_188_reset = reset; // @[:@25425.4]
  assign RetimeWrapper_188_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25427.4]
  assign RetimeWrapper_188_io_in = _T_2789 & io_rPort_15_en_0; // @[package.scala 94:16:@25426.4]
  assign RetimeWrapper_189_clock = clock; // @[:@25432.4]
  assign RetimeWrapper_189_reset = reset; // @[:@25433.4]
  assign RetimeWrapper_189_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25435.4]
  assign RetimeWrapper_189_io_in = _T_2973 & io_rPort_15_en_0; // @[package.scala 94:16:@25434.4]
  assign RetimeWrapper_190_clock = clock; // @[:@25440.4]
  assign RetimeWrapper_190_reset = reset; // @[:@25441.4]
  assign RetimeWrapper_190_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25443.4]
  assign RetimeWrapper_190_io_in = _T_3157 & io_rPort_15_en_0; // @[package.scala 94:16:@25442.4]
  assign RetimeWrapper_191_clock = clock; // @[:@25448.4]
  assign RetimeWrapper_191_reset = reset; // @[:@25449.4]
  assign RetimeWrapper_191_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25451.4]
  assign RetimeWrapper_191_io_in = _T_3341 & io_rPort_15_en_0; // @[package.scala 94:16:@25450.4]
  assign RetimeWrapper_192_clock = clock; // @[:@25504.4]
  assign RetimeWrapper_192_reset = reset; // @[:@25505.4]
  assign RetimeWrapper_192_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25507.4]
  assign RetimeWrapper_192_io_in = _T_1231 & io_rPort_16_en_0; // @[package.scala 94:16:@25506.4]
  assign RetimeWrapper_193_clock = clock; // @[:@25512.4]
  assign RetimeWrapper_193_reset = reset; // @[:@25513.4]
  assign RetimeWrapper_193_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25515.4]
  assign RetimeWrapper_193_io_in = _T_1415 & io_rPort_16_en_0; // @[package.scala 94:16:@25514.4]
  assign RetimeWrapper_194_clock = clock; // @[:@25520.4]
  assign RetimeWrapper_194_reset = reset; // @[:@25521.4]
  assign RetimeWrapper_194_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25523.4]
  assign RetimeWrapper_194_io_in = _T_1599 & io_rPort_16_en_0; // @[package.scala 94:16:@25522.4]
  assign RetimeWrapper_195_clock = clock; // @[:@25528.4]
  assign RetimeWrapper_195_reset = reset; // @[:@25529.4]
  assign RetimeWrapper_195_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25531.4]
  assign RetimeWrapper_195_io_in = _T_1783 & io_rPort_16_en_0; // @[package.scala 94:16:@25530.4]
  assign RetimeWrapper_196_clock = clock; // @[:@25536.4]
  assign RetimeWrapper_196_reset = reset; // @[:@25537.4]
  assign RetimeWrapper_196_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25539.4]
  assign RetimeWrapper_196_io_in = _T_1967 & io_rPort_16_en_0; // @[package.scala 94:16:@25538.4]
  assign RetimeWrapper_197_clock = clock; // @[:@25544.4]
  assign RetimeWrapper_197_reset = reset; // @[:@25545.4]
  assign RetimeWrapper_197_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25547.4]
  assign RetimeWrapper_197_io_in = _T_2151 & io_rPort_16_en_0; // @[package.scala 94:16:@25546.4]
  assign RetimeWrapper_198_clock = clock; // @[:@25552.4]
  assign RetimeWrapper_198_reset = reset; // @[:@25553.4]
  assign RetimeWrapper_198_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25555.4]
  assign RetimeWrapper_198_io_in = _T_2335 & io_rPort_16_en_0; // @[package.scala 94:16:@25554.4]
  assign RetimeWrapper_199_clock = clock; // @[:@25560.4]
  assign RetimeWrapper_199_reset = reset; // @[:@25561.4]
  assign RetimeWrapper_199_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25563.4]
  assign RetimeWrapper_199_io_in = _T_2519 & io_rPort_16_en_0; // @[package.scala 94:16:@25562.4]
  assign RetimeWrapper_200_clock = clock; // @[:@25568.4]
  assign RetimeWrapper_200_reset = reset; // @[:@25569.4]
  assign RetimeWrapper_200_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25571.4]
  assign RetimeWrapper_200_io_in = _T_2703 & io_rPort_16_en_0; // @[package.scala 94:16:@25570.4]
  assign RetimeWrapper_201_clock = clock; // @[:@25576.4]
  assign RetimeWrapper_201_reset = reset; // @[:@25577.4]
  assign RetimeWrapper_201_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25579.4]
  assign RetimeWrapper_201_io_in = _T_2887 & io_rPort_16_en_0; // @[package.scala 94:16:@25578.4]
  assign RetimeWrapper_202_clock = clock; // @[:@25584.4]
  assign RetimeWrapper_202_reset = reset; // @[:@25585.4]
  assign RetimeWrapper_202_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25587.4]
  assign RetimeWrapper_202_io_in = _T_3071 & io_rPort_16_en_0; // @[package.scala 94:16:@25586.4]
  assign RetimeWrapper_203_clock = clock; // @[:@25592.4]
  assign RetimeWrapper_203_reset = reset; // @[:@25593.4]
  assign RetimeWrapper_203_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25595.4]
  assign RetimeWrapper_203_io_in = _T_3255 & io_rPort_16_en_0; // @[package.scala 94:16:@25594.4]
  assign RetimeWrapper_204_clock = clock; // @[:@25648.4]
  assign RetimeWrapper_204_reset = reset; // @[:@25649.4]
  assign RetimeWrapper_204_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25651.4]
  assign RetimeWrapper_204_io_in = _T_1323 & io_rPort_17_en_0; // @[package.scala 94:16:@25650.4]
  assign RetimeWrapper_205_clock = clock; // @[:@25656.4]
  assign RetimeWrapper_205_reset = reset; // @[:@25657.4]
  assign RetimeWrapper_205_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25659.4]
  assign RetimeWrapper_205_io_in = _T_1507 & io_rPort_17_en_0; // @[package.scala 94:16:@25658.4]
  assign RetimeWrapper_206_clock = clock; // @[:@25664.4]
  assign RetimeWrapper_206_reset = reset; // @[:@25665.4]
  assign RetimeWrapper_206_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25667.4]
  assign RetimeWrapper_206_io_in = _T_1691 & io_rPort_17_en_0; // @[package.scala 94:16:@25666.4]
  assign RetimeWrapper_207_clock = clock; // @[:@25672.4]
  assign RetimeWrapper_207_reset = reset; // @[:@25673.4]
  assign RetimeWrapper_207_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25675.4]
  assign RetimeWrapper_207_io_in = _T_1875 & io_rPort_17_en_0; // @[package.scala 94:16:@25674.4]
  assign RetimeWrapper_208_clock = clock; // @[:@25680.4]
  assign RetimeWrapper_208_reset = reset; // @[:@25681.4]
  assign RetimeWrapper_208_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25683.4]
  assign RetimeWrapper_208_io_in = _T_2059 & io_rPort_17_en_0; // @[package.scala 94:16:@25682.4]
  assign RetimeWrapper_209_clock = clock; // @[:@25688.4]
  assign RetimeWrapper_209_reset = reset; // @[:@25689.4]
  assign RetimeWrapper_209_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25691.4]
  assign RetimeWrapper_209_io_in = _T_2243 & io_rPort_17_en_0; // @[package.scala 94:16:@25690.4]
  assign RetimeWrapper_210_clock = clock; // @[:@25696.4]
  assign RetimeWrapper_210_reset = reset; // @[:@25697.4]
  assign RetimeWrapper_210_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25699.4]
  assign RetimeWrapper_210_io_in = _T_2427 & io_rPort_17_en_0; // @[package.scala 94:16:@25698.4]
  assign RetimeWrapper_211_clock = clock; // @[:@25704.4]
  assign RetimeWrapper_211_reset = reset; // @[:@25705.4]
  assign RetimeWrapper_211_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25707.4]
  assign RetimeWrapper_211_io_in = _T_2611 & io_rPort_17_en_0; // @[package.scala 94:16:@25706.4]
  assign RetimeWrapper_212_clock = clock; // @[:@25712.4]
  assign RetimeWrapper_212_reset = reset; // @[:@25713.4]
  assign RetimeWrapper_212_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25715.4]
  assign RetimeWrapper_212_io_in = _T_2795 & io_rPort_17_en_0; // @[package.scala 94:16:@25714.4]
  assign RetimeWrapper_213_clock = clock; // @[:@25720.4]
  assign RetimeWrapper_213_reset = reset; // @[:@25721.4]
  assign RetimeWrapper_213_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25723.4]
  assign RetimeWrapper_213_io_in = _T_2979 & io_rPort_17_en_0; // @[package.scala 94:16:@25722.4]
  assign RetimeWrapper_214_clock = clock; // @[:@25728.4]
  assign RetimeWrapper_214_reset = reset; // @[:@25729.4]
  assign RetimeWrapper_214_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25731.4]
  assign RetimeWrapper_214_io_in = _T_3163 & io_rPort_17_en_0; // @[package.scala 94:16:@25730.4]
  assign RetimeWrapper_215_clock = clock; // @[:@25736.4]
  assign RetimeWrapper_215_reset = reset; // @[:@25737.4]
  assign RetimeWrapper_215_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25739.4]
  assign RetimeWrapper_215_io_in = _T_3347 & io_rPort_17_en_0; // @[package.scala 94:16:@25738.4]
endmodule
module Modulo( // @[:@25768.2]
  input         clock, // @[:@25769.4]
  input         io_flow, // @[:@25771.4]
  input  [31:0] io_dividend, // @[:@25771.4]
  input  [31:0] io_divisor, // @[:@25771.4]
  output [31:0] io_out // @[:@25771.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  div_32_32_16_Unsigned_Remainder m ( // @[ZynqBlackBoxes.scala 48:19:@25773.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign io_out = m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 56:12:@25789.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 54:31:@25787.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 53:32:@25786.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 52:32:@25785.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 51:33:@25784.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 50:17:@25783.4 ZynqBlackBoxes.scala 55:17:@25788.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 49:15:@25782.4]
endmodule
module fix2fixBox_38( // @[:@25791.2]
  input  [63:0] io_a, // @[:@25794.4]
  output [31:0] io_b // @[:@25794.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@25807.4]
endmodule
module x403( // @[:@25809.2]
  input         clock, // @[:@25810.4]
  input  [31:0] io_a, // @[:@25812.4]
  input         io_flow, // @[:@25812.4]
  output [31:0] io_result // @[:@25812.4]
);
  wire  x403_clock; // @[BigIPZynq.scala 35:21:@25820.4]
  wire  x403_io_flow; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [31:0] x403_io_dividend; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [31:0] x403_io_divisor; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [31:0] x403_io_out; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@25827.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@25827.4]
  Modulo x403 ( // @[BigIPZynq.scala 35:21:@25820.4]
    .clock(x403_clock),
    .io_flow(x403_io_flow),
    .io_dividend(x403_io_dividend),
    .io_divisor(x403_io_divisor),
    .io_out(x403_io_out)
  );
  fix2fixBox_38 fix2fixBox ( // @[Math.scala 357:30:@25827.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@25835.4]
  assign x403_clock = clock; // @[:@25821.4]
  assign x403_io_flow = io_flow; // @[BigIPZynq.scala 38:17:@25825.4]
  assign x403_io_dividend = io_a; // @[BigIPZynq.scala 36:21:@25823.4]
  assign x403_io_divisor = 32'h6; // @[BigIPZynq.scala 37:20:@25824.4]
  assign fix2fixBox_io_a = {{32'd0}, x403_io_out}; // @[Math.scala 358:23:@25830.4]
endmodule
module Divider( // @[:@26029.2]
  input         clock, // @[:@26030.4]
  input         io_flow, // @[:@26032.4]
  input  [31:0] io_dividend, // @[:@26032.4]
  input  [31:0] io_divisor, // @[:@26032.4]
  output [31:0] io_out // @[:@26032.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire [29:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@26050.4]
  div_32_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@26034.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[31:2]; // @[ZynqBlackBoxes.scala 34:37:@26050.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@26051.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@26048.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@26047.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@26046.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@26045.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@26044.4 ZynqBlackBoxes.scala 33:17:@26049.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@26043.4]
endmodule
module x406_div( // @[:@26089.2]
  input         clock, // @[:@26090.4]
  input  [31:0] io_a, // @[:@26092.4]
  input         io_flow, // @[:@26092.4]
  output [31:0] io_result // @[:@26092.4]
);
  wire  x406_div_clock; // @[BigIPZynq.scala 25:21:@26100.4]
  wire  x406_div_io_flow; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] x406_div_io_dividend; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] x406_div_io_divisor; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] x406_div_io_out; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@26113.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@26113.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@26098.4]
  wire [31:0] _T_19; // @[BigIPZynq.scala 29:16:@26108.4]
  Divider x406_div ( // @[BigIPZynq.scala 25:21:@26100.4]
    .clock(x406_div_clock),
    .io_flow(x406_div_io_flow),
    .io_dividend(x406_div_io_dividend),
    .io_divisor(x406_div_io_divisor),
    .io_out(x406_div_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@26113.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@26098.4]
  assign _T_19 = $signed(x406_div_io_out); // @[BigIPZynq.scala 29:16:@26108.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@26121.4]
  assign x406_div_clock = clock; // @[:@26101.4]
  assign x406_div_io_flow = io_flow; // @[BigIPZynq.scala 28:17:@26107.4]
  assign x406_div_io_dividend = $unsigned(_T_15); // @[BigIPZynq.scala 26:21:@26104.4]
  assign x406_div_io_divisor = 32'h6; // @[BigIPZynq.scala 27:20:@26106.4]
  assign __io_b = $unsigned(_T_19); // @[Math.scala 721:17:@26116.4]
endmodule
module RetimeWrapper_298( // @[:@26135.2]
  input         clock, // @[:@26136.4]
  input         reset, // @[:@26137.4]
  input         io_flow, // @[:@26138.4]
  input  [31:0] io_in, // @[:@26138.4]
  output [31:0] io_out // @[:@26138.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@26140.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26153.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26152.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26151.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26150.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26149.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26147.4]
endmodule
module RetimeWrapper_300( // @[:@26346.2]
  input         clock, // @[:@26347.4]
  input         reset, // @[:@26348.4]
  input         io_flow, // @[:@26349.4]
  input  [31:0] io_in, // @[:@26349.4]
  output [31:0] io_out // @[:@26349.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26351.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26364.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26363.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26362.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26361.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26360.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26358.4]
endmodule
module RetimeWrapper_301( // @[:@26378.2]
  input         clock, // @[:@26379.4]
  input         reset, // @[:@26380.4]
  input         io_flow, // @[:@26381.4]
  input  [31:0] io_in, // @[:@26381.4]
  output [31:0] io_out // @[:@26381.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@26383.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26396.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26395.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26394.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26393.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26392.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26390.4]
endmodule
module RetimeWrapper_302( // @[:@26410.2]
  input         clock, // @[:@26411.4]
  input         reset, // @[:@26412.4]
  input         io_flow, // @[:@26413.4]
  input  [31:0] io_in, // @[:@26413.4]
  output [31:0] io_out // @[:@26413.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@26415.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26428.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26427.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26426.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26425.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26424.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26422.4]
endmodule
module RetimeWrapper_303( // @[:@26442.2]
  input   clock, // @[:@26443.4]
  input   reset, // @[:@26444.4]
  input   io_flow, // @[:@26445.4]
  input   io_in, // @[:@26445.4]
  output  io_out // @[:@26445.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@26447.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26460.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26459.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@26458.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26457.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26456.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26454.4]
endmodule
module RetimeWrapper_304( // @[:@26474.2]
  input         clock, // @[:@26475.4]
  input         reset, // @[:@26476.4]
  input         io_flow, // @[:@26477.4]
  input  [31:0] io_in, // @[:@26477.4]
  output [31:0] io_out // @[:@26477.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26479.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26479.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26479.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26479.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26479.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26479.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@26479.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26492.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26491.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26490.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26489.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26488.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26486.4]
endmodule
module RetimeWrapper_308( // @[:@26938.2]
  input         clock, // @[:@26939.4]
  input         reset, // @[:@26940.4]
  input         io_flow, // @[:@26941.4]
  input  [31:0] io_in, // @[:@26941.4]
  output [31:0] io_out // @[:@26941.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@26943.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26956.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26955.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26954.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26953.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26952.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26950.4]
endmodule
module RetimeWrapper_310( // @[:@27149.2]
  input         clock, // @[:@27150.4]
  input         reset, // @[:@27151.4]
  input         io_flow, // @[:@27152.4]
  input  [31:0] io_in, // @[:@27152.4]
  output [31:0] io_out // @[:@27152.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@27154.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27167.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27166.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27165.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27164.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27163.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27161.4]
endmodule
module RetimeWrapper_311( // @[:@27181.2]
  input         clock, // @[:@27182.4]
  input         reset, // @[:@27183.4]
  input         io_flow, // @[:@27184.4]
  input  [31:0] io_in, // @[:@27184.4]
  output [31:0] io_out // @[:@27184.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@27186.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27199.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27198.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27197.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27196.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27195.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27193.4]
endmodule
module RetimeWrapper_326( // @[:@28627.2]
  input         clock, // @[:@28628.4]
  input         reset, // @[:@28629.4]
  input         io_flow, // @[:@28630.4]
  input  [31:0] io_in, // @[:@28630.4]
  output [31:0] io_out // @[:@28630.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@28632.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28645.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28644.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@28643.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28642.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28641.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28639.4]
endmodule
module RetimeWrapper_331( // @[:@28787.2]
  input         clock, // @[:@28788.4]
  input         reset, // @[:@28789.4]
  input         io_flow, // @[:@28790.4]
  input  [31:0] io_in, // @[:@28790.4]
  output [31:0] io_out // @[:@28790.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@28792.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@28792.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@28792.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28792.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28792.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28792.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@28792.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28805.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28804.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@28803.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28802.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28801.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28799.4]
endmodule
module RetimeWrapper_333( // @[:@28851.2]
  input         clock, // @[:@28852.4]
  input         reset, // @[:@28853.4]
  input         io_flow, // @[:@28854.4]
  input  [31:0] io_in, // @[:@28854.4]
  output [31:0] io_out // @[:@28854.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(31)) sr ( // @[RetimeShiftRegister.scala 15:20:@28856.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28869.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28868.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@28867.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28866.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28865.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28863.4]
endmodule
module RetimeWrapper_334( // @[:@28883.2]
  input   clock, // @[:@28884.4]
  input   reset, // @[:@28885.4]
  input   io_flow, // @[:@28886.4]
  input   io_in, // @[:@28886.4]
  output  io_out // @[:@28886.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@28888.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28901.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28900.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@28899.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28898.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28897.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28895.4]
endmodule
module RetimeWrapper_335( // @[:@28915.2]
  input   clock, // @[:@28916.4]
  input   reset, // @[:@28917.4]
  input   io_flow, // @[:@28918.4]
  input   io_in, // @[:@28918.4]
  output  io_out // @[:@28918.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@28920.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@28920.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@28920.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28920.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28920.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28920.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@28920.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28933.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28932.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@28931.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28930.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28929.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28927.4]
endmodule
module RetimeWrapper_352( // @[:@29459.2]
  input         clock, // @[:@29460.4]
  input         reset, // @[:@29461.4]
  input         io_flow, // @[:@29462.4]
  input  [31:0] io_in, // @[:@29462.4]
  output [31:0] io_out // @[:@29462.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@29464.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29477.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29476.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29475.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29474.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29473.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29471.4]
endmodule
module RetimeWrapper_353( // @[:@29491.2]
  input         clock, // @[:@29492.4]
  input         reset, // @[:@29493.4]
  input         io_flow, // @[:@29494.4]
  input  [31:0] io_in, // @[:@29494.4]
  output [31:0] io_out // @[:@29494.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(32)) sr ( // @[RetimeShiftRegister.scala 15:20:@29496.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29509.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29508.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29507.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29506.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29505.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29503.4]
endmodule
module RetimeWrapper_354( // @[:@29523.2]
  input   clock, // @[:@29524.4]
  input   reset, // @[:@29525.4]
  input   io_flow, // @[:@29526.4]
  input   io_in, // @[:@29526.4]
  output  io_out // @[:@29526.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@29528.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29541.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29540.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29539.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29538.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29537.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29535.4]
endmodule
module RetimeWrapper_358( // @[:@29987.2]
  input         clock, // @[:@29988.4]
  input         reset, // @[:@29989.4]
  input         io_flow, // @[:@29990.4]
  input  [31:0] io_in, // @[:@29990.4]
  output [31:0] io_out // @[:@29990.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(46)) sr ( // @[RetimeShiftRegister.scala 15:20:@29992.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30005.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30004.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30003.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30002.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30001.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29999.4]
endmodule
module RetimeWrapper_360( // @[:@30198.2]
  input         clock, // @[:@30199.4]
  input         reset, // @[:@30200.4]
  input         io_flow, // @[:@30201.4]
  input  [31:0] io_in, // @[:@30201.4]
  output [31:0] io_out // @[:@30201.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@30203.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30216.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30215.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30214.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30213.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30212.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30210.4]
endmodule
module RetimeWrapper_374( // @[:@31424.2]
  input         clock, // @[:@31425.4]
  input         reset, // @[:@31426.4]
  input         io_flow, // @[:@31427.4]
  input  [31:0] io_in, // @[:@31427.4]
  output [31:0] io_out // @[:@31427.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@31429.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31442.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31441.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31440.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31439.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31438.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31436.4]
endmodule
module RetimeWrapper_390( // @[:@32377.2]
  input         clock, // @[:@32378.4]
  input         reset, // @[:@32379.4]
  input         io_flow, // @[:@32380.4]
  input  [31:0] io_in, // @[:@32380.4]
  output [31:0] io_out // @[:@32380.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@32382.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@32395.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@32394.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@32393.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@32392.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@32391.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@32389.4]
endmodule
module fix2fixBox_134( // @[:@35199.2]
  input  [31:0] io_a, // @[:@35202.4]
  output [32:0] io_b // @[:@35202.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@35216.4]
endmodule
module __86( // @[:@35218.2]
  input  [31:0] io_b, // @[:@35221.4]
  output [32:0] io_result // @[:@35221.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@35226.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@35226.4]
  fix2fixBox_134 fix2fixBox ( // @[BigIPZynq.scala 219:30:@35226.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@35234.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@35229.4]
endmodule
module x544_x13( // @[:@35330.2]
  input         clock, // @[:@35331.4]
  input         reset, // @[:@35332.4]
  input  [31:0] io_a, // @[:@35333.4]
  input  [31:0] io_b, // @[:@35333.4]
  input         io_flow, // @[:@35333.4]
  output [31:0] io_result // @[:@35333.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@35341.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@35341.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@35348.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@35348.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@35358.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@35358.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@35358.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@35358.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@35358.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@35346.4 Math.scala 724:14:@35347.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@35353.4 Math.scala 724:14:@35354.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@35355.4]
  __86 _ ( // @[Math.scala 720:24:@35341.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __86 __1 ( // @[Math.scala 720:24:@35348.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@35358.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@35346.4 Math.scala 724:14:@35347.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@35353.4 Math.scala 724:14:@35354.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@35355.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@35366.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@35344.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@35351.4]
  assign fix2fixBox_clock = clock; // @[:@35359.4]
  assign fix2fixBox_reset = reset; // @[:@35360.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@35361.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@35364.4]
endmodule
module fix2fixBox_158( // @[:@36583.2]
  input  [31:0] io_a, // @[:@36586.4]
  output [31:0] io_b // @[:@36586.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@36596.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@36596.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@36599.4]
endmodule
module x552( // @[:@36601.2]
  input  [31:0] io_b, // @[:@36604.4]
  output [31:0] io_result // @[:@36604.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@36609.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@36609.4]
  fix2fixBox_158 fix2fixBox ( // @[BigIPZynq.scala 219:30:@36609.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@36617.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@36612.4]
endmodule
module Multiplier( // @[:@36629.2]
  input         clock, // @[:@36630.4]
  input         io_flow, // @[:@36632.4]
  input  [38:0] io_a, // @[:@36632.4]
  input  [38:0] io_b, // @[:@36632.4]
  output [38:0] io_out // @[:@36632.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@36634.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@36634.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@36634.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@36634.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@36634.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@36634.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@36644.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@36642.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@36641.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@36643.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@36640.4]
endmodule
module fix2fixBox_159( // @[:@36646.2]
  input  [38:0] io_a, // @[:@36649.4]
  output [31:0] io_b // @[:@36649.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@36657.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@36660.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@36657.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@36660.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@36663.4]
endmodule
module x553_mul( // @[:@36665.2]
  input         clock, // @[:@36666.4]
  input  [31:0] io_a, // @[:@36668.4]
  input  [31:0] io_b, // @[:@36668.4]
  input         io_flow, // @[:@36668.4]
  output [31:0] io_result // @[:@36668.4]
);
  wire  x553_mul_clock; // @[BigIPZynq.scala 63:21:@36683.4]
  wire  x553_mul_io_flow; // @[BigIPZynq.scala 63:21:@36683.4]
  wire [38:0] x553_mul_io_a; // @[BigIPZynq.scala 63:21:@36683.4]
  wire [38:0] x553_mul_io_b; // @[BigIPZynq.scala 63:21:@36683.4]
  wire [38:0] x553_mul_io_out; // @[BigIPZynq.scala 63:21:@36683.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@36691.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@36691.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@36675.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@36677.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@36679.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@36681.4]
  Multiplier x553_mul ( // @[BigIPZynq.scala 63:21:@36683.4]
    .clock(x553_mul_clock),
    .io_flow(x553_mul_io_flow),
    .io_a(x553_mul_io_a),
    .io_b(x553_mul_io_b),
    .io_out(x553_mul_io_out)
  );
  fix2fixBox_159 fix2fixBox ( // @[Math.scala 253:30:@36691.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@36675.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@36677.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@36679.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@36681.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@36699.4]
  assign x553_mul_clock = clock; // @[:@36684.4]
  assign x553_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@36688.4]
  assign x553_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@36686.4]
  assign x553_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@36687.4]
  assign fix2fixBox_io_a = x553_mul_io_out; // @[Math.scala 254:23:@36694.4]
endmodule
module fix2fixBox_160( // @[:@36701.2]
  input  [31:0] io_a, // @[:@36704.4]
  output [31:0] io_b // @[:@36704.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@36716.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@36716.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@36719.4]
endmodule
module x554( // @[:@36721.2]
  input  [31:0] io_b, // @[:@36724.4]
  output [31:0] io_result // @[:@36724.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@36729.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@36729.4]
  fix2fixBox_160 fix2fixBox ( // @[BigIPZynq.scala 219:30:@36729.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@36737.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@36732.4]
endmodule
module RetimeWrapper_437( // @[:@36751.2]
  input         clock, // @[:@36752.4]
  input         reset, // @[:@36753.4]
  input         io_flow, // @[:@36754.4]
  input  [31:0] io_in, // @[:@36754.4]
  output [31:0] io_out // @[:@36754.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36756.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36756.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36756.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36756.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36756.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36756.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(10)) sr ( // @[RetimeShiftRegister.scala 15:20:@36756.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36769.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36768.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@36767.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36766.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36765.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36763.4]
endmodule
module x555_sub( // @[:@36902.2]
  input         clock, // @[:@36903.4]
  input         reset, // @[:@36904.4]
  input  [31:0] io_a, // @[:@36905.4]
  input  [31:0] io_b, // @[:@36905.4]
  input         io_flow, // @[:@36905.4]
  output [31:0] io_result // @[:@36905.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@36913.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@36913.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@36920.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@36920.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@36931.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@36931.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@36931.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@36931.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@36931.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@36918.4 Math.scala 724:14:@36919.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@36925.4 Math.scala 724:14:@36926.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@36927.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@36928.4]
  __86 _ ( // @[Math.scala 720:24:@36913.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __86 __1 ( // @[Math.scala 720:24:@36920.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@36931.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@36918.4 Math.scala 724:14:@36919.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@36925.4 Math.scala 724:14:@36926.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@36927.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@36928.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@36939.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@36916.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@36923.4]
  assign fix2fixBox_clock = clock; // @[:@36932.4]
  assign fix2fixBox_reset = reset; // @[:@36933.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@36934.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@36937.4]
endmodule
module RetimeWrapper_496( // @[:@44671.2]
  input          clock, // @[:@44672.4]
  input          reset, // @[:@44673.4]
  input          io_flow, // @[:@44674.4]
  input  [127:0] io_in, // @[:@44674.4]
  output [127:0] io_out // @[:@44674.4]
);
  wire [127:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@44676.4]
  wire [127:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@44676.4]
  wire [127:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@44676.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@44676.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@44676.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@44676.4]
  RetimeShiftRegister #(.WIDTH(128), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@44676.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@44689.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@44688.4]
  assign sr_init = 128'h0; // @[RetimeShiftRegister.scala 19:16:@44687.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@44686.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@44685.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@44683.4]
endmodule
module x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@44787.2]
  input          clock, // @[:@44788.4]
  input          reset, // @[:@44789.4]
  output         io_in_x353_TREADY, // @[:@44790.4]
  input  [255:0] io_in_x353_TDATA, // @[:@44790.4]
  input  [7:0]   io_in_x353_TID, // @[:@44790.4]
  input  [7:0]   io_in_x353_TDEST, // @[:@44790.4]
  output         io_in_x354_TVALID, // @[:@44790.4]
  input          io_in_x354_TREADY, // @[:@44790.4]
  output [255:0] io_in_x354_TDATA, // @[:@44790.4]
  input          io_sigsIn_backpressure, // @[:@44790.4]
  input          io_sigsIn_datapathEn, // @[:@44790.4]
  input          io_sigsIn_break, // @[:@44790.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@44790.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@44790.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@44790.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@44790.4]
  input          io_rr // @[:@44790.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@44804.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@44804.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@44816.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@44816.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@44839.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@44839.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@44839.4]
  wire [127:0] RetimeWrapper_io_in; // @[package.scala 93:22:@44839.4]
  wire [127:0] RetimeWrapper_io_out; // @[package.scala 93:22:@44839.4]
  wire  x398_lb_0_clock; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_reset; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_17_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_17_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_17_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_17_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_17_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_17_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_16_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_16_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_16_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_16_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_16_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_16_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_15_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_15_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_15_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_15_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_15_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_15_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_14_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_14_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_14_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_14_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_14_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_14_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_13_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_13_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_13_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_13_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_13_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_13_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_12_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_12_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_12_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_12_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_12_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_12_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_11_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_11_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_11_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_11_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_11_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_11_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_10_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_10_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_10_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_10_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_10_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_10_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_9_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_9_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_9_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_9_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_9_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_9_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_8_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_8_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_8_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_8_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_8_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_8_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_7_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_7_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_7_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_7_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_7_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_7_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_6_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_6_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_6_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_6_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_6_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_6_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_5_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_5_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_5_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_5_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_5_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_5_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_4_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_4_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_4_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_4_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_4_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_4_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_3_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_3_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_3_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_3_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_3_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_3_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_2_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_2_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_2_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_2_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_2_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_2_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_1_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_1_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_1_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_1_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_1_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_1_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_0_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_rPort_0_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_rPort_0_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_0_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_rPort_0_backpressure; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_rPort_0_output_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_3_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_3_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_wPort_3_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_wPort_3_data_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_wPort_3_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_2_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_2_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_wPort_2_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_wPort_2_data_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_wPort_2_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_1_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_1_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_wPort_1_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_wPort_1_data_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_wPort_1_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_0_banks_1; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [2:0] x398_lb_0_io_wPort_0_banks_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [8:0] x398_lb_0_io_wPort_0_ofs_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire [31:0] x398_lb_0_io_wPort_0_data_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x398_lb_0_io_wPort_0_en_0; // @[m_x398_lb_0.scala 47:17:@44849.4]
  wire  x403_1_clock; // @[Math.scala 366:24:@45032.4]
  wire [31:0] x403_1_io_a; // @[Math.scala 366:24:@45032.4]
  wire  x403_1_io_flow; // @[Math.scala 366:24:@45032.4]
  wire [31:0] x403_1_io_result; // @[Math.scala 366:24:@45032.4]
  wire  x713_sum_1_clock; // @[Math.scala 150:24:@45069.4]
  wire  x713_sum_1_reset; // @[Math.scala 150:24:@45069.4]
  wire [31:0] x713_sum_1_io_a; // @[Math.scala 150:24:@45069.4]
  wire [31:0] x713_sum_1_io_b; // @[Math.scala 150:24:@45069.4]
  wire  x713_sum_1_io_flow; // @[Math.scala 150:24:@45069.4]
  wire [31:0] x713_sum_1_io_result; // @[Math.scala 150:24:@45069.4]
  wire  x406_div_1_clock; // @[Math.scala 327:24:@45081.4]
  wire [31:0] x406_div_1_io_a; // @[Math.scala 327:24:@45081.4]
  wire  x406_div_1_io_flow; // @[Math.scala 327:24:@45081.4]
  wire [31:0] x406_div_1_io_result; // @[Math.scala 327:24:@45081.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45091.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45091.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45091.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@45091.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@45091.4]
  wire  x407_sum_1_clock; // @[Math.scala 150:24:@45100.4]
  wire  x407_sum_1_reset; // @[Math.scala 150:24:@45100.4]
  wire [31:0] x407_sum_1_io_a; // @[Math.scala 150:24:@45100.4]
  wire [31:0] x407_sum_1_io_b; // @[Math.scala 150:24:@45100.4]
  wire  x407_sum_1_io_flow; // @[Math.scala 150:24:@45100.4]
  wire [31:0] x407_sum_1_io_result; // @[Math.scala 150:24:@45100.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@45110.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@45110.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@45110.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@45110.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@45110.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@45119.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@45119.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@45119.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@45119.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@45119.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@45128.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@45128.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@45128.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@45128.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@45128.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@45137.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@45137.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@45137.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@45137.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@45137.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@45146.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@45146.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@45155.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@45155.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@45155.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@45155.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@45155.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@45166.4]
  wire  x409_rdcol_1_clock; // @[Math.scala 150:24:@45189.4]
  wire  x409_rdcol_1_reset; // @[Math.scala 150:24:@45189.4]
  wire [31:0] x409_rdcol_1_io_a; // @[Math.scala 150:24:@45189.4]
  wire [31:0] x409_rdcol_1_io_b; // @[Math.scala 150:24:@45189.4]
  wire  x409_rdcol_1_io_flow; // @[Math.scala 150:24:@45189.4]
  wire [31:0] x409_rdcol_1_io_result; // @[Math.scala 150:24:@45189.4]
  wire  x411_1_clock; // @[Math.scala 366:24:@45203.4]
  wire [31:0] x411_1_io_a; // @[Math.scala 366:24:@45203.4]
  wire  x411_1_io_flow; // @[Math.scala 366:24:@45203.4]
  wire [31:0] x411_1_io_result; // @[Math.scala 366:24:@45203.4]
  wire  x412_div_1_clock; // @[Math.scala 327:24:@45215.4]
  wire [31:0] x412_div_1_io_a; // @[Math.scala 327:24:@45215.4]
  wire  x412_div_1_io_flow; // @[Math.scala 327:24:@45215.4]
  wire [31:0] x412_div_1_io_result; // @[Math.scala 327:24:@45215.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@45225.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@45225.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@45225.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@45225.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@45225.4]
  wire  x413_sum_1_clock; // @[Math.scala 150:24:@45234.4]
  wire  x413_sum_1_reset; // @[Math.scala 150:24:@45234.4]
  wire [31:0] x413_sum_1_io_a; // @[Math.scala 150:24:@45234.4]
  wire [31:0] x413_sum_1_io_b; // @[Math.scala 150:24:@45234.4]
  wire  x413_sum_1_io_flow; // @[Math.scala 150:24:@45234.4]
  wire [31:0] x413_sum_1_io_result; // @[Math.scala 150:24:@45234.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@45244.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@45244.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@45244.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@45244.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@45244.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@45253.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@45253.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@45253.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@45253.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@45253.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@45262.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@45262.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@45262.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@45262.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@45262.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@45273.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@45273.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@45273.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@45273.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@45273.4]
  wire  x415_rdcol_1_clock; // @[Math.scala 150:24:@45296.4]
  wire  x415_rdcol_1_reset; // @[Math.scala 150:24:@45296.4]
  wire [31:0] x415_rdcol_1_io_a; // @[Math.scala 150:24:@45296.4]
  wire [31:0] x415_rdcol_1_io_b; // @[Math.scala 150:24:@45296.4]
  wire  x415_rdcol_1_io_flow; // @[Math.scala 150:24:@45296.4]
  wire [31:0] x415_rdcol_1_io_result; // @[Math.scala 150:24:@45296.4]
  wire  x417_1_clock; // @[Math.scala 366:24:@45310.4]
  wire [31:0] x417_1_io_a; // @[Math.scala 366:24:@45310.4]
  wire  x417_1_io_flow; // @[Math.scala 366:24:@45310.4]
  wire [31:0] x417_1_io_result; // @[Math.scala 366:24:@45310.4]
  wire  x418_div_1_clock; // @[Math.scala 327:24:@45322.4]
  wire [31:0] x418_div_1_io_a; // @[Math.scala 327:24:@45322.4]
  wire  x418_div_1_io_flow; // @[Math.scala 327:24:@45322.4]
  wire [31:0] x418_div_1_io_result; // @[Math.scala 327:24:@45322.4]
  wire  x419_sum_1_clock; // @[Math.scala 150:24:@45332.4]
  wire  x419_sum_1_reset; // @[Math.scala 150:24:@45332.4]
  wire [31:0] x419_sum_1_io_a; // @[Math.scala 150:24:@45332.4]
  wire [31:0] x419_sum_1_io_b; // @[Math.scala 150:24:@45332.4]
  wire  x419_sum_1_io_flow; // @[Math.scala 150:24:@45332.4]
  wire [31:0] x419_sum_1_io_result; // @[Math.scala 150:24:@45332.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@45342.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@45342.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@45342.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@45342.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@45342.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@45351.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@45351.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@45351.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@45351.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@45351.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@45360.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@45360.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@45360.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@45360.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@45360.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@45371.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@45371.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@45371.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@45371.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@45371.4]
  wire  x421_rdcol_1_clock; // @[Math.scala 150:24:@45394.4]
  wire  x421_rdcol_1_reset; // @[Math.scala 150:24:@45394.4]
  wire [31:0] x421_rdcol_1_io_a; // @[Math.scala 150:24:@45394.4]
  wire [31:0] x421_rdcol_1_io_b; // @[Math.scala 150:24:@45394.4]
  wire  x421_rdcol_1_io_flow; // @[Math.scala 150:24:@45394.4]
  wire [31:0] x421_rdcol_1_io_result; // @[Math.scala 150:24:@45394.4]
  wire  x423_1_clock; // @[Math.scala 366:24:@45408.4]
  wire [31:0] x423_1_io_a; // @[Math.scala 366:24:@45408.4]
  wire  x423_1_io_flow; // @[Math.scala 366:24:@45408.4]
  wire [31:0] x423_1_io_result; // @[Math.scala 366:24:@45408.4]
  wire  x424_div_1_clock; // @[Math.scala 327:24:@45420.4]
  wire [31:0] x424_div_1_io_a; // @[Math.scala 327:24:@45420.4]
  wire  x424_div_1_io_flow; // @[Math.scala 327:24:@45420.4]
  wire [31:0] x424_div_1_io_result; // @[Math.scala 327:24:@45420.4]
  wire  x425_sum_1_clock; // @[Math.scala 150:24:@45430.4]
  wire  x425_sum_1_reset; // @[Math.scala 150:24:@45430.4]
  wire [31:0] x425_sum_1_io_a; // @[Math.scala 150:24:@45430.4]
  wire [31:0] x425_sum_1_io_b; // @[Math.scala 150:24:@45430.4]
  wire  x425_sum_1_io_flow; // @[Math.scala 150:24:@45430.4]
  wire [31:0] x425_sum_1_io_result; // @[Math.scala 150:24:@45430.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@45440.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@45440.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@45440.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@45440.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@45440.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@45449.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@45449.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@45449.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@45449.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@45449.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@45458.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@45458.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@45458.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@45458.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@45458.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@45469.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@45469.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@45469.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@45469.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@45469.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@45490.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@45490.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@45490.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@45490.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@45490.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@45506.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@45506.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@45506.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@45506.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@45506.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@45515.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@45515.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@45515.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@45515.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@45515.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@45529.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@45529.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@45529.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@45529.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@45529.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@45538.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@45538.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@45538.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@45538.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@45538.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@45553.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@45553.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@45553.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@45553.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@45553.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@45562.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@45562.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@45562.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@45562.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@45562.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@45571.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@45571.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@45571.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@45571.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@45571.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@45580.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@45580.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@45580.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@45580.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@45580.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@45589.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@45589.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@45589.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@45589.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@45589.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@45598.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@45598.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@45598.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@45598.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@45598.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@45610.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@45610.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@45610.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@45610.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@45610.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@45631.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@45631.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@45645.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@45645.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@45645.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@45645.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@45645.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@45660.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@45660.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@45660.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@45660.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@45660.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@45669.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@45669.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@45669.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@45669.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@45669.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@45678.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@45678.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@45678.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@45678.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@45678.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@45690.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@45690.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@45690.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@45690.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@45690.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@45711.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@45711.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@45711.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@45711.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@45711.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@45725.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@45725.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@45725.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@45725.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@45725.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@45740.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@45740.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@45740.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@45740.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@45740.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@45749.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@45749.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@45749.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@45749.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@45749.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@45758.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@45758.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@45758.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@45758.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@45758.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@45770.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@45770.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@45770.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@45770.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@45770.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@45791.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@45791.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@45791.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@45791.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@45791.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@45805.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@45805.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@45805.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@45805.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@45805.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@45820.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@45820.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@45820.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@45820.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@45820.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@45829.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@45829.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@45829.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@45829.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@45829.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@45838.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@45838.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@45838.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@45838.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@45838.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@45850.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@45850.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@45850.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@45850.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@45850.4]
  wire  x449_rdcol_1_clock; // @[Math.scala 150:24:@45873.4]
  wire  x449_rdcol_1_reset; // @[Math.scala 150:24:@45873.4]
  wire [31:0] x449_rdcol_1_io_a; // @[Math.scala 150:24:@45873.4]
  wire [31:0] x449_rdcol_1_io_b; // @[Math.scala 150:24:@45873.4]
  wire  x449_rdcol_1_io_flow; // @[Math.scala 150:24:@45873.4]
  wire [31:0] x449_rdcol_1_io_result; // @[Math.scala 150:24:@45873.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@45888.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@45888.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@45888.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@45888.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@45888.4]
  wire  x453_1_clock; // @[Math.scala 366:24:@45907.4]
  wire [31:0] x453_1_io_a; // @[Math.scala 366:24:@45907.4]
  wire  x453_1_io_flow; // @[Math.scala 366:24:@45907.4]
  wire [31:0] x453_1_io_result; // @[Math.scala 366:24:@45907.4]
  wire  x454_div_1_clock; // @[Math.scala 327:24:@45919.4]
  wire [31:0] x454_div_1_io_a; // @[Math.scala 327:24:@45919.4]
  wire  x454_div_1_io_flow; // @[Math.scala 327:24:@45919.4]
  wire [31:0] x454_div_1_io_result; // @[Math.scala 327:24:@45919.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@45929.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@45929.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@45929.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@45929.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@45929.4]
  wire  x455_sum_1_clock; // @[Math.scala 150:24:@45938.4]
  wire  x455_sum_1_reset; // @[Math.scala 150:24:@45938.4]
  wire [31:0] x455_sum_1_io_a; // @[Math.scala 150:24:@45938.4]
  wire [31:0] x455_sum_1_io_b; // @[Math.scala 150:24:@45938.4]
  wire  x455_sum_1_io_flow; // @[Math.scala 150:24:@45938.4]
  wire [31:0] x455_sum_1_io_result; // @[Math.scala 150:24:@45938.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@45948.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@45948.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@45948.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@45948.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@45948.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@45957.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@45957.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@45957.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@45957.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@45957.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@45969.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@45969.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@45969.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@45969.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@45969.4]
  wire  x458_rdcol_1_clock; // @[Math.scala 150:24:@45992.4]
  wire  x458_rdcol_1_reset; // @[Math.scala 150:24:@45992.4]
  wire [31:0] x458_rdcol_1_io_a; // @[Math.scala 150:24:@45992.4]
  wire [31:0] x458_rdcol_1_io_b; // @[Math.scala 150:24:@45992.4]
  wire  x458_rdcol_1_io_flow; // @[Math.scala 150:24:@45992.4]
  wire [31:0] x458_rdcol_1_io_result; // @[Math.scala 150:24:@45992.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@46007.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@46007.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@46007.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@46007.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@46007.4]
  wire  x462_1_clock; // @[Math.scala 366:24:@46024.4]
  wire [31:0] x462_1_io_a; // @[Math.scala 366:24:@46024.4]
  wire  x462_1_io_flow; // @[Math.scala 366:24:@46024.4]
  wire [31:0] x462_1_io_result; // @[Math.scala 366:24:@46024.4]
  wire  x463_div_1_clock; // @[Math.scala 327:24:@46036.4]
  wire [31:0] x463_div_1_io_a; // @[Math.scala 327:24:@46036.4]
  wire  x463_div_1_io_flow; // @[Math.scala 327:24:@46036.4]
  wire [31:0] x463_div_1_io_result; // @[Math.scala 327:24:@46036.4]
  wire  x464_sum_1_clock; // @[Math.scala 150:24:@46046.4]
  wire  x464_sum_1_reset; // @[Math.scala 150:24:@46046.4]
  wire [31:0] x464_sum_1_io_a; // @[Math.scala 150:24:@46046.4]
  wire [31:0] x464_sum_1_io_b; // @[Math.scala 150:24:@46046.4]
  wire  x464_sum_1_io_flow; // @[Math.scala 150:24:@46046.4]
  wire [31:0] x464_sum_1_io_result; // @[Math.scala 150:24:@46046.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@46056.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@46056.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@46056.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@46056.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@46056.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@46065.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@46065.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@46065.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@46065.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@46065.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@46077.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@46077.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@46077.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@46077.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@46077.4]
  wire  x467_rdrow_1_clock; // @[Math.scala 191:24:@46100.4]
  wire  x467_rdrow_1_reset; // @[Math.scala 191:24:@46100.4]
  wire [31:0] x467_rdrow_1_io_a; // @[Math.scala 191:24:@46100.4]
  wire [31:0] x467_rdrow_1_io_b; // @[Math.scala 191:24:@46100.4]
  wire  x467_rdrow_1_io_flow; // @[Math.scala 191:24:@46100.4]
  wire [31:0] x467_rdrow_1_io_result; // @[Math.scala 191:24:@46100.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@46126.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@46126.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@46126.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@46126.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@46126.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@46148.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@46148.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@46148.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@46148.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@46148.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@46174.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@46174.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@46174.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@46174.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@46174.4]
  wire  x718_sum_1_clock; // @[Math.scala 150:24:@46195.4]
  wire  x718_sum_1_reset; // @[Math.scala 150:24:@46195.4]
  wire [31:0] x718_sum_1_io_a; // @[Math.scala 150:24:@46195.4]
  wire [31:0] x718_sum_1_io_b; // @[Math.scala 150:24:@46195.4]
  wire  x718_sum_1_io_flow; // @[Math.scala 150:24:@46195.4]
  wire [31:0] x718_sum_1_io_result; // @[Math.scala 150:24:@46195.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@46205.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@46205.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@46205.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@46205.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@46205.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@46214.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@46214.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@46214.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@46214.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@46214.4]
  wire  x475_sum_1_clock; // @[Math.scala 150:24:@46223.4]
  wire  x475_sum_1_reset; // @[Math.scala 150:24:@46223.4]
  wire [31:0] x475_sum_1_io_a; // @[Math.scala 150:24:@46223.4]
  wire [31:0] x475_sum_1_io_b; // @[Math.scala 150:24:@46223.4]
  wire  x475_sum_1_io_flow; // @[Math.scala 150:24:@46223.4]
  wire [31:0] x475_sum_1_io_result; // @[Math.scala 150:24:@46223.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@46233.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@46233.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@46233.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@46233.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@46233.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@46242.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@46242.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@46242.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@46242.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@46242.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@46254.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@46254.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@46254.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@46254.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@46254.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@46281.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@46281.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@46281.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@46281.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@46281.4]
  wire  x480_sum_1_clock; // @[Math.scala 150:24:@46290.4]
  wire  x480_sum_1_reset; // @[Math.scala 150:24:@46290.4]
  wire [31:0] x480_sum_1_io_a; // @[Math.scala 150:24:@46290.4]
  wire [31:0] x480_sum_1_io_b; // @[Math.scala 150:24:@46290.4]
  wire  x480_sum_1_io_flow; // @[Math.scala 150:24:@46290.4]
  wire [31:0] x480_sum_1_io_result; // @[Math.scala 150:24:@46290.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@46300.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@46300.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@46300.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@46300.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@46300.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@46339.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@46339.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@46339.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@46339.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@46339.4]
  wire  x485_sum_1_clock; // @[Math.scala 150:24:@46348.4]
  wire  x485_sum_1_reset; // @[Math.scala 150:24:@46348.4]
  wire [31:0] x485_sum_1_io_a; // @[Math.scala 150:24:@46348.4]
  wire [31:0] x485_sum_1_io_b; // @[Math.scala 150:24:@46348.4]
  wire  x485_sum_1_io_flow; // @[Math.scala 150:24:@46348.4]
  wire [31:0] x485_sum_1_io_result; // @[Math.scala 150:24:@46348.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@46358.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@46358.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@46358.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@46358.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@46358.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@46370.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@46370.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@46370.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@46370.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@46370.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@46391.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@46391.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@46391.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@46391.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@46391.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@46406.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@46406.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@46406.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@46406.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@46406.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@46415.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@46415.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@46415.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@46415.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@46415.4]
  wire  x490_sum_1_clock; // @[Math.scala 150:24:@46426.4]
  wire  x490_sum_1_reset; // @[Math.scala 150:24:@46426.4]
  wire [31:0] x490_sum_1_io_a; // @[Math.scala 150:24:@46426.4]
  wire [31:0] x490_sum_1_io_b; // @[Math.scala 150:24:@46426.4]
  wire  x490_sum_1_io_flow; // @[Math.scala 150:24:@46426.4]
  wire [31:0] x490_sum_1_io_result; // @[Math.scala 150:24:@46426.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@46436.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@46436.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@46436.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@46436.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@46436.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@46445.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@46445.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@46445.4]
  wire [31:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@46445.4]
  wire [31:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@46445.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@46457.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@46457.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@46457.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@46457.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@46457.4]
  wire  x495_sum_1_clock; // @[Math.scala 150:24:@46484.4]
  wire  x495_sum_1_reset; // @[Math.scala 150:24:@46484.4]
  wire [31:0] x495_sum_1_io_a; // @[Math.scala 150:24:@46484.4]
  wire [31:0] x495_sum_1_io_b; // @[Math.scala 150:24:@46484.4]
  wire  x495_sum_1_io_flow; // @[Math.scala 150:24:@46484.4]
  wire [31:0] x495_sum_1_io_result; // @[Math.scala 150:24:@46484.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@46494.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@46494.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@46494.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@46494.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@46494.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@46506.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@46506.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@46506.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@46506.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@46506.4]
  wire  x500_sum_1_clock; // @[Math.scala 150:24:@46533.4]
  wire  x500_sum_1_reset; // @[Math.scala 150:24:@46533.4]
  wire [31:0] x500_sum_1_io_a; // @[Math.scala 150:24:@46533.4]
  wire [31:0] x500_sum_1_io_b; // @[Math.scala 150:24:@46533.4]
  wire  x500_sum_1_io_flow; // @[Math.scala 150:24:@46533.4]
  wire [31:0] x500_sum_1_io_result; // @[Math.scala 150:24:@46533.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@46543.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@46543.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@46543.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@46543.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@46543.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@46555.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@46555.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@46555.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@46555.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@46555.4]
  wire  x503_rdrow_1_clock; // @[Math.scala 191:24:@46578.4]
  wire  x503_rdrow_1_reset; // @[Math.scala 191:24:@46578.4]
  wire [31:0] x503_rdrow_1_io_a; // @[Math.scala 191:24:@46578.4]
  wire [31:0] x503_rdrow_1_io_b; // @[Math.scala 191:24:@46578.4]
  wire  x503_rdrow_1_io_flow; // @[Math.scala 191:24:@46578.4]
  wire [31:0] x503_rdrow_1_io_result; // @[Math.scala 191:24:@46578.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@46604.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@46604.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@46604.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@46604.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@46604.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@46626.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@46626.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@46626.4]
  wire [31:0] RetimeWrapper_86_io_in; // @[package.scala 93:22:@46626.4]
  wire [31:0] RetimeWrapper_86_io_out; // @[package.scala 93:22:@46626.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@46652.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@46652.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@46652.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@46652.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@46652.4]
  wire  x723_sum_1_clock; // @[Math.scala 150:24:@46673.4]
  wire  x723_sum_1_reset; // @[Math.scala 150:24:@46673.4]
  wire [31:0] x723_sum_1_io_a; // @[Math.scala 150:24:@46673.4]
  wire [31:0] x723_sum_1_io_b; // @[Math.scala 150:24:@46673.4]
  wire  x723_sum_1_io_flow; // @[Math.scala 150:24:@46673.4]
  wire [31:0] x723_sum_1_io_result; // @[Math.scala 150:24:@46673.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@46683.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@46683.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@46683.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@46683.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@46683.4]
  wire  x511_sum_1_clock; // @[Math.scala 150:24:@46692.4]
  wire  x511_sum_1_reset; // @[Math.scala 150:24:@46692.4]
  wire [31:0] x511_sum_1_io_a; // @[Math.scala 150:24:@46692.4]
  wire [31:0] x511_sum_1_io_b; // @[Math.scala 150:24:@46692.4]
  wire  x511_sum_1_io_flow; // @[Math.scala 150:24:@46692.4]
  wire [31:0] x511_sum_1_io_result; // @[Math.scala 150:24:@46692.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@46702.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@46702.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@46702.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@46702.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@46702.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@46711.4]
  wire [31:0] RetimeWrapper_90_io_in; // @[package.scala 93:22:@46711.4]
  wire [31:0] RetimeWrapper_90_io_out; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@46723.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@46723.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@46723.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@46723.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@46723.4]
  wire  x516_sum_1_clock; // @[Math.scala 150:24:@46750.4]
  wire  x516_sum_1_reset; // @[Math.scala 150:24:@46750.4]
  wire [31:0] x516_sum_1_io_a; // @[Math.scala 150:24:@46750.4]
  wire [31:0] x516_sum_1_io_b; // @[Math.scala 150:24:@46750.4]
  wire  x516_sum_1_io_flow; // @[Math.scala 150:24:@46750.4]
  wire [31:0] x516_sum_1_io_result; // @[Math.scala 150:24:@46750.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@46760.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@46760.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@46760.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@46760.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@46760.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@46772.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@46772.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@46772.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@46772.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@46772.4]
  wire  x521_sum_1_clock; // @[Math.scala 150:24:@46799.4]
  wire  x521_sum_1_reset; // @[Math.scala 150:24:@46799.4]
  wire [31:0] x521_sum_1_io_a; // @[Math.scala 150:24:@46799.4]
  wire [31:0] x521_sum_1_io_b; // @[Math.scala 150:24:@46799.4]
  wire  x521_sum_1_io_flow; // @[Math.scala 150:24:@46799.4]
  wire [31:0] x521_sum_1_io_result; // @[Math.scala 150:24:@46799.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@46809.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@46809.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@46809.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@46809.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@46809.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@46848.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@46848.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@46848.4]
  wire [31:0] RetimeWrapper_96_io_in; // @[package.scala 93:22:@46848.4]
  wire [31:0] RetimeWrapper_96_io_out; // @[package.scala 93:22:@46848.4]
  wire  x526_sum_1_clock; // @[Math.scala 150:24:@46859.4]
  wire  x526_sum_1_reset; // @[Math.scala 150:24:@46859.4]
  wire [31:0] x526_sum_1_io_a; // @[Math.scala 150:24:@46859.4]
  wire [31:0] x526_sum_1_io_b; // @[Math.scala 150:24:@46859.4]
  wire  x526_sum_1_io_flow; // @[Math.scala 150:24:@46859.4]
  wire [31:0] x526_sum_1_io_result; // @[Math.scala 150:24:@46859.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@46869.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@46869.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@46869.4]
  wire [31:0] RetimeWrapper_97_io_in; // @[package.scala 93:22:@46869.4]
  wire [31:0] RetimeWrapper_97_io_out; // @[package.scala 93:22:@46869.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@46878.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@46878.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@46878.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@46878.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@46878.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@46890.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@46890.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@46890.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@46890.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@46890.4]
  wire  x531_sum_1_clock; // @[Math.scala 150:24:@46917.4]
  wire  x531_sum_1_reset; // @[Math.scala 150:24:@46917.4]
  wire [31:0] x531_sum_1_io_a; // @[Math.scala 150:24:@46917.4]
  wire [31:0] x531_sum_1_io_b; // @[Math.scala 150:24:@46917.4]
  wire  x531_sum_1_io_flow; // @[Math.scala 150:24:@46917.4]
  wire [31:0] x531_sum_1_io_result; // @[Math.scala 150:24:@46917.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@46927.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@46927.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@46927.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@46927.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@46927.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@46939.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@46939.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@46939.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@46939.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@46939.4]
  wire  x536_sum_1_clock; // @[Math.scala 150:24:@46966.4]
  wire  x536_sum_1_reset; // @[Math.scala 150:24:@46966.4]
  wire [31:0] x536_sum_1_io_a; // @[Math.scala 150:24:@46966.4]
  wire [31:0] x536_sum_1_io_b; // @[Math.scala 150:24:@46966.4]
  wire  x536_sum_1_io_flow; // @[Math.scala 150:24:@46966.4]
  wire [31:0] x536_sum_1_io_result; // @[Math.scala 150:24:@46966.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@46976.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@46976.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@46976.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@46976.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@46976.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@46988.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@46988.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@46988.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@46988.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@46988.4]
  wire  x544_x13_1_clock; // @[Math.scala 150:24:@47034.4]
  wire  x544_x13_1_reset; // @[Math.scala 150:24:@47034.4]
  wire [31:0] x544_x13_1_io_a; // @[Math.scala 150:24:@47034.4]
  wire [31:0] x544_x13_1_io_b; // @[Math.scala 150:24:@47034.4]
  wire  x544_x13_1_io_flow; // @[Math.scala 150:24:@47034.4]
  wire [31:0] x544_x13_1_io_result; // @[Math.scala 150:24:@47034.4]
  wire  x545_x14_1_clock; // @[Math.scala 150:24:@47044.4]
  wire  x545_x14_1_reset; // @[Math.scala 150:24:@47044.4]
  wire [31:0] x545_x14_1_io_a; // @[Math.scala 150:24:@47044.4]
  wire [31:0] x545_x14_1_io_b; // @[Math.scala 150:24:@47044.4]
  wire  x545_x14_1_io_flow; // @[Math.scala 150:24:@47044.4]
  wire [31:0] x545_x14_1_io_result; // @[Math.scala 150:24:@47044.4]
  wire  x546_x13_1_clock; // @[Math.scala 150:24:@47054.4]
  wire  x546_x13_1_reset; // @[Math.scala 150:24:@47054.4]
  wire [31:0] x546_x13_1_io_a; // @[Math.scala 150:24:@47054.4]
  wire [31:0] x546_x13_1_io_b; // @[Math.scala 150:24:@47054.4]
  wire  x546_x13_1_io_flow; // @[Math.scala 150:24:@47054.4]
  wire [31:0] x546_x13_1_io_result; // @[Math.scala 150:24:@47054.4]
  wire  x547_x14_1_clock; // @[Math.scala 150:24:@47064.4]
  wire  x547_x14_1_reset; // @[Math.scala 150:24:@47064.4]
  wire [31:0] x547_x14_1_io_a; // @[Math.scala 150:24:@47064.4]
  wire [31:0] x547_x14_1_io_b; // @[Math.scala 150:24:@47064.4]
  wire  x547_x14_1_io_flow; // @[Math.scala 150:24:@47064.4]
  wire [31:0] x547_x14_1_io_result; // @[Math.scala 150:24:@47064.4]
  wire  x548_x13_1_clock; // @[Math.scala 150:24:@47074.4]
  wire  x548_x13_1_reset; // @[Math.scala 150:24:@47074.4]
  wire [31:0] x548_x13_1_io_a; // @[Math.scala 150:24:@47074.4]
  wire [31:0] x548_x13_1_io_b; // @[Math.scala 150:24:@47074.4]
  wire  x548_x13_1_io_flow; // @[Math.scala 150:24:@47074.4]
  wire [31:0] x548_x13_1_io_result; // @[Math.scala 150:24:@47074.4]
  wire  x549_x14_1_clock; // @[Math.scala 150:24:@47084.4]
  wire  x549_x14_1_reset; // @[Math.scala 150:24:@47084.4]
  wire [31:0] x549_x14_1_io_a; // @[Math.scala 150:24:@47084.4]
  wire [31:0] x549_x14_1_io_b; // @[Math.scala 150:24:@47084.4]
  wire  x549_x14_1_io_flow; // @[Math.scala 150:24:@47084.4]
  wire [31:0] x549_x14_1_io_result; // @[Math.scala 150:24:@47084.4]
  wire  x550_x13_1_clock; // @[Math.scala 150:24:@47094.4]
  wire  x550_x13_1_reset; // @[Math.scala 150:24:@47094.4]
  wire [31:0] x550_x13_1_io_a; // @[Math.scala 150:24:@47094.4]
  wire [31:0] x550_x13_1_io_b; // @[Math.scala 150:24:@47094.4]
  wire  x550_x13_1_io_flow; // @[Math.scala 150:24:@47094.4]
  wire [31:0] x550_x13_1_io_result; // @[Math.scala 150:24:@47094.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@47104.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@47104.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@47104.4]
  wire [31:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@47104.4]
  wire [31:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@47104.4]
  wire  x551_sum_1_clock; // @[Math.scala 150:24:@47113.4]
  wire  x551_sum_1_reset; // @[Math.scala 150:24:@47113.4]
  wire [31:0] x551_sum_1_io_a; // @[Math.scala 150:24:@47113.4]
  wire [31:0] x551_sum_1_io_b; // @[Math.scala 150:24:@47113.4]
  wire  x551_sum_1_io_flow; // @[Math.scala 150:24:@47113.4]
  wire [31:0] x551_sum_1_io_result; // @[Math.scala 150:24:@47113.4]
  wire [31:0] x552_1_io_b; // @[Math.scala 720:24:@47123.4]
  wire [31:0] x552_1_io_result; // @[Math.scala 720:24:@47123.4]
  wire  x553_mul_1_clock; // @[Math.scala 262:24:@47134.4]
  wire [31:0] x553_mul_1_io_a; // @[Math.scala 262:24:@47134.4]
  wire [31:0] x553_mul_1_io_b; // @[Math.scala 262:24:@47134.4]
  wire  x553_mul_1_io_flow; // @[Math.scala 262:24:@47134.4]
  wire [31:0] x553_mul_1_io_result; // @[Math.scala 262:24:@47134.4]
  wire [31:0] x554_1_io_b; // @[Math.scala 720:24:@47144.4]
  wire [31:0] x554_1_io_result; // @[Math.scala 720:24:@47144.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@47153.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@47153.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@47153.4]
  wire [31:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@47153.4]
  wire [31:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@47153.4]
  wire  x555_sub_1_clock; // @[Math.scala 191:24:@47162.4]
  wire  x555_sub_1_reset; // @[Math.scala 191:24:@47162.4]
  wire [31:0] x555_sub_1_io_a; // @[Math.scala 191:24:@47162.4]
  wire [31:0] x555_sub_1_io_b; // @[Math.scala 191:24:@47162.4]
  wire  x555_sub_1_io_flow; // @[Math.scala 191:24:@47162.4]
  wire [31:0] x555_sub_1_io_result; // @[Math.scala 191:24:@47162.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@47175.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@47175.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@47175.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@47175.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@47175.4]
  wire  x557_sub_1_clock; // @[Math.scala 191:24:@47184.4]
  wire  x557_sub_1_reset; // @[Math.scala 191:24:@47184.4]
  wire [31:0] x557_sub_1_io_a; // @[Math.scala 191:24:@47184.4]
  wire [31:0] x557_sub_1_io_b; // @[Math.scala 191:24:@47184.4]
  wire  x557_sub_1_io_flow; // @[Math.scala 191:24:@47184.4]
  wire [31:0] x557_sub_1_io_result; // @[Math.scala 191:24:@47184.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@47197.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@47197.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@47197.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@47197.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@47197.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@47209.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@47209.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@47209.4]
  wire [31:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@47209.4]
  wire [31:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@47209.4]
  wire [31:0] x561_1_io_b; // @[Math.scala 720:24:@47223.4]
  wire [31:0] x561_1_io_result; // @[Math.scala 720:24:@47223.4]
  wire  x562_mul_1_clock; // @[Math.scala 262:24:@47234.4]
  wire [31:0] x562_mul_1_io_a; // @[Math.scala 262:24:@47234.4]
  wire [31:0] x562_mul_1_io_b; // @[Math.scala 262:24:@47234.4]
  wire  x562_mul_1_io_flow; // @[Math.scala 262:24:@47234.4]
  wire [31:0] x562_mul_1_io_result; // @[Math.scala 262:24:@47234.4]
  wire [31:0] x563_1_io_b; // @[Math.scala 720:24:@47246.4]
  wire [31:0] x563_1_io_result; // @[Math.scala 720:24:@47246.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@47255.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@47255.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@47255.4]
  wire [31:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@47255.4]
  wire [31:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@47255.4]
  wire  x564_sum_1_clock; // @[Math.scala 150:24:@47264.4]
  wire  x564_sum_1_reset; // @[Math.scala 150:24:@47264.4]
  wire [31:0] x564_sum_1_io_a; // @[Math.scala 150:24:@47264.4]
  wire [31:0] x564_sum_1_io_b; // @[Math.scala 150:24:@47264.4]
  wire  x564_sum_1_io_flow; // @[Math.scala 150:24:@47264.4]
  wire [31:0] x564_sum_1_io_result; // @[Math.scala 150:24:@47264.4]
  wire  x570_x13_1_clock; // @[Math.scala 150:24:@47299.4]
  wire  x570_x13_1_reset; // @[Math.scala 150:24:@47299.4]
  wire [31:0] x570_x13_1_io_a; // @[Math.scala 150:24:@47299.4]
  wire [31:0] x570_x13_1_io_b; // @[Math.scala 150:24:@47299.4]
  wire  x570_x13_1_io_flow; // @[Math.scala 150:24:@47299.4]
  wire [31:0] x570_x13_1_io_result; // @[Math.scala 150:24:@47299.4]
  wire  x571_x14_1_clock; // @[Math.scala 150:24:@47309.4]
  wire  x571_x14_1_reset; // @[Math.scala 150:24:@47309.4]
  wire [31:0] x571_x14_1_io_a; // @[Math.scala 150:24:@47309.4]
  wire [31:0] x571_x14_1_io_b; // @[Math.scala 150:24:@47309.4]
  wire  x571_x14_1_io_flow; // @[Math.scala 150:24:@47309.4]
  wire [31:0] x571_x14_1_io_result; // @[Math.scala 150:24:@47309.4]
  wire  x572_x13_1_clock; // @[Math.scala 150:24:@47319.4]
  wire  x572_x13_1_reset; // @[Math.scala 150:24:@47319.4]
  wire [31:0] x572_x13_1_io_a; // @[Math.scala 150:24:@47319.4]
  wire [31:0] x572_x13_1_io_b; // @[Math.scala 150:24:@47319.4]
  wire  x572_x13_1_io_flow; // @[Math.scala 150:24:@47319.4]
  wire [31:0] x572_x13_1_io_result; // @[Math.scala 150:24:@47319.4]
  wire  x573_x14_1_clock; // @[Math.scala 150:24:@47329.4]
  wire  x573_x14_1_reset; // @[Math.scala 150:24:@47329.4]
  wire [31:0] x573_x14_1_io_a; // @[Math.scala 150:24:@47329.4]
  wire [31:0] x573_x14_1_io_b; // @[Math.scala 150:24:@47329.4]
  wire  x573_x14_1_io_flow; // @[Math.scala 150:24:@47329.4]
  wire [31:0] x573_x14_1_io_result; // @[Math.scala 150:24:@47329.4]
  wire  x574_x13_1_clock; // @[Math.scala 150:24:@47339.4]
  wire  x574_x13_1_reset; // @[Math.scala 150:24:@47339.4]
  wire [31:0] x574_x13_1_io_a; // @[Math.scala 150:24:@47339.4]
  wire [31:0] x574_x13_1_io_b; // @[Math.scala 150:24:@47339.4]
  wire  x574_x13_1_io_flow; // @[Math.scala 150:24:@47339.4]
  wire [31:0] x574_x13_1_io_result; // @[Math.scala 150:24:@47339.4]
  wire  x575_x14_1_clock; // @[Math.scala 150:24:@47349.4]
  wire  x575_x14_1_reset; // @[Math.scala 150:24:@47349.4]
  wire [31:0] x575_x14_1_io_a; // @[Math.scala 150:24:@47349.4]
  wire [31:0] x575_x14_1_io_b; // @[Math.scala 150:24:@47349.4]
  wire  x575_x14_1_io_flow; // @[Math.scala 150:24:@47349.4]
  wire [31:0] x575_x14_1_io_result; // @[Math.scala 150:24:@47349.4]
  wire  x576_x13_1_clock; // @[Math.scala 150:24:@47359.4]
  wire  x576_x13_1_reset; // @[Math.scala 150:24:@47359.4]
  wire [31:0] x576_x13_1_io_a; // @[Math.scala 150:24:@47359.4]
  wire [31:0] x576_x13_1_io_b; // @[Math.scala 150:24:@47359.4]
  wire  x576_x13_1_io_flow; // @[Math.scala 150:24:@47359.4]
  wire [31:0] x576_x13_1_io_result; // @[Math.scala 150:24:@47359.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@47369.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@47369.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@47369.4]
  wire [31:0] RetimeWrapper_110_io_in; // @[package.scala 93:22:@47369.4]
  wire [31:0] RetimeWrapper_110_io_out; // @[package.scala 93:22:@47369.4]
  wire  x577_sum_1_clock; // @[Math.scala 150:24:@47378.4]
  wire  x577_sum_1_reset; // @[Math.scala 150:24:@47378.4]
  wire [31:0] x577_sum_1_io_a; // @[Math.scala 150:24:@47378.4]
  wire [31:0] x577_sum_1_io_b; // @[Math.scala 150:24:@47378.4]
  wire  x577_sum_1_io_flow; // @[Math.scala 150:24:@47378.4]
  wire [31:0] x577_sum_1_io_result; // @[Math.scala 150:24:@47378.4]
  wire [31:0] x578_1_io_b; // @[Math.scala 720:24:@47388.4]
  wire [31:0] x578_1_io_result; // @[Math.scala 720:24:@47388.4]
  wire  x579_mul_1_clock; // @[Math.scala 262:24:@47399.4]
  wire [31:0] x579_mul_1_io_a; // @[Math.scala 262:24:@47399.4]
  wire [31:0] x579_mul_1_io_b; // @[Math.scala 262:24:@47399.4]
  wire  x579_mul_1_io_flow; // @[Math.scala 262:24:@47399.4]
  wire [31:0] x579_mul_1_io_result; // @[Math.scala 262:24:@47399.4]
  wire [31:0] x580_1_io_b; // @[Math.scala 720:24:@47409.4]
  wire [31:0] x580_1_io_result; // @[Math.scala 720:24:@47409.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@47418.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@47418.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@47418.4]
  wire [31:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@47418.4]
  wire [31:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@47418.4]
  wire  x581_sub_1_clock; // @[Math.scala 191:24:@47427.4]
  wire  x581_sub_1_reset; // @[Math.scala 191:24:@47427.4]
  wire [31:0] x581_sub_1_io_a; // @[Math.scala 191:24:@47427.4]
  wire [31:0] x581_sub_1_io_b; // @[Math.scala 191:24:@47427.4]
  wire  x581_sub_1_io_flow; // @[Math.scala 191:24:@47427.4]
  wire [31:0] x581_sub_1_io_result; // @[Math.scala 191:24:@47427.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@47440.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@47440.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@47440.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@47440.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@47440.4]
  wire  x583_sub_1_clock; // @[Math.scala 191:24:@47449.4]
  wire  x583_sub_1_reset; // @[Math.scala 191:24:@47449.4]
  wire [31:0] x583_sub_1_io_a; // @[Math.scala 191:24:@47449.4]
  wire [31:0] x583_sub_1_io_b; // @[Math.scala 191:24:@47449.4]
  wire  x583_sub_1_io_flow; // @[Math.scala 191:24:@47449.4]
  wire [31:0] x583_sub_1_io_result; // @[Math.scala 191:24:@47449.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@47462.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@47462.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@47462.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@47462.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@47462.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@47474.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@47474.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@47474.4]
  wire [31:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@47474.4]
  wire [31:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@47474.4]
  wire [31:0] x587_1_io_b; // @[Math.scala 720:24:@47488.4]
  wire [31:0] x587_1_io_result; // @[Math.scala 720:24:@47488.4]
  wire  x588_mul_1_clock; // @[Math.scala 262:24:@47499.4]
  wire [31:0] x588_mul_1_io_a; // @[Math.scala 262:24:@47499.4]
  wire [31:0] x588_mul_1_io_b; // @[Math.scala 262:24:@47499.4]
  wire  x588_mul_1_io_flow; // @[Math.scala 262:24:@47499.4]
  wire [31:0] x588_mul_1_io_result; // @[Math.scala 262:24:@47499.4]
  wire [31:0] x589_1_io_b; // @[Math.scala 720:24:@47509.4]
  wire [31:0] x589_1_io_result; // @[Math.scala 720:24:@47509.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@47518.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@47518.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@47518.4]
  wire [31:0] RetimeWrapper_115_io_in; // @[package.scala 93:22:@47518.4]
  wire [31:0] RetimeWrapper_115_io_out; // @[package.scala 93:22:@47518.4]
  wire  x590_sum_1_clock; // @[Math.scala 150:24:@47527.4]
  wire  x590_sum_1_reset; // @[Math.scala 150:24:@47527.4]
  wire [31:0] x590_sum_1_io_a; // @[Math.scala 150:24:@47527.4]
  wire [31:0] x590_sum_1_io_b; // @[Math.scala 150:24:@47527.4]
  wire  x590_sum_1_io_flow; // @[Math.scala 150:24:@47527.4]
  wire [31:0] x590_sum_1_io_result; // @[Math.scala 150:24:@47527.4]
  wire  x595_x13_1_clock; // @[Math.scala 150:24:@47557.4]
  wire  x595_x13_1_reset; // @[Math.scala 150:24:@47557.4]
  wire [31:0] x595_x13_1_io_a; // @[Math.scala 150:24:@47557.4]
  wire [31:0] x595_x13_1_io_b; // @[Math.scala 150:24:@47557.4]
  wire  x595_x13_1_io_flow; // @[Math.scala 150:24:@47557.4]
  wire [31:0] x595_x13_1_io_result; // @[Math.scala 150:24:@47557.4]
  wire  x596_x14_1_clock; // @[Math.scala 150:24:@47567.4]
  wire  x596_x14_1_reset; // @[Math.scala 150:24:@47567.4]
  wire [31:0] x596_x14_1_io_a; // @[Math.scala 150:24:@47567.4]
  wire [31:0] x596_x14_1_io_b; // @[Math.scala 150:24:@47567.4]
  wire  x596_x14_1_io_flow; // @[Math.scala 150:24:@47567.4]
  wire [31:0] x596_x14_1_io_result; // @[Math.scala 150:24:@47567.4]
  wire  x597_x13_1_clock; // @[Math.scala 150:24:@47577.4]
  wire  x597_x13_1_reset; // @[Math.scala 150:24:@47577.4]
  wire [31:0] x597_x13_1_io_a; // @[Math.scala 150:24:@47577.4]
  wire [31:0] x597_x13_1_io_b; // @[Math.scala 150:24:@47577.4]
  wire  x597_x13_1_io_flow; // @[Math.scala 150:24:@47577.4]
  wire [31:0] x597_x13_1_io_result; // @[Math.scala 150:24:@47577.4]
  wire  x598_x14_1_clock; // @[Math.scala 150:24:@47587.4]
  wire  x598_x14_1_reset; // @[Math.scala 150:24:@47587.4]
  wire [31:0] x598_x14_1_io_a; // @[Math.scala 150:24:@47587.4]
  wire [31:0] x598_x14_1_io_b; // @[Math.scala 150:24:@47587.4]
  wire  x598_x14_1_io_flow; // @[Math.scala 150:24:@47587.4]
  wire [31:0] x598_x14_1_io_result; // @[Math.scala 150:24:@47587.4]
  wire  x599_x13_1_clock; // @[Math.scala 150:24:@47597.4]
  wire  x599_x13_1_reset; // @[Math.scala 150:24:@47597.4]
  wire [31:0] x599_x13_1_io_a; // @[Math.scala 150:24:@47597.4]
  wire [31:0] x599_x13_1_io_b; // @[Math.scala 150:24:@47597.4]
  wire  x599_x13_1_io_flow; // @[Math.scala 150:24:@47597.4]
  wire [31:0] x599_x13_1_io_result; // @[Math.scala 150:24:@47597.4]
  wire  x600_x14_1_clock; // @[Math.scala 150:24:@47607.4]
  wire  x600_x14_1_reset; // @[Math.scala 150:24:@47607.4]
  wire [31:0] x600_x14_1_io_a; // @[Math.scala 150:24:@47607.4]
  wire [31:0] x600_x14_1_io_b; // @[Math.scala 150:24:@47607.4]
  wire  x600_x14_1_io_flow; // @[Math.scala 150:24:@47607.4]
  wire [31:0] x600_x14_1_io_result; // @[Math.scala 150:24:@47607.4]
  wire  x601_x13_1_clock; // @[Math.scala 150:24:@47617.4]
  wire  x601_x13_1_reset; // @[Math.scala 150:24:@47617.4]
  wire [31:0] x601_x13_1_io_a; // @[Math.scala 150:24:@47617.4]
  wire [31:0] x601_x13_1_io_b; // @[Math.scala 150:24:@47617.4]
  wire  x601_x13_1_io_flow; // @[Math.scala 150:24:@47617.4]
  wire [31:0] x601_x13_1_io_result; // @[Math.scala 150:24:@47617.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@47627.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@47627.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@47627.4]
  wire [31:0] RetimeWrapper_116_io_in; // @[package.scala 93:22:@47627.4]
  wire [31:0] RetimeWrapper_116_io_out; // @[package.scala 93:22:@47627.4]
  wire  x602_sum_1_clock; // @[Math.scala 150:24:@47636.4]
  wire  x602_sum_1_reset; // @[Math.scala 150:24:@47636.4]
  wire [31:0] x602_sum_1_io_a; // @[Math.scala 150:24:@47636.4]
  wire [31:0] x602_sum_1_io_b; // @[Math.scala 150:24:@47636.4]
  wire  x602_sum_1_io_flow; // @[Math.scala 150:24:@47636.4]
  wire [31:0] x602_sum_1_io_result; // @[Math.scala 150:24:@47636.4]
  wire [31:0] x603_1_io_b; // @[Math.scala 720:24:@47646.4]
  wire [31:0] x603_1_io_result; // @[Math.scala 720:24:@47646.4]
  wire  x604_mul_1_clock; // @[Math.scala 262:24:@47657.4]
  wire [31:0] x604_mul_1_io_a; // @[Math.scala 262:24:@47657.4]
  wire [31:0] x604_mul_1_io_b; // @[Math.scala 262:24:@47657.4]
  wire  x604_mul_1_io_flow; // @[Math.scala 262:24:@47657.4]
  wire [31:0] x604_mul_1_io_result; // @[Math.scala 262:24:@47657.4]
  wire [31:0] x605_1_io_b; // @[Math.scala 720:24:@47667.4]
  wire [31:0] x605_1_io_result; // @[Math.scala 720:24:@47667.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@47676.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@47676.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@47676.4]
  wire [31:0] RetimeWrapper_117_io_in; // @[package.scala 93:22:@47676.4]
  wire [31:0] RetimeWrapper_117_io_out; // @[package.scala 93:22:@47676.4]
  wire  x606_sub_1_clock; // @[Math.scala 191:24:@47687.4]
  wire  x606_sub_1_reset; // @[Math.scala 191:24:@47687.4]
  wire [31:0] x606_sub_1_io_a; // @[Math.scala 191:24:@47687.4]
  wire [31:0] x606_sub_1_io_b; // @[Math.scala 191:24:@47687.4]
  wire  x606_sub_1_io_flow; // @[Math.scala 191:24:@47687.4]
  wire [31:0] x606_sub_1_io_result; // @[Math.scala 191:24:@47687.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@47700.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@47700.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@47700.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@47700.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@47700.4]
  wire  x608_sub_1_clock; // @[Math.scala 191:24:@47709.4]
  wire  x608_sub_1_reset; // @[Math.scala 191:24:@47709.4]
  wire [31:0] x608_sub_1_io_a; // @[Math.scala 191:24:@47709.4]
  wire [31:0] x608_sub_1_io_b; // @[Math.scala 191:24:@47709.4]
  wire  x608_sub_1_io_flow; // @[Math.scala 191:24:@47709.4]
  wire [31:0] x608_sub_1_io_result; // @[Math.scala 191:24:@47709.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@47722.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@47722.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@47722.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@47722.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@47722.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@47734.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@47734.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@47734.4]
  wire [31:0] RetimeWrapper_120_io_in; // @[package.scala 93:22:@47734.4]
  wire [31:0] RetimeWrapper_120_io_out; // @[package.scala 93:22:@47734.4]
  wire [31:0] x612_1_io_b; // @[Math.scala 720:24:@47748.4]
  wire [31:0] x612_1_io_result; // @[Math.scala 720:24:@47748.4]
  wire  x613_mul_1_clock; // @[Math.scala 262:24:@47759.4]
  wire [31:0] x613_mul_1_io_a; // @[Math.scala 262:24:@47759.4]
  wire [31:0] x613_mul_1_io_b; // @[Math.scala 262:24:@47759.4]
  wire  x613_mul_1_io_flow; // @[Math.scala 262:24:@47759.4]
  wire [31:0] x613_mul_1_io_result; // @[Math.scala 262:24:@47759.4]
  wire [31:0] x614_1_io_b; // @[Math.scala 720:24:@47769.4]
  wire [31:0] x614_1_io_result; // @[Math.scala 720:24:@47769.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@47778.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@47778.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@47778.4]
  wire [31:0] RetimeWrapper_121_io_in; // @[package.scala 93:22:@47778.4]
  wire [31:0] RetimeWrapper_121_io_out; // @[package.scala 93:22:@47778.4]
  wire  x615_sum_1_clock; // @[Math.scala 150:24:@47787.4]
  wire  x615_sum_1_reset; // @[Math.scala 150:24:@47787.4]
  wire [31:0] x615_sum_1_io_a; // @[Math.scala 150:24:@47787.4]
  wire [31:0] x615_sum_1_io_b; // @[Math.scala 150:24:@47787.4]
  wire  x615_sum_1_io_flow; // @[Math.scala 150:24:@47787.4]
  wire [31:0] x615_sum_1_io_result; // @[Math.scala 150:24:@47787.4]
  wire  x620_x13_1_clock; // @[Math.scala 150:24:@47817.4]
  wire  x620_x13_1_reset; // @[Math.scala 150:24:@47817.4]
  wire [31:0] x620_x13_1_io_a; // @[Math.scala 150:24:@47817.4]
  wire [31:0] x620_x13_1_io_b; // @[Math.scala 150:24:@47817.4]
  wire  x620_x13_1_io_flow; // @[Math.scala 150:24:@47817.4]
  wire [31:0] x620_x13_1_io_result; // @[Math.scala 150:24:@47817.4]
  wire  x621_x14_1_clock; // @[Math.scala 150:24:@47827.4]
  wire  x621_x14_1_reset; // @[Math.scala 150:24:@47827.4]
  wire [31:0] x621_x14_1_io_a; // @[Math.scala 150:24:@47827.4]
  wire [31:0] x621_x14_1_io_b; // @[Math.scala 150:24:@47827.4]
  wire  x621_x14_1_io_flow; // @[Math.scala 150:24:@47827.4]
  wire [31:0] x621_x14_1_io_result; // @[Math.scala 150:24:@47827.4]
  wire  x622_x13_1_clock; // @[Math.scala 150:24:@47837.4]
  wire  x622_x13_1_reset; // @[Math.scala 150:24:@47837.4]
  wire [31:0] x622_x13_1_io_a; // @[Math.scala 150:24:@47837.4]
  wire [31:0] x622_x13_1_io_b; // @[Math.scala 150:24:@47837.4]
  wire  x622_x13_1_io_flow; // @[Math.scala 150:24:@47837.4]
  wire [31:0] x622_x13_1_io_result; // @[Math.scala 150:24:@47837.4]
  wire  x623_x14_1_clock; // @[Math.scala 150:24:@47847.4]
  wire  x623_x14_1_reset; // @[Math.scala 150:24:@47847.4]
  wire [31:0] x623_x14_1_io_a; // @[Math.scala 150:24:@47847.4]
  wire [31:0] x623_x14_1_io_b; // @[Math.scala 150:24:@47847.4]
  wire  x623_x14_1_io_flow; // @[Math.scala 150:24:@47847.4]
  wire [31:0] x623_x14_1_io_result; // @[Math.scala 150:24:@47847.4]
  wire  x624_x13_1_clock; // @[Math.scala 150:24:@47857.4]
  wire  x624_x13_1_reset; // @[Math.scala 150:24:@47857.4]
  wire [31:0] x624_x13_1_io_a; // @[Math.scala 150:24:@47857.4]
  wire [31:0] x624_x13_1_io_b; // @[Math.scala 150:24:@47857.4]
  wire  x624_x13_1_io_flow; // @[Math.scala 150:24:@47857.4]
  wire [31:0] x624_x13_1_io_result; // @[Math.scala 150:24:@47857.4]
  wire  x625_x14_1_clock; // @[Math.scala 150:24:@47867.4]
  wire  x625_x14_1_reset; // @[Math.scala 150:24:@47867.4]
  wire [31:0] x625_x14_1_io_a; // @[Math.scala 150:24:@47867.4]
  wire [31:0] x625_x14_1_io_b; // @[Math.scala 150:24:@47867.4]
  wire  x625_x14_1_io_flow; // @[Math.scala 150:24:@47867.4]
  wire [31:0] x625_x14_1_io_result; // @[Math.scala 150:24:@47867.4]
  wire  x626_x13_1_clock; // @[Math.scala 150:24:@47877.4]
  wire  x626_x13_1_reset; // @[Math.scala 150:24:@47877.4]
  wire [31:0] x626_x13_1_io_a; // @[Math.scala 150:24:@47877.4]
  wire [31:0] x626_x13_1_io_b; // @[Math.scala 150:24:@47877.4]
  wire  x626_x13_1_io_flow; // @[Math.scala 150:24:@47877.4]
  wire [31:0] x626_x13_1_io_result; // @[Math.scala 150:24:@47877.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@47887.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@47887.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@47887.4]
  wire [31:0] RetimeWrapper_122_io_in; // @[package.scala 93:22:@47887.4]
  wire [31:0] RetimeWrapper_122_io_out; // @[package.scala 93:22:@47887.4]
  wire  x627_sum_1_clock; // @[Math.scala 150:24:@47896.4]
  wire  x627_sum_1_reset; // @[Math.scala 150:24:@47896.4]
  wire [31:0] x627_sum_1_io_a; // @[Math.scala 150:24:@47896.4]
  wire [31:0] x627_sum_1_io_b; // @[Math.scala 150:24:@47896.4]
  wire  x627_sum_1_io_flow; // @[Math.scala 150:24:@47896.4]
  wire [31:0] x627_sum_1_io_result; // @[Math.scala 150:24:@47896.4]
  wire [31:0] x628_1_io_b; // @[Math.scala 720:24:@47906.4]
  wire [31:0] x628_1_io_result; // @[Math.scala 720:24:@47906.4]
  wire  x629_mul_1_clock; // @[Math.scala 262:24:@47917.4]
  wire [31:0] x629_mul_1_io_a; // @[Math.scala 262:24:@47917.4]
  wire [31:0] x629_mul_1_io_b; // @[Math.scala 262:24:@47917.4]
  wire  x629_mul_1_io_flow; // @[Math.scala 262:24:@47917.4]
  wire [31:0] x629_mul_1_io_result; // @[Math.scala 262:24:@47917.4]
  wire [31:0] x630_1_io_b; // @[Math.scala 720:24:@47927.4]
  wire [31:0] x630_1_io_result; // @[Math.scala 720:24:@47927.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@47936.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@47936.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@47936.4]
  wire [31:0] RetimeWrapper_123_io_in; // @[package.scala 93:22:@47936.4]
  wire [31:0] RetimeWrapper_123_io_out; // @[package.scala 93:22:@47936.4]
  wire  x631_sub_1_clock; // @[Math.scala 191:24:@47945.4]
  wire  x631_sub_1_reset; // @[Math.scala 191:24:@47945.4]
  wire [31:0] x631_sub_1_io_a; // @[Math.scala 191:24:@47945.4]
  wire [31:0] x631_sub_1_io_b; // @[Math.scala 191:24:@47945.4]
  wire  x631_sub_1_io_flow; // @[Math.scala 191:24:@47945.4]
  wire [31:0] x631_sub_1_io_result; // @[Math.scala 191:24:@47945.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@47958.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@47958.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@47958.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@47958.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@47958.4]
  wire  x633_sub_1_clock; // @[Math.scala 191:24:@47967.4]
  wire  x633_sub_1_reset; // @[Math.scala 191:24:@47967.4]
  wire [31:0] x633_sub_1_io_a; // @[Math.scala 191:24:@47967.4]
  wire [31:0] x633_sub_1_io_b; // @[Math.scala 191:24:@47967.4]
  wire  x633_sub_1_io_flow; // @[Math.scala 191:24:@47967.4]
  wire [31:0] x633_sub_1_io_result; // @[Math.scala 191:24:@47967.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@47980.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@47980.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@47980.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@47980.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@47980.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@47992.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@47992.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@47992.4]
  wire [31:0] RetimeWrapper_126_io_in; // @[package.scala 93:22:@47992.4]
  wire [31:0] RetimeWrapper_126_io_out; // @[package.scala 93:22:@47992.4]
  wire [31:0] x637_1_io_b; // @[Math.scala 720:24:@48006.4]
  wire [31:0] x637_1_io_result; // @[Math.scala 720:24:@48006.4]
  wire  x638_mul_1_clock; // @[Math.scala 262:24:@48017.4]
  wire [31:0] x638_mul_1_io_a; // @[Math.scala 262:24:@48017.4]
  wire [31:0] x638_mul_1_io_b; // @[Math.scala 262:24:@48017.4]
  wire  x638_mul_1_io_flow; // @[Math.scala 262:24:@48017.4]
  wire [31:0] x638_mul_1_io_result; // @[Math.scala 262:24:@48017.4]
  wire [31:0] x639_1_io_b; // @[Math.scala 720:24:@48027.4]
  wire [31:0] x639_1_io_result; // @[Math.scala 720:24:@48027.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@48036.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@48036.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@48036.4]
  wire [31:0] RetimeWrapper_127_io_in; // @[package.scala 93:22:@48036.4]
  wire [31:0] RetimeWrapper_127_io_out; // @[package.scala 93:22:@48036.4]
  wire  x640_sum_1_clock; // @[Math.scala 150:24:@48045.4]
  wire  x640_sum_1_reset; // @[Math.scala 150:24:@48045.4]
  wire [31:0] x640_sum_1_io_a; // @[Math.scala 150:24:@48045.4]
  wire [31:0] x640_sum_1_io_b; // @[Math.scala 150:24:@48045.4]
  wire  x640_sum_1_io_flow; // @[Math.scala 150:24:@48045.4]
  wire [31:0] x640_sum_1_io_result; // @[Math.scala 150:24:@48045.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@48065.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@48065.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@48065.4]
  wire [127:0] RetimeWrapper_128_io_in; // @[package.scala 93:22:@48065.4]
  wire [127:0] RetimeWrapper_128_io_out; // @[package.scala 93:22:@48065.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@48074.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@48074.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@48074.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@48074.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@48074.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@48083.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@48083.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@48083.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@48083.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@48083.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@48092.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@48092.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@48092.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@48092.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@48092.4]
  wire  b394; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 62:18:@44824.4]
  wire  b395; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 63:18:@44825.4]
  wire  _T_205; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 67:30:@44827.4]
  wire  _T_206; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 67:37:@44828.4]
  wire  _T_210; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 69:76:@44833.4]
  wire  _T_211; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 69:62:@44834.4]
  wire  _T_213; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 69:101:@44835.4]
  wire [127:0] x729_x396_D1_0_number; // @[package.scala 96:25:@44844.4 package.scala 96:25:@44845.4]
  wire [31:0] b392_number; // @[Math.scala 723:22:@44809.4 Math.scala 724:14:@44810.4]
  wire [31:0] _T_247; // @[Math.scala 406:49:@45009.4]
  wire [31:0] _T_249; // @[Math.scala 406:56:@45011.4]
  wire [31:0] _T_250; // @[Math.scala 406:56:@45012.4]
  wire [31:0] x709_number; // @[implicits.scala 133:21:@45013.4]
  wire [31:0] _T_260; // @[Math.scala 406:49:@45022.4]
  wire [31:0] _T_262; // @[Math.scala 406:56:@45024.4]
  wire [31:0] _T_263; // @[Math.scala 406:56:@45025.4]
  wire  _T_274; // @[FixedPoint.scala 50:25:@45043.4]
  wire [1:0] _T_278; // @[Bitwise.scala 72:12:@45045.4]
  wire [29:0] _T_279; // @[FixedPoint.scala 18:52:@45046.4]
  wire  _T_285; // @[Math.scala 451:55:@45048.4]
  wire [1:0] _T_286; // @[FixedPoint.scala 18:52:@45049.4]
  wire  _T_292; // @[Math.scala 451:110:@45051.4]
  wire  _T_293; // @[Math.scala 451:94:@45052.4]
  wire [31:0] _T_295; // @[Cat.scala 30:58:@45054.4]
  wire [31:0] x404_1_number; // @[Math.scala 454:20:@45055.4]
  wire [39:0] _GEN_0; // @[Math.scala 461:32:@45060.4]
  wire [39:0] _T_300; // @[Math.scala 461:32:@45060.4]
  wire [37:0] _GEN_1; // @[Math.scala 461:32:@45065.4]
  wire [37:0] _T_303; // @[Math.scala 461:32:@45065.4]
  wire  _T_339; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:101:@45163.4]
  wire  _T_343; // @[package.scala 96:25:@45171.4 package.scala 96:25:@45172.4]
  wire  _T_345; // @[implicits.scala 55:10:@45173.4]
  wire  _T_346; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:118:@45174.4]
  wire  _T_348; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:207:@45176.4]
  wire  _T_349; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:226:@45177.4]
  wire  x734_b394_D24; // @[package.scala 96:25:@45142.4 package.scala 96:25:@45143.4]
  wire  _T_350; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:252:@45178.4]
  wire  x736_b395_D24; // @[package.scala 96:25:@45160.4 package.scala 96:25:@45161.4]
  wire  _T_394; // @[package.scala 96:25:@45278.4 package.scala 96:25:@45279.4]
  wire  _T_396; // @[implicits.scala 55:10:@45280.4]
  wire  _T_397; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:118:@45281.4]
  wire  _T_399; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:207:@45283.4]
  wire  _T_400; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:226:@45284.4]
  wire  _T_401; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:252:@45285.4]
  wire  _T_442; // @[package.scala 96:25:@45376.4 package.scala 96:25:@45377.4]
  wire  _T_444; // @[implicits.scala 55:10:@45378.4]
  wire  _T_445; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:118:@45379.4]
  wire  _T_447; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:207:@45381.4]
  wire  _T_448; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:226:@45382.4]
  wire  _T_449; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:252:@45383.4]
  wire  _T_490; // @[package.scala 96:25:@45474.4 package.scala 96:25:@45475.4]
  wire  _T_492; // @[implicits.scala 55:10:@45476.4]
  wire  _T_493; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:166:@45477.4]
  wire  _T_495; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:255:@45479.4]
  wire  _T_496; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:274:@45480.4]
  wire  _T_497; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:300:@45481.4]
  wire [31:0] x747_b392_D26_number; // @[package.scala 96:25:@45495.4 package.scala 96:25:@45496.4]
  wire [31:0] _T_509; // @[Math.scala 476:37:@45503.4]
  wire [31:0] x748_x421_rdcol_D26_number; // @[package.scala 96:25:@45520.4 package.scala 96:25:@45521.4]
  wire [31:0] _T_522; // @[Math.scala 476:37:@45526.4]
  wire  x749_x428_D1; // @[package.scala 96:25:@45543.4 package.scala 96:25:@45544.4]
  wire  x429; // @[package.scala 96:25:@45534.4 package.scala 96:25:@45535.4]
  wire  x430; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 203:24:@45547.4]
  wire  _T_563; // @[package.scala 96:25:@45615.4 package.scala 96:25:@45616.4]
  wire  _T_565; // @[implicits.scala 55:10:@45617.4]
  wire  _T_566; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 222:194:@45618.4]
  wire  x754_x431_D20; // @[package.scala 96:25:@45594.4 package.scala 96:25:@45595.4]
  wire  _T_567; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 222:283:@45619.4]
  wire  x753_b394_D48; // @[package.scala 96:25:@45585.4 package.scala 96:25:@45586.4]
  wire  _T_568; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 222:291:@45620.4]
  wire  x755_b395_D48; // @[package.scala 96:25:@45603.4 package.scala 96:25:@45604.4]
  wire [31:0] x756_x415_rdcol_D26_number; // @[package.scala 96:25:@45636.4 package.scala 96:25:@45637.4]
  wire [31:0] _T_579; // @[Math.scala 476:37:@45642.4]
  wire  x434; // @[package.scala 96:25:@45650.4 package.scala 96:25:@45651.4]
  wire  x435; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 230:24:@45654.4]
  wire  _T_608; // @[package.scala 96:25:@45695.4 package.scala 96:25:@45696.4]
  wire  _T_610; // @[implicits.scala 55:10:@45697.4]
  wire  _T_611; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:194:@45698.4]
  wire  x758_x436_D20; // @[package.scala 96:25:@45674.4 package.scala 96:25:@45675.4]
  wire  _T_612; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:283:@45699.4]
  wire  _T_613; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:291:@45700.4]
  wire [31:0] x760_x409_rdcol_D26_number; // @[package.scala 96:25:@45716.4 package.scala 96:25:@45717.4]
  wire [31:0] _T_624; // @[Math.scala 476:37:@45722.4]
  wire  x439; // @[package.scala 96:25:@45730.4 package.scala 96:25:@45731.4]
  wire  x440; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 251:24:@45734.4]
  wire  _T_653; // @[package.scala 96:25:@45775.4 package.scala 96:25:@45776.4]
  wire  _T_655; // @[implicits.scala 55:10:@45777.4]
  wire  _T_656; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:194:@45778.4]
  wire  x763_x441_D20; // @[package.scala 96:25:@45763.4 package.scala 96:25:@45764.4]
  wire  _T_657; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:283:@45779.4]
  wire  _T_658; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:291:@45780.4]
  wire [31:0] x764_b393_D26_number; // @[package.scala 96:25:@45796.4 package.scala 96:25:@45797.4]
  wire [31:0] _T_669; // @[Math.scala 476:37:@45802.4]
  wire  x428; // @[package.scala 96:25:@45511.4 package.scala 96:25:@45512.4]
  wire  x444; // @[package.scala 96:25:@45810.4 package.scala 96:25:@45811.4]
  wire  x445; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 272:24:@45814.4]
  wire  _T_698; // @[package.scala 96:25:@45855.4 package.scala 96:25:@45856.4]
  wire  _T_700; // @[implicits.scala 55:10:@45857.4]
  wire  _T_701; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:194:@45858.4]
  wire  x767_x446_D21; // @[package.scala 96:25:@45843.4 package.scala 96:25:@45844.4]
  wire  _T_702; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:283:@45859.4]
  wire  _T_703; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:291:@45860.4]
  wire [31:0] x449_rdcol_number; // @[Math.scala 154:22:@45879.4 Math.scala 155:14:@45880.4]
  wire [31:0] _T_718; // @[Math.scala 476:37:@45885.4]
  wire  x450; // @[package.scala 96:25:@45893.4 package.scala 96:25:@45894.4]
  wire  x451; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 293:24:@45897.4]
  wire  _T_766; // @[package.scala 96:25:@45974.4 package.scala 96:25:@45975.4]
  wire  _T_768; // @[implicits.scala 55:10:@45976.4]
  wire  _T_769; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:194:@45977.4]
  wire  x770_x452_D20; // @[package.scala 96:25:@45962.4 package.scala 96:25:@45963.4]
  wire  _T_770; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:283:@45978.4]
  wire  _T_771; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:291:@45979.4]
  wire [31:0] x458_rdcol_number; // @[Math.scala 154:22:@45998.4 Math.scala 155:14:@45999.4]
  wire [31:0] _T_786; // @[Math.scala 476:37:@46004.4]
  wire  x459; // @[package.scala 96:25:@46012.4 package.scala 96:25:@46013.4]
  wire  x460; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 328:59:@46016.4]
  wire  _T_829; // @[package.scala 96:25:@46082.4 package.scala 96:25:@46083.4]
  wire  _T_831; // @[implicits.scala 55:10:@46084.4]
  wire  _T_832; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 345:194:@46085.4]
  wire  x771_x461_D20; // @[package.scala 96:25:@46061.4 package.scala 96:25:@46062.4]
  wire  _T_833; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 345:283:@46086.4]
  wire  _T_834; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 345:291:@46087.4]
  wire [31:0] x467_rdrow_number; // @[Math.scala 195:22:@46106.4 Math.scala 196:14:@46107.4]
  wire [31:0] _T_851; // @[Math.scala 406:49:@46113.4]
  wire [31:0] _T_853; // @[Math.scala 406:56:@46115.4]
  wire [31:0] _T_854; // @[Math.scala 406:56:@46116.4]
  wire [31:0] x714_number; // @[implicits.scala 133:21:@46117.4]
  wire  x469; // @[package.scala 96:25:@46131.4 package.scala 96:25:@46132.4]
  wire  x470; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 355:24:@46135.4]
  wire [31:0] _T_877; // @[Math.scala 406:49:@46144.4]
  wire [31:0] _T_879; // @[Math.scala 406:56:@46146.4]
  wire [31:0] _T_880; // @[Math.scala 406:56:@46147.4]
  wire [31:0] _T_884; // @[package.scala 96:25:@46155.4]
  wire  _T_888; // @[FixedPoint.scala 50:25:@46162.4]
  wire [1:0] _T_892; // @[Bitwise.scala 72:12:@46164.4]
  wire [29:0] _T_893; // @[FixedPoint.scala 18:52:@46165.4]
  wire  _T_899; // @[Math.scala 451:55:@46167.4]
  wire [1:0] _T_900; // @[FixedPoint.scala 18:52:@46168.4]
  wire  _T_906; // @[Math.scala 451:110:@46170.4]
  wire  _T_907; // @[Math.scala 451:94:@46171.4]
  wire [31:0] _T_911; // @[package.scala 96:25:@46179.4 package.scala 96:25:@46180.4]
  wire [31:0] x473_1_number; // @[Math.scala 454:20:@46181.4]
  wire [39:0] _GEN_2; // @[Math.scala 461:32:@46186.4]
  wire [39:0] _T_916; // @[Math.scala 461:32:@46186.4]
  wire [37:0] _GEN_3; // @[Math.scala 461:32:@46191.4]
  wire [37:0] _T_919; // @[Math.scala 461:32:@46191.4]
  wire  _T_949; // @[package.scala 96:25:@46259.4 package.scala 96:25:@46260.4]
  wire  _T_951; // @[implicits.scala 55:10:@46261.4]
  wire  _T_952; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:194:@46262.4]
  wire  x776_x471_D20; // @[package.scala 96:25:@46247.4 package.scala 96:25:@46248.4]
  wire  _T_953; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:283:@46263.4]
  wire  _T_954; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:291:@46264.4]
  wire  x478; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 386:24:@46275.4]
  wire  _T_981; // @[package.scala 96:25:@46317.4 package.scala 96:25:@46318.4]
  wire  _T_983; // @[implicits.scala 55:10:@46319.4]
  wire  _T_984; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:194:@46320.4]
  wire  x778_x479_D20; // @[package.scala 96:25:@46305.4 package.scala 96:25:@46306.4]
  wire  _T_985; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:283:@46321.4]
  wire  _T_986; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:291:@46322.4]
  wire  x483; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 403:24:@46333.4]
  wire  _T_1013; // @[package.scala 96:25:@46375.4 package.scala 96:25:@46376.4]
  wire  _T_1015; // @[implicits.scala 55:10:@46377.4]
  wire  _T_1016; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:194:@46378.4]
  wire  x780_x484_D20; // @[package.scala 96:25:@46363.4 package.scala 96:25:@46364.4]
  wire  _T_1017; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:283:@46379.4]
  wire  _T_1018; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:291:@46380.4]
  wire  x781_x444_D1; // @[package.scala 96:25:@46396.4 package.scala 96:25:@46397.4]
  wire  x488; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 428:59:@46400.4]
  wire  _T_1056; // @[package.scala 96:25:@46462.4 package.scala 96:25:@46463.4]
  wire  _T_1058; // @[implicits.scala 55:10:@46464.4]
  wire  _T_1059; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:194:@46465.4]
  wire  x784_x489_D20; // @[package.scala 96:25:@46441.4 package.scala 96:25:@46442.4]
  wire  _T_1060; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:283:@46466.4]
  wire  _T_1061; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:291:@46467.4]
  wire  x493; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 451:59:@46478.4]
  wire  _T_1085; // @[package.scala 96:25:@46511.4 package.scala 96:25:@46512.4]
  wire  _T_1087; // @[implicits.scala 55:10:@46513.4]
  wire  _T_1088; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:194:@46514.4]
  wire  x786_x494_D20; // @[package.scala 96:25:@46499.4 package.scala 96:25:@46500.4]
  wire  _T_1089; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:283:@46515.4]
  wire  _T_1090; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:291:@46516.4]
  wire  x498; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 466:59:@46527.4]
  wire  _T_1114; // @[package.scala 96:25:@46560.4 package.scala 96:25:@46561.4]
  wire  _T_1116; // @[implicits.scala 55:10:@46562.4]
  wire  _T_1117; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:194:@46563.4]
  wire  x787_x499_D20; // @[package.scala 96:25:@46548.4 package.scala 96:25:@46549.4]
  wire  _T_1118; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:283:@46564.4]
  wire  _T_1119; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:291:@46565.4]
  wire [31:0] x503_rdrow_number; // @[Math.scala 195:22:@46584.4 Math.scala 196:14:@46585.4]
  wire [31:0] _T_1136; // @[Math.scala 406:49:@46591.4]
  wire [31:0] _T_1138; // @[Math.scala 406:56:@46593.4]
  wire [31:0] _T_1139; // @[Math.scala 406:56:@46594.4]
  wire [31:0] x719_number; // @[implicits.scala 133:21:@46595.4]
  wire  x505; // @[package.scala 96:25:@46609.4 package.scala 96:25:@46610.4]
  wire  x506; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 487:24:@46613.4]
  wire [31:0] _T_1162; // @[Math.scala 406:49:@46622.4]
  wire [31:0] _T_1164; // @[Math.scala 406:56:@46624.4]
  wire [31:0] _T_1165; // @[Math.scala 406:56:@46625.4]
  wire [31:0] _T_1169; // @[package.scala 96:25:@46633.4]
  wire  _T_1173; // @[FixedPoint.scala 50:25:@46640.4]
  wire [1:0] _T_1177; // @[Bitwise.scala 72:12:@46642.4]
  wire [29:0] _T_1178; // @[FixedPoint.scala 18:52:@46643.4]
  wire  _T_1184; // @[Math.scala 451:55:@46645.4]
  wire [1:0] _T_1185; // @[FixedPoint.scala 18:52:@46646.4]
  wire  _T_1191; // @[Math.scala 451:110:@46648.4]
  wire  _T_1192; // @[Math.scala 451:94:@46649.4]
  wire [31:0] _T_1196; // @[package.scala 96:25:@46657.4 package.scala 96:25:@46658.4]
  wire [31:0] x509_1_number; // @[Math.scala 454:20:@46659.4]
  wire [39:0] _GEN_4; // @[Math.scala 461:32:@46664.4]
  wire [39:0] _T_1201; // @[Math.scala 461:32:@46664.4]
  wire [37:0] _GEN_5; // @[Math.scala 461:32:@46669.4]
  wire [37:0] _T_1204; // @[Math.scala 461:32:@46669.4]
  wire  _T_1231; // @[package.scala 96:25:@46728.4 package.scala 96:25:@46729.4]
  wire  _T_1233; // @[implicits.scala 55:10:@46730.4]
  wire  _T_1234; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 512:194:@46731.4]
  wire  x789_x507_D20; // @[package.scala 96:25:@46707.4 package.scala 96:25:@46708.4]
  wire  _T_1235; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 512:283:@46732.4]
  wire  _T_1236; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 512:291:@46733.4]
  wire  x514; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 516:24:@46744.4]
  wire  _T_1260; // @[package.scala 96:25:@46777.4 package.scala 96:25:@46778.4]
  wire  _T_1262; // @[implicits.scala 55:10:@46779.4]
  wire  _T_1263; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:194:@46780.4]
  wire  x791_x515_D20; // @[package.scala 96:25:@46765.4 package.scala 96:25:@46766.4]
  wire  _T_1264; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:283:@46781.4]
  wire  _T_1265; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:291:@46782.4]
  wire  x519; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 531:24:@46793.4]
  wire  _T_1289; // @[package.scala 96:25:@46826.4 package.scala 96:25:@46827.4]
  wire  _T_1291; // @[implicits.scala 55:10:@46828.4]
  wire  _T_1292; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:194:@46829.4]
  wire  x792_x520_D20; // @[package.scala 96:25:@46814.4 package.scala 96:25:@46815.4]
  wire  _T_1293; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:283:@46830.4]
  wire  _T_1294; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:326:@46831.4]
  wire  x524; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 552:59:@46842.4]
  wire  _T_1326; // @[package.scala 96:25:@46895.4 package.scala 96:25:@46896.4]
  wire  _T_1328; // @[implicits.scala 55:10:@46897.4]
  wire  _T_1329; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:194:@46898.4]
  wire  x795_x525_D20; // @[package.scala 96:25:@46883.4 package.scala 96:25:@46884.4]
  wire  _T_1330; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:283:@46899.4]
  wire  _T_1331; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:291:@46900.4]
  wire  x529; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 573:59:@46911.4]
  wire  _T_1355; // @[package.scala 96:25:@46944.4 package.scala 96:25:@46945.4]
  wire  _T_1357; // @[implicits.scala 55:10:@46946.4]
  wire  _T_1358; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:194:@46947.4]
  wire  x796_x530_D20; // @[package.scala 96:25:@46932.4 package.scala 96:25:@46933.4]
  wire  _T_1359; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:283:@46948.4]
  wire  _T_1360; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:291:@46949.4]
  wire  x534; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 588:59:@46960.4]
  wire  _T_1384; // @[package.scala 96:25:@46993.4 package.scala 96:25:@46994.4]
  wire  _T_1386; // @[implicits.scala 55:10:@46995.4]
  wire  _T_1387; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 599:194:@46996.4]
  wire  x797_x535_D20; // @[package.scala 96:25:@46981.4 package.scala 96:25:@46982.4]
  wire  _T_1388; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 599:283:@46997.4]
  wire  _T_1389; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 599:291:@46998.4]
  wire [31:0] x437_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 239:29:@45686.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:338:@45707.4]
  wire [32:0] _GEN_6; // @[Math.scala 461:32:@47010.4]
  wire [32:0] _T_1394; // @[Math.scala 461:32:@47010.4]
  wire [31:0] x476_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 378:29:@46250.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:408:@46271.4]
  wire [32:0] _GEN_7; // @[Math.scala 461:32:@47015.4]
  wire [32:0] _T_1397; // @[Math.scala 461:32:@47015.4]
  wire [31:0] x481_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 395:29:@46308.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:408:@46329.4]
  wire [33:0] _GEN_8; // @[Math.scala 461:32:@47020.4]
  wire [33:0] _T_1400; // @[Math.scala 461:32:@47020.4]
  wire [31:0] x486_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 412:29:@46366.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:408:@46387.4]
  wire [32:0] _GEN_9; // @[Math.scala 461:32:@47025.4]
  wire [32:0] _T_1403; // @[Math.scala 461:32:@47025.4]
  wire [31:0] x517_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 523:29:@46768.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:408:@46789.4]
  wire [32:0] _GEN_10; // @[Math.scala 461:32:@47030.4]
  wire [32:0] _T_1406; // @[Math.scala 461:32:@47030.4]
  wire [31:0] x555_sub_number; // @[Math.scala 195:22:@47168.4 Math.scala 196:14:@47169.4]
  wire [31:0] x557_sub_number; // @[Math.scala 195:22:@47190.4 Math.scala 196:14:@47191.4]
  wire  x556; // @[package.scala 96:25:@47180.4 package.scala 96:25:@47181.4]
  wire  x558; // @[package.scala 96:25:@47202.4 package.scala 96:25:@47203.4]
  wire  x559; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 647:24:@47206.4]
  wire [31:0] x800_x555_sub_D1_number; // @[package.scala 96:25:@47214.4 package.scala 96:25:@47215.4]
  wire [31:0] x442_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 260:29:@45766.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:338:@45787.4]
  wire [32:0] _GEN_11; // @[Math.scala 461:32:@47275.4]
  wire [32:0] _T_1506; // @[Math.scala 461:32:@47275.4]
  wire [32:0] _GEN_12; // @[Math.scala 461:32:@47280.4]
  wire [32:0] _T_1509; // @[Math.scala 461:32:@47280.4]
  wire [33:0] _GEN_13; // @[Math.scala 461:32:@47285.4]
  wire [33:0] _T_1512; // @[Math.scala 461:32:@47285.4]
  wire [31:0] x491_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 443:29:@46453.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:408:@46474.4]
  wire [32:0] _GEN_14; // @[Math.scala 461:32:@47290.4]
  wire [32:0] _T_1515; // @[Math.scala 461:32:@47290.4]
  wire [31:0] x522_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 544:29:@46817.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:443:@46838.4]
  wire [32:0] _GEN_15; // @[Math.scala 461:32:@47295.4]
  wire [32:0] _T_1518; // @[Math.scala 461:32:@47295.4]
  wire [31:0] x581_sub_number; // @[Math.scala 195:22:@47433.4 Math.scala 196:14:@47434.4]
  wire [31:0] x583_sub_number; // @[Math.scala 195:22:@47455.4 Math.scala 196:14:@47456.4]
  wire  x582; // @[package.scala 96:25:@47445.4 package.scala 96:25:@47446.4]
  wire  x584; // @[package.scala 96:25:@47467.4 package.scala 96:25:@47468.4]
  wire  x585; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 715:24:@47471.4]
  wire [31:0] x804_x581_sub_D1_number; // @[package.scala 96:25:@47479.4 package.scala 96:25:@47480.4]
  wire [31:0] x447_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 281:29:@45846.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:338:@45867.4]
  wire [32:0] _GEN_16; // @[Math.scala 461:32:@47538.4]
  wire [32:0] _T_1616; // @[Math.scala 461:32:@47538.4]
  wire [33:0] _GEN_17; // @[Math.scala 461:32:@47543.4]
  wire [33:0] _T_1619; // @[Math.scala 461:32:@47543.4]
  wire [31:0] x496_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 458:29:@46502.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:408:@46523.4]
  wire [32:0] _GEN_18; // @[Math.scala 461:32:@47548.4]
  wire [32:0] _T_1622; // @[Math.scala 461:32:@47548.4]
  wire [31:0] x527_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 565:29:@46886.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:408:@46907.4]
  wire [32:0] _GEN_19; // @[Math.scala 461:32:@47553.4]
  wire [32:0] _T_1625; // @[Math.scala 461:32:@47553.4]
  wire [31:0] x606_sub_number; // @[Math.scala 195:22:@47693.4 Math.scala 196:14:@47694.4]
  wire [31:0] x608_sub_number; // @[Math.scala 195:22:@47715.4 Math.scala 196:14:@47716.4]
  wire  x607; // @[package.scala 96:25:@47705.4 package.scala 96:25:@47706.4]
  wire  x609; // @[package.scala 96:25:@47727.4 package.scala 96:25:@47728.4]
  wire  x610; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 781:24:@47731.4]
  wire [31:0] x808_x606_sub_D1_number; // @[package.scala 96:25:@47739.4 package.scala 96:25:@47740.4]
  wire [31:0] x456_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 316:29:@45965.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:408:@45986.4]
  wire [32:0] _GEN_20; // @[Math.scala 461:32:@47798.4]
  wire [32:0] _T_1725; // @[Math.scala 461:32:@47798.4]
  wire [33:0] _GEN_21; // @[Math.scala 461:32:@47803.4]
  wire [33:0] _T_1728; // @[Math.scala 461:32:@47803.4]
  wire [31:0] x501_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 473:29:@46551.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:408:@46572.4]
  wire [32:0] _GEN_22; // @[Math.scala 461:32:@47808.4]
  wire [32:0] _T_1731; // @[Math.scala 461:32:@47808.4]
  wire [31:0] x532_rd_0_number; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 580:29:@46935.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:408:@46956.4]
  wire [32:0] _GEN_23; // @[Math.scala 461:32:@47813.4]
  wire [32:0] _T_1734; // @[Math.scala 461:32:@47813.4]
  wire [31:0] x631_sub_number; // @[Math.scala 195:22:@47951.4 Math.scala 196:14:@47952.4]
  wire [31:0] x633_sub_number; // @[Math.scala 195:22:@47973.4 Math.scala 196:14:@47974.4]
  wire  x632; // @[package.scala 96:25:@47963.4 package.scala 96:25:@47964.4]
  wire  x634; // @[package.scala 96:25:@47985.4 package.scala 96:25:@47986.4]
  wire  x635; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 839:24:@47989.4]
  wire [31:0] x812_x631_sub_D1_number; // @[package.scala 96:25:@47997.4 package.scala 96:25:@47998.4]
  wire [31:0] x615_sum_number; // @[Math.scala 154:22:@47793.4 Math.scala 155:14:@47794.4]
  wire [31:0] x640_sum_number; // @[Math.scala 154:22:@48051.4 Math.scala 155:14:@48052.4]
  wire [63:0] _T_1841; // @[Cat.scala 30:58:@48060.4]
  wire [31:0] x564_sum_number; // @[Math.scala 154:22:@47270.4 Math.scala 155:14:@47271.4]
  wire [31:0] x590_sum_number; // @[Math.scala 154:22:@47533.4 Math.scala 155:14:@47534.4]
  wire [63:0] _T_1842; // @[Cat.scala 30:58:@48061.4]
  wire  _T_1855; // @[package.scala 96:25:@48097.4 package.scala 96:25:@48098.4]
  wire  _T_1857; // @[implicits.scala 55:10:@48099.4]
  wire  x815_b394_D72; // @[package.scala 96:25:@48088.4 package.scala 96:25:@48089.4]
  wire  _T_1858; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 863:117:@48100.4]
  wire  x814_b395_D72; // @[package.scala 96:25:@48079.4 package.scala 96:25:@48080.4]
  wire  _T_1859; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 863:123:@48101.4]
  wire [31:0] x731_x407_sum_D3_number; // @[package.scala 96:25:@45115.4 package.scala 96:25:@45116.4]
  wire [31:0] x732_x710_D24_number; // @[package.scala 96:25:@45124.4 package.scala 96:25:@45125.4]
  wire [31:0] x733_x403_D8_number; // @[package.scala 96:25:@45133.4 package.scala 96:25:@45134.4]
  wire [31:0] x738_x411_D7_number; // @[package.scala 96:25:@45249.4 package.scala 96:25:@45250.4]
  wire [31:0] x739_x413_sum_D2_number; // @[package.scala 96:25:@45258.4 package.scala 96:25:@45259.4]
  wire [31:0] x741_x417_D7_number; // @[package.scala 96:25:@45347.4 package.scala 96:25:@45348.4]
  wire [31:0] x743_x419_sum_D2_number; // @[package.scala 96:25:@45365.4 package.scala 96:25:@45366.4]
  wire [31:0] x744_x425_sum_D2_number; // @[package.scala 96:25:@45445.4 package.scala 96:25:@45446.4]
  wire [31:0] x745_x423_D7_number; // @[package.scala 96:25:@45454.4 package.scala 96:25:@45455.4]
  wire [31:0] x750_x710_D48_number; // @[package.scala 96:25:@45558.4 package.scala 96:25:@45559.4]
  wire [31:0] x751_x425_sum_D26_number; // @[package.scala 96:25:@45567.4 package.scala 96:25:@45568.4]
  wire [31:0] x752_x423_D31_number; // @[package.scala 96:25:@45576.4 package.scala 96:25:@45577.4]
  wire [31:0] x757_x417_D31_number; // @[package.scala 96:25:@45665.4 package.scala 96:25:@45666.4]
  wire [31:0] x759_x419_sum_D26_number; // @[package.scala 96:25:@45683.4 package.scala 96:25:@45684.4]
  wire [31:0] x761_x411_D31_number; // @[package.scala 96:25:@45745.4 package.scala 96:25:@45746.4]
  wire [31:0] x762_x413_sum_D26_number; // @[package.scala 96:25:@45754.4 package.scala 96:25:@45755.4]
  wire [31:0] x765_x407_sum_D27_number; // @[package.scala 96:25:@45825.4 package.scala 96:25:@45826.4]
  wire [31:0] x766_x403_D32_number; // @[package.scala 96:25:@45834.4 package.scala 96:25:@45835.4]
  wire [31:0] x455_sum_number; // @[Math.scala 154:22:@45944.4 Math.scala 155:14:@45945.4]
  wire [31:0] x769_x453_D5_number; // @[package.scala 96:25:@45953.4 package.scala 96:25:@45954.4]
  wire [31:0] x464_sum_number; // @[Math.scala 154:22:@46052.4 Math.scala 155:14:@46053.4]
  wire [31:0] x772_x462_D5_number; // @[package.scala 96:25:@46070.4 package.scala 96:25:@46071.4]
  wire [31:0] x475_sum_number; // @[Math.scala 154:22:@46229.4 Math.scala 155:14:@46230.4]
  wire [31:0] x775_x715_D20_number; // @[package.scala 96:25:@46238.4 package.scala 96:25:@46239.4]
  wire [31:0] x480_sum_number; // @[Math.scala 154:22:@46296.4 Math.scala 155:14:@46297.4]
  wire [31:0] x485_sum_number; // @[Math.scala 154:22:@46354.4 Math.scala 155:14:@46355.4]
  wire [31:0] x785_x490_sum_D1_number; // @[package.scala 96:25:@46450.4 package.scala 96:25:@46451.4]
  wire [31:0] x495_sum_number; // @[Math.scala 154:22:@46490.4 Math.scala 155:14:@46491.4]
  wire [31:0] x500_sum_number; // @[Math.scala 154:22:@46539.4 Math.scala 155:14:@46540.4]
  wire [31:0] x511_sum_number; // @[Math.scala 154:22:@46698.4 Math.scala 155:14:@46699.4]
  wire [31:0] x790_x720_D20_number; // @[package.scala 96:25:@46716.4 package.scala 96:25:@46717.4]
  wire [31:0] x516_sum_number; // @[Math.scala 154:22:@46756.4 Math.scala 155:14:@46757.4]
  wire [31:0] x521_sum_number; // @[Math.scala 154:22:@46805.4 Math.scala 155:14:@46806.4]
  wire [31:0] x794_x526_sum_D1_number; // @[package.scala 96:25:@46874.4 package.scala 96:25:@46875.4]
  wire [31:0] x531_sum_number; // @[Math.scala 154:22:@46923.4 Math.scala 155:14:@46924.4]
  wire [31:0] x536_sum_number; // @[Math.scala 154:22:@46972.4 Math.scala 155:14:@46973.4]
  _ _ ( // @[Math.scala 720:24:@44804.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@44816.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_56 RetimeWrapper ( // @[package.scala 93:22:@44839.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x398_lb_0 x398_lb_0 ( // @[m_x398_lb_0.scala 47:17:@44849.4]
    .clock(x398_lb_0_clock),
    .reset(x398_lb_0_reset),
    .io_rPort_17_banks_1(x398_lb_0_io_rPort_17_banks_1),
    .io_rPort_17_banks_0(x398_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x398_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x398_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x398_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x398_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_1(x398_lb_0_io_rPort_16_banks_1),
    .io_rPort_16_banks_0(x398_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x398_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x398_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x398_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x398_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_1(x398_lb_0_io_rPort_15_banks_1),
    .io_rPort_15_banks_0(x398_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x398_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x398_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x398_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x398_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_1(x398_lb_0_io_rPort_14_banks_1),
    .io_rPort_14_banks_0(x398_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x398_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x398_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x398_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x398_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_1(x398_lb_0_io_rPort_13_banks_1),
    .io_rPort_13_banks_0(x398_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x398_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x398_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x398_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x398_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_1(x398_lb_0_io_rPort_12_banks_1),
    .io_rPort_12_banks_0(x398_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x398_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x398_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x398_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x398_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_1(x398_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x398_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x398_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x398_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x398_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x398_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x398_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x398_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x398_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x398_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x398_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x398_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x398_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x398_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x398_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x398_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x398_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x398_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x398_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x398_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x398_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x398_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x398_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x398_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x398_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x398_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x398_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x398_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x398_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x398_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x398_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x398_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x398_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x398_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x398_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x398_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x398_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x398_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x398_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x398_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x398_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x398_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x398_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x398_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x398_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x398_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x398_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x398_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x398_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x398_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x398_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x398_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x398_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x398_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x398_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x398_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x398_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x398_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x398_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x398_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x398_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x398_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x398_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x398_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x398_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x398_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x398_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x398_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x398_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x398_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x398_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x398_lb_0_io_rPort_0_output_0),
    .io_wPort_3_banks_1(x398_lb_0_io_wPort_3_banks_1),
    .io_wPort_3_banks_0(x398_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x398_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x398_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x398_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_1(x398_lb_0_io_wPort_2_banks_1),
    .io_wPort_2_banks_0(x398_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x398_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x398_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x398_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_1(x398_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x398_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x398_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x398_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x398_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x398_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x398_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x398_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x398_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x398_lb_0_io_wPort_0_en_0)
  );
  x403 x403_1 ( // @[Math.scala 366:24:@45032.4]
    .clock(x403_1_clock),
    .io_a(x403_1_io_a),
    .io_flow(x403_1_io_flow),
    .io_result(x403_1_io_result)
  );
  x367_sum x713_sum_1 ( // @[Math.scala 150:24:@45069.4]
    .clock(x713_sum_1_clock),
    .reset(x713_sum_1_reset),
    .io_a(x713_sum_1_io_a),
    .io_b(x713_sum_1_io_b),
    .io_flow(x713_sum_1_io_flow),
    .io_result(x713_sum_1_io_result)
  );
  x406_div x406_div_1 ( // @[Math.scala 327:24:@45081.4]
    .clock(x406_div_1_clock),
    .io_a(x406_div_1_io_a),
    .io_flow(x406_div_1_io_flow),
    .io_result(x406_div_1_io_result)
  );
  RetimeWrapper_298 RetimeWrapper_1 ( // @[package.scala 93:22:@45091.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x367_sum x407_sum_1 ( // @[Math.scala 150:24:@45100.4]
    .clock(x407_sum_1_clock),
    .reset(x407_sum_1_reset),
    .io_a(x407_sum_1_io_a),
    .io_b(x407_sum_1_io_b),
    .io_flow(x407_sum_1_io_flow),
    .io_result(x407_sum_1_io_result)
  );
  RetimeWrapper_300 RetimeWrapper_2 ( // @[package.scala 93:22:@45110.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_301 RetimeWrapper_3 ( // @[package.scala 93:22:@45119.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_302 RetimeWrapper_4 ( // @[package.scala 93:22:@45128.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_5 ( // @[package.scala 93:22:@45137.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_304 RetimeWrapper_6 ( // @[package.scala 93:22:@45146.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_7 ( // @[package.scala 93:22:@45155.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_8 ( // @[package.scala 93:22:@45166.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x367_sum x409_rdcol_1 ( // @[Math.scala 150:24:@45189.4]
    .clock(x409_rdcol_1_clock),
    .reset(x409_rdcol_1_reset),
    .io_a(x409_rdcol_1_io_a),
    .io_b(x409_rdcol_1_io_b),
    .io_flow(x409_rdcol_1_io_flow),
    .io_result(x409_rdcol_1_io_result)
  );
  x403 x411_1 ( // @[Math.scala 366:24:@45203.4]
    .clock(x411_1_clock),
    .io_a(x411_1_io_a),
    .io_flow(x411_1_io_flow),
    .io_result(x411_1_io_result)
  );
  x406_div x412_div_1 ( // @[Math.scala 327:24:@45215.4]
    .clock(x412_div_1_clock),
    .io_a(x412_div_1_io_a),
    .io_flow(x412_div_1_io_flow),
    .io_result(x412_div_1_io_result)
  );
  RetimeWrapper_308 RetimeWrapper_9 ( // @[package.scala 93:22:@45225.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  x367_sum x413_sum_1 ( // @[Math.scala 150:24:@45234.4]
    .clock(x413_sum_1_clock),
    .reset(x413_sum_1_reset),
    .io_a(x413_sum_1_io_a),
    .io_b(x413_sum_1_io_b),
    .io_flow(x413_sum_1_io_flow),
    .io_result(x413_sum_1_io_result)
  );
  RetimeWrapper_310 RetimeWrapper_10 ( // @[package.scala 93:22:@45244.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_11 ( // @[package.scala 93:22:@45253.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_304 RetimeWrapper_12 ( // @[package.scala 93:22:@45262.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_13 ( // @[package.scala 93:22:@45273.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x367_sum x415_rdcol_1 ( // @[Math.scala 150:24:@45296.4]
    .clock(x415_rdcol_1_clock),
    .reset(x415_rdcol_1_reset),
    .io_a(x415_rdcol_1_io_a),
    .io_b(x415_rdcol_1_io_b),
    .io_flow(x415_rdcol_1_io_flow),
    .io_result(x415_rdcol_1_io_result)
  );
  x403 x417_1 ( // @[Math.scala 366:24:@45310.4]
    .clock(x417_1_clock),
    .io_a(x417_1_io_a),
    .io_flow(x417_1_io_flow),
    .io_result(x417_1_io_result)
  );
  x406_div x418_div_1 ( // @[Math.scala 327:24:@45322.4]
    .clock(x418_div_1_clock),
    .io_a(x418_div_1_io_a),
    .io_flow(x418_div_1_io_flow),
    .io_result(x418_div_1_io_result)
  );
  x367_sum x419_sum_1 ( // @[Math.scala 150:24:@45332.4]
    .clock(x419_sum_1_clock),
    .reset(x419_sum_1_reset),
    .io_a(x419_sum_1_io_a),
    .io_b(x419_sum_1_io_b),
    .io_flow(x419_sum_1_io_flow),
    .io_result(x419_sum_1_io_result)
  );
  RetimeWrapper_310 RetimeWrapper_14 ( // @[package.scala 93:22:@45342.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_304 RetimeWrapper_15 ( // @[package.scala 93:22:@45351.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_16 ( // @[package.scala 93:22:@45360.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_17 ( // @[package.scala 93:22:@45371.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x367_sum x421_rdcol_1 ( // @[Math.scala 150:24:@45394.4]
    .clock(x421_rdcol_1_clock),
    .reset(x421_rdcol_1_reset),
    .io_a(x421_rdcol_1_io_a),
    .io_b(x421_rdcol_1_io_b),
    .io_flow(x421_rdcol_1_io_flow),
    .io_result(x421_rdcol_1_io_result)
  );
  x403 x423_1 ( // @[Math.scala 366:24:@45408.4]
    .clock(x423_1_clock),
    .io_a(x423_1_io_a),
    .io_flow(x423_1_io_flow),
    .io_result(x423_1_io_result)
  );
  x406_div x424_div_1 ( // @[Math.scala 327:24:@45420.4]
    .clock(x424_div_1_clock),
    .io_a(x424_div_1_io_a),
    .io_flow(x424_div_1_io_flow),
    .io_result(x424_div_1_io_result)
  );
  x367_sum x425_sum_1 ( // @[Math.scala 150:24:@45430.4]
    .clock(x425_sum_1_clock),
    .reset(x425_sum_1_reset),
    .io_a(x425_sum_1_io_a),
    .io_b(x425_sum_1_io_b),
    .io_flow(x425_sum_1_io_flow),
    .io_result(x425_sum_1_io_result)
  );
  RetimeWrapper_311 RetimeWrapper_18 ( // @[package.scala 93:22:@45440.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_310 RetimeWrapper_19 ( // @[package.scala 93:22:@45449.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_304 RetimeWrapper_20 ( // @[package.scala 93:22:@45458.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_21 ( // @[package.scala 93:22:@45469.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_22 ( // @[package.scala 93:22:@45490.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@45506.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_24 ( // @[package.scala 93:22:@45515.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@45529.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@45538.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_331 RetimeWrapper_27 ( // @[package.scala 93:22:@45553.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_28 ( // @[package.scala 93:22:@45562.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_29 ( // @[package.scala 93:22:@45571.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_30 ( // @[package.scala 93:22:@45580.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_31 ( // @[package.scala 93:22:@45589.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_32 ( // @[package.scala 93:22:@45598.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_33 ( // @[package.scala 93:22:@45610.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_34 ( // @[package.scala 93:22:@45631.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@45645.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_36 ( // @[package.scala 93:22:@45660.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_37 ( // @[package.scala 93:22:@45669.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_38 ( // @[package.scala 93:22:@45678.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_39 ( // @[package.scala 93:22:@45690.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_40 ( // @[package.scala 93:22:@45711.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@45725.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_42 ( // @[package.scala 93:22:@45740.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_43 ( // @[package.scala 93:22:@45749.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_44 ( // @[package.scala 93:22:@45758.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_45 ( // @[package.scala 93:22:@45770.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_46 ( // @[package.scala 93:22:@45791.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper RetimeWrapper_47 ( // @[package.scala 93:22:@45805.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_48 ( // @[package.scala 93:22:@45820.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_353 RetimeWrapper_49 ( // @[package.scala 93:22:@45829.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_354 RetimeWrapper_50 ( // @[package.scala 93:22:@45838.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_51 ( // @[package.scala 93:22:@45850.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x367_sum x449_rdcol_1 ( // @[Math.scala 150:24:@45873.4]
    .clock(x449_rdcol_1_clock),
    .reset(x449_rdcol_1_reset),
    .io_a(x449_rdcol_1_io_a),
    .io_b(x449_rdcol_1_io_b),
    .io_flow(x449_rdcol_1_io_flow),
    .io_result(x449_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_52 ( // @[package.scala 93:22:@45888.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x403 x453_1 ( // @[Math.scala 366:24:@45907.4]
    .clock(x453_1_clock),
    .io_a(x453_1_io_a),
    .io_flow(x453_1_io_flow),
    .io_result(x453_1_io_result)
  );
  x406_div x454_div_1 ( // @[Math.scala 327:24:@45919.4]
    .clock(x454_div_1_clock),
    .io_a(x454_div_1_io_a),
    .io_flow(x454_div_1_io_flow),
    .io_result(x454_div_1_io_result)
  );
  RetimeWrapper_358 RetimeWrapper_53 ( // @[package.scala 93:22:@45929.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x367_sum x455_sum_1 ( // @[Math.scala 150:24:@45938.4]
    .clock(x455_sum_1_clock),
    .reset(x455_sum_1_reset),
    .io_a(x455_sum_1_io_a),
    .io_b(x455_sum_1_io_b),
    .io_flow(x455_sum_1_io_flow),
    .io_result(x455_sum_1_io_result)
  );
  RetimeWrapper_360 RetimeWrapper_54 ( // @[package.scala 93:22:@45948.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_55 ( // @[package.scala 93:22:@45957.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_56 ( // @[package.scala 93:22:@45969.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x367_sum x458_rdcol_1 ( // @[Math.scala 150:24:@45992.4]
    .clock(x458_rdcol_1_clock),
    .reset(x458_rdcol_1_reset),
    .io_a(x458_rdcol_1_io_a),
    .io_b(x458_rdcol_1_io_b),
    .io_flow(x458_rdcol_1_io_flow),
    .io_result(x458_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@46007.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x403 x462_1 ( // @[Math.scala 366:24:@46024.4]
    .clock(x462_1_clock),
    .io_a(x462_1_io_a),
    .io_flow(x462_1_io_flow),
    .io_result(x462_1_io_result)
  );
  x406_div x463_div_1 ( // @[Math.scala 327:24:@46036.4]
    .clock(x463_div_1_clock),
    .io_a(x463_div_1_io_a),
    .io_flow(x463_div_1_io_flow),
    .io_result(x463_div_1_io_result)
  );
  x367_sum x464_sum_1 ( // @[Math.scala 150:24:@46046.4]
    .clock(x464_sum_1_clock),
    .reset(x464_sum_1_reset),
    .io_a(x464_sum_1_io_a),
    .io_b(x464_sum_1_io_b),
    .io_flow(x464_sum_1_io_flow),
    .io_result(x464_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_58 ( // @[package.scala 93:22:@46056.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_360 RetimeWrapper_59 ( // @[package.scala 93:22:@46065.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_60 ( // @[package.scala 93:22:@46077.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x696_sub x467_rdrow_1 ( // @[Math.scala 191:24:@46100.4]
    .clock(x467_rdrow_1_clock),
    .reset(x467_rdrow_1_reset),
    .io_a(x467_rdrow_1_io_a),
    .io_b(x467_rdrow_1_io_b),
    .io_flow(x467_rdrow_1_io_flow),
    .io_result(x467_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_61 ( // @[package.scala 93:22:@46126.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_62 ( // @[package.scala 93:22:@46148.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_63 ( // @[package.scala 93:22:@46174.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x367_sum x718_sum_1 ( // @[Math.scala 150:24:@46195.4]
    .clock(x718_sum_1_clock),
    .reset(x718_sum_1_reset),
    .io_a(x718_sum_1_io_a),
    .io_b(x718_sum_1_io_b),
    .io_flow(x718_sum_1_io_flow),
    .io_result(x718_sum_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_64 ( // @[package.scala 93:22:@46205.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_65 ( // @[package.scala 93:22:@46214.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x367_sum x475_sum_1 ( // @[Math.scala 150:24:@46223.4]
    .clock(x475_sum_1_clock),
    .reset(x475_sum_1_reset),
    .io_a(x475_sum_1_io_a),
    .io_b(x475_sum_1_io_b),
    .io_flow(x475_sum_1_io_flow),
    .io_result(x475_sum_1_io_result)
  );
  RetimeWrapper_308 RetimeWrapper_66 ( // @[package.scala 93:22:@46233.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_67 ( // @[package.scala 93:22:@46242.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_68 ( // @[package.scala 93:22:@46254.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_69 ( // @[package.scala 93:22:@46281.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x367_sum x480_sum_1 ( // @[Math.scala 150:24:@46290.4]
    .clock(x480_sum_1_clock),
    .reset(x480_sum_1_reset),
    .io_a(x480_sum_1_io_a),
    .io_b(x480_sum_1_io_b),
    .io_flow(x480_sum_1_io_flow),
    .io_result(x480_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_70 ( // @[package.scala 93:22:@46300.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_71 ( // @[package.scala 93:22:@46312.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_72 ( // @[package.scala 93:22:@46339.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x367_sum x485_sum_1 ( // @[Math.scala 150:24:@46348.4]
    .clock(x485_sum_1_clock),
    .reset(x485_sum_1_reset),
    .io_a(x485_sum_1_io_a),
    .io_b(x485_sum_1_io_b),
    .io_flow(x485_sum_1_io_flow),
    .io_result(x485_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_73 ( // @[package.scala 93:22:@46358.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_74 ( // @[package.scala 93:22:@46370.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper RetimeWrapper_75 ( // @[package.scala 93:22:@46391.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_76 ( // @[package.scala 93:22:@46406.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_390 RetimeWrapper_77 ( // @[package.scala 93:22:@46415.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x367_sum x490_sum_1 ( // @[Math.scala 150:24:@46426.4]
    .clock(x490_sum_1_clock),
    .reset(x490_sum_1_reset),
    .io_a(x490_sum_1_io_a),
    .io_b(x490_sum_1_io_b),
    .io_flow(x490_sum_1_io_flow),
    .io_result(x490_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_78 ( // @[package.scala 93:22:@46436.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_79 ( // @[package.scala 93:22:@46445.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_80 ( // @[package.scala 93:22:@46457.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x367_sum x495_sum_1 ( // @[Math.scala 150:24:@46484.4]
    .clock(x495_sum_1_clock),
    .reset(x495_sum_1_reset),
    .io_a(x495_sum_1_io_a),
    .io_b(x495_sum_1_io_b),
    .io_flow(x495_sum_1_io_flow),
    .io_result(x495_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_81 ( // @[package.scala 93:22:@46494.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_82 ( // @[package.scala 93:22:@46506.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x367_sum x500_sum_1 ( // @[Math.scala 150:24:@46533.4]
    .clock(x500_sum_1_clock),
    .reset(x500_sum_1_reset),
    .io_a(x500_sum_1_io_a),
    .io_b(x500_sum_1_io_b),
    .io_flow(x500_sum_1_io_flow),
    .io_result(x500_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_83 ( // @[package.scala 93:22:@46543.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_84 ( // @[package.scala 93:22:@46555.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  x696_sub x503_rdrow_1 ( // @[Math.scala 191:24:@46578.4]
    .clock(x503_rdrow_1_clock),
    .reset(x503_rdrow_1_reset),
    .io_a(x503_rdrow_1_io_a),
    .io_b(x503_rdrow_1_io_b),
    .io_flow(x503_rdrow_1_io_flow),
    .io_result(x503_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_85 ( // @[package.scala 93:22:@46604.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_86 ( // @[package.scala 93:22:@46626.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_87 ( // @[package.scala 93:22:@46652.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  x367_sum x723_sum_1 ( // @[Math.scala 150:24:@46673.4]
    .clock(x723_sum_1_clock),
    .reset(x723_sum_1_reset),
    .io_a(x723_sum_1_io_a),
    .io_b(x723_sum_1_io_b),
    .io_flow(x723_sum_1_io_flow),
    .io_result(x723_sum_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_88 ( // @[package.scala 93:22:@46683.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  x367_sum x511_sum_1 ( // @[Math.scala 150:24:@46692.4]
    .clock(x511_sum_1_clock),
    .reset(x511_sum_1_reset),
    .io_a(x511_sum_1_io_a),
    .io_b(x511_sum_1_io_b),
    .io_flow(x511_sum_1_io_flow),
    .io_result(x511_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_89 ( // @[package.scala 93:22:@46702.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_308 RetimeWrapper_90 ( // @[package.scala 93:22:@46711.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_91 ( // @[package.scala 93:22:@46723.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  x367_sum x516_sum_1 ( // @[Math.scala 150:24:@46750.4]
    .clock(x516_sum_1_clock),
    .reset(x516_sum_1_reset),
    .io_a(x516_sum_1_io_a),
    .io_b(x516_sum_1_io_b),
    .io_flow(x516_sum_1_io_flow),
    .io_result(x516_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_92 ( // @[package.scala 93:22:@46760.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_93 ( // @[package.scala 93:22:@46772.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  x367_sum x521_sum_1 ( // @[Math.scala 150:24:@46799.4]
    .clock(x521_sum_1_clock),
    .reset(x521_sum_1_reset),
    .io_a(x521_sum_1_io_a),
    .io_b(x521_sum_1_io_b),
    .io_flow(x521_sum_1_io_flow),
    .io_result(x521_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_94 ( // @[package.scala 93:22:@46809.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_95 ( // @[package.scala 93:22:@46821.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_390 RetimeWrapper_96 ( // @[package.scala 93:22:@46848.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  x367_sum x526_sum_1 ( // @[Math.scala 150:24:@46859.4]
    .clock(x526_sum_1_clock),
    .reset(x526_sum_1_reset),
    .io_a(x526_sum_1_io_a),
    .io_b(x526_sum_1_io_b),
    .io_flow(x526_sum_1_io_flow),
    .io_result(x526_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_97 ( // @[package.scala 93:22:@46869.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_98 ( // @[package.scala 93:22:@46878.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_99 ( // @[package.scala 93:22:@46890.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  x367_sum x531_sum_1 ( // @[Math.scala 150:24:@46917.4]
    .clock(x531_sum_1_clock),
    .reset(x531_sum_1_reset),
    .io_a(x531_sum_1_io_a),
    .io_b(x531_sum_1_io_b),
    .io_flow(x531_sum_1_io_flow),
    .io_result(x531_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_100 ( // @[package.scala 93:22:@46927.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_101 ( // @[package.scala 93:22:@46939.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  x367_sum x536_sum_1 ( // @[Math.scala 150:24:@46966.4]
    .clock(x536_sum_1_clock),
    .reset(x536_sum_1_reset),
    .io_a(x536_sum_1_io_a),
    .io_b(x536_sum_1_io_b),
    .io_flow(x536_sum_1_io_flow),
    .io_result(x536_sum_1_io_result)
  );
  RetimeWrapper_335 RetimeWrapper_102 ( // @[package.scala 93:22:@46976.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_103 ( // @[package.scala 93:22:@46988.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  x544_x13 x544_x13_1 ( // @[Math.scala 150:24:@47034.4]
    .clock(x544_x13_1_clock),
    .reset(x544_x13_1_reset),
    .io_a(x544_x13_1_io_a),
    .io_b(x544_x13_1_io_b),
    .io_flow(x544_x13_1_io_flow),
    .io_result(x544_x13_1_io_result)
  );
  x544_x13 x545_x14_1 ( // @[Math.scala 150:24:@47044.4]
    .clock(x545_x14_1_clock),
    .reset(x545_x14_1_reset),
    .io_a(x545_x14_1_io_a),
    .io_b(x545_x14_1_io_b),
    .io_flow(x545_x14_1_io_flow),
    .io_result(x545_x14_1_io_result)
  );
  x544_x13 x546_x13_1 ( // @[Math.scala 150:24:@47054.4]
    .clock(x546_x13_1_clock),
    .reset(x546_x13_1_reset),
    .io_a(x546_x13_1_io_a),
    .io_b(x546_x13_1_io_b),
    .io_flow(x546_x13_1_io_flow),
    .io_result(x546_x13_1_io_result)
  );
  x544_x13 x547_x14_1 ( // @[Math.scala 150:24:@47064.4]
    .clock(x547_x14_1_clock),
    .reset(x547_x14_1_reset),
    .io_a(x547_x14_1_io_a),
    .io_b(x547_x14_1_io_b),
    .io_flow(x547_x14_1_io_flow),
    .io_result(x547_x14_1_io_result)
  );
  x544_x13 x548_x13_1 ( // @[Math.scala 150:24:@47074.4]
    .clock(x548_x13_1_clock),
    .reset(x548_x13_1_reset),
    .io_a(x548_x13_1_io_a),
    .io_b(x548_x13_1_io_b),
    .io_flow(x548_x13_1_io_flow),
    .io_result(x548_x13_1_io_result)
  );
  x544_x13 x549_x14_1 ( // @[Math.scala 150:24:@47084.4]
    .clock(x549_x14_1_clock),
    .reset(x549_x14_1_reset),
    .io_a(x549_x14_1_io_a),
    .io_b(x549_x14_1_io_b),
    .io_flow(x549_x14_1_io_flow),
    .io_result(x549_x14_1_io_result)
  );
  x544_x13 x550_x13_1 ( // @[Math.scala 150:24:@47094.4]
    .clock(x550_x13_1_clock),
    .reset(x550_x13_1_reset),
    .io_a(x550_x13_1_io_a),
    .io_b(x550_x13_1_io_b),
    .io_flow(x550_x13_1_io_flow),
    .io_result(x550_x13_1_io_result)
  );
  RetimeWrapper_300 RetimeWrapper_104 ( // @[package.scala 93:22:@47104.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  x544_x13 x551_sum_1 ( // @[Math.scala 150:24:@47113.4]
    .clock(x551_sum_1_clock),
    .reset(x551_sum_1_reset),
    .io_a(x551_sum_1_io_a),
    .io_b(x551_sum_1_io_b),
    .io_flow(x551_sum_1_io_flow),
    .io_result(x551_sum_1_io_result)
  );
  x552 x552_1 ( // @[Math.scala 720:24:@47123.4]
    .io_b(x552_1_io_b),
    .io_result(x552_1_io_result)
  );
  x553_mul x553_mul_1 ( // @[Math.scala 262:24:@47134.4]
    .clock(x553_mul_1_clock),
    .io_a(x553_mul_1_io_a),
    .io_b(x553_mul_1_io_b),
    .io_flow(x553_mul_1_io_flow),
    .io_result(x553_mul_1_io_result)
  );
  x554 x554_1 ( // @[Math.scala 720:24:@47144.4]
    .io_b(x554_1_io_b),
    .io_result(x554_1_io_result)
  );
  RetimeWrapper_437 RetimeWrapper_105 ( // @[package.scala 93:22:@47153.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  x555_sub x555_sub_1 ( // @[Math.scala 191:24:@47162.4]
    .clock(x555_sub_1_clock),
    .reset(x555_sub_1_reset),
    .io_a(x555_sub_1_io_a),
    .io_b(x555_sub_1_io_b),
    .io_flow(x555_sub_1_io_flow),
    .io_result(x555_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_106 ( // @[package.scala 93:22:@47175.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  x555_sub x557_sub_1 ( // @[Math.scala 191:24:@47184.4]
    .clock(x557_sub_1_clock),
    .reset(x557_sub_1_reset),
    .io_a(x557_sub_1_io_a),
    .io_b(x557_sub_1_io_b),
    .io_flow(x557_sub_1_io_flow),
    .io_result(x557_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_107 ( // @[package.scala 93:22:@47197.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_108 ( // @[package.scala 93:22:@47209.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  x552 x561_1 ( // @[Math.scala 720:24:@47223.4]
    .io_b(x561_1_io_b),
    .io_result(x561_1_io_result)
  );
  x553_mul x562_mul_1 ( // @[Math.scala 262:24:@47234.4]
    .clock(x562_mul_1_clock),
    .io_a(x562_mul_1_io_a),
    .io_b(x562_mul_1_io_b),
    .io_flow(x562_mul_1_io_flow),
    .io_result(x562_mul_1_io_result)
  );
  x554 x563_1 ( // @[Math.scala 720:24:@47246.4]
    .io_b(x563_1_io_b),
    .io_result(x563_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_109 ( // @[package.scala 93:22:@47255.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  x544_x13 x564_sum_1 ( // @[Math.scala 150:24:@47264.4]
    .clock(x564_sum_1_clock),
    .reset(x564_sum_1_reset),
    .io_a(x564_sum_1_io_a),
    .io_b(x564_sum_1_io_b),
    .io_flow(x564_sum_1_io_flow),
    .io_result(x564_sum_1_io_result)
  );
  x544_x13 x570_x13_1 ( // @[Math.scala 150:24:@47299.4]
    .clock(x570_x13_1_clock),
    .reset(x570_x13_1_reset),
    .io_a(x570_x13_1_io_a),
    .io_b(x570_x13_1_io_b),
    .io_flow(x570_x13_1_io_flow),
    .io_result(x570_x13_1_io_result)
  );
  x544_x13 x571_x14_1 ( // @[Math.scala 150:24:@47309.4]
    .clock(x571_x14_1_clock),
    .reset(x571_x14_1_reset),
    .io_a(x571_x14_1_io_a),
    .io_b(x571_x14_1_io_b),
    .io_flow(x571_x14_1_io_flow),
    .io_result(x571_x14_1_io_result)
  );
  x544_x13 x572_x13_1 ( // @[Math.scala 150:24:@47319.4]
    .clock(x572_x13_1_clock),
    .reset(x572_x13_1_reset),
    .io_a(x572_x13_1_io_a),
    .io_b(x572_x13_1_io_b),
    .io_flow(x572_x13_1_io_flow),
    .io_result(x572_x13_1_io_result)
  );
  x544_x13 x573_x14_1 ( // @[Math.scala 150:24:@47329.4]
    .clock(x573_x14_1_clock),
    .reset(x573_x14_1_reset),
    .io_a(x573_x14_1_io_a),
    .io_b(x573_x14_1_io_b),
    .io_flow(x573_x14_1_io_flow),
    .io_result(x573_x14_1_io_result)
  );
  x544_x13 x574_x13_1 ( // @[Math.scala 150:24:@47339.4]
    .clock(x574_x13_1_clock),
    .reset(x574_x13_1_reset),
    .io_a(x574_x13_1_io_a),
    .io_b(x574_x13_1_io_b),
    .io_flow(x574_x13_1_io_flow),
    .io_result(x574_x13_1_io_result)
  );
  x544_x13 x575_x14_1 ( // @[Math.scala 150:24:@47349.4]
    .clock(x575_x14_1_clock),
    .reset(x575_x14_1_reset),
    .io_a(x575_x14_1_io_a),
    .io_b(x575_x14_1_io_b),
    .io_flow(x575_x14_1_io_flow),
    .io_result(x575_x14_1_io_result)
  );
  x544_x13 x576_x13_1 ( // @[Math.scala 150:24:@47359.4]
    .clock(x576_x13_1_clock),
    .reset(x576_x13_1_reset),
    .io_a(x576_x13_1_io_a),
    .io_b(x576_x13_1_io_b),
    .io_flow(x576_x13_1_io_flow),
    .io_result(x576_x13_1_io_result)
  );
  RetimeWrapper_300 RetimeWrapper_110 ( // @[package.scala 93:22:@47369.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  x544_x13 x577_sum_1 ( // @[Math.scala 150:24:@47378.4]
    .clock(x577_sum_1_clock),
    .reset(x577_sum_1_reset),
    .io_a(x577_sum_1_io_a),
    .io_b(x577_sum_1_io_b),
    .io_flow(x577_sum_1_io_flow),
    .io_result(x577_sum_1_io_result)
  );
  x552 x578_1 ( // @[Math.scala 720:24:@47388.4]
    .io_b(x578_1_io_b),
    .io_result(x578_1_io_result)
  );
  x553_mul x579_mul_1 ( // @[Math.scala 262:24:@47399.4]
    .clock(x579_mul_1_clock),
    .io_a(x579_mul_1_io_a),
    .io_b(x579_mul_1_io_b),
    .io_flow(x579_mul_1_io_flow),
    .io_result(x579_mul_1_io_result)
  );
  x554 x580_1 ( // @[Math.scala 720:24:@47409.4]
    .io_b(x580_1_io_b),
    .io_result(x580_1_io_result)
  );
  RetimeWrapper_437 RetimeWrapper_111 ( // @[package.scala 93:22:@47418.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  x555_sub x581_sub_1 ( // @[Math.scala 191:24:@47427.4]
    .clock(x581_sub_1_clock),
    .reset(x581_sub_1_reset),
    .io_a(x581_sub_1_io_a),
    .io_b(x581_sub_1_io_b),
    .io_flow(x581_sub_1_io_flow),
    .io_result(x581_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_112 ( // @[package.scala 93:22:@47440.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  x555_sub x583_sub_1 ( // @[Math.scala 191:24:@47449.4]
    .clock(x583_sub_1_clock),
    .reset(x583_sub_1_reset),
    .io_a(x583_sub_1_io_a),
    .io_b(x583_sub_1_io_b),
    .io_flow(x583_sub_1_io_flow),
    .io_result(x583_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_113 ( // @[package.scala 93:22:@47462.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_114 ( // @[package.scala 93:22:@47474.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  x552 x587_1 ( // @[Math.scala 720:24:@47488.4]
    .io_b(x587_1_io_b),
    .io_result(x587_1_io_result)
  );
  x553_mul x588_mul_1 ( // @[Math.scala 262:24:@47499.4]
    .clock(x588_mul_1_clock),
    .io_a(x588_mul_1_io_a),
    .io_b(x588_mul_1_io_b),
    .io_flow(x588_mul_1_io_flow),
    .io_result(x588_mul_1_io_result)
  );
  x554 x589_1 ( // @[Math.scala 720:24:@47509.4]
    .io_b(x589_1_io_b),
    .io_result(x589_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_115 ( // @[package.scala 93:22:@47518.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  x544_x13 x590_sum_1 ( // @[Math.scala 150:24:@47527.4]
    .clock(x590_sum_1_clock),
    .reset(x590_sum_1_reset),
    .io_a(x590_sum_1_io_a),
    .io_b(x590_sum_1_io_b),
    .io_flow(x590_sum_1_io_flow),
    .io_result(x590_sum_1_io_result)
  );
  x544_x13 x595_x13_1 ( // @[Math.scala 150:24:@47557.4]
    .clock(x595_x13_1_clock),
    .reset(x595_x13_1_reset),
    .io_a(x595_x13_1_io_a),
    .io_b(x595_x13_1_io_b),
    .io_flow(x595_x13_1_io_flow),
    .io_result(x595_x13_1_io_result)
  );
  x544_x13 x596_x14_1 ( // @[Math.scala 150:24:@47567.4]
    .clock(x596_x14_1_clock),
    .reset(x596_x14_1_reset),
    .io_a(x596_x14_1_io_a),
    .io_b(x596_x14_1_io_b),
    .io_flow(x596_x14_1_io_flow),
    .io_result(x596_x14_1_io_result)
  );
  x544_x13 x597_x13_1 ( // @[Math.scala 150:24:@47577.4]
    .clock(x597_x13_1_clock),
    .reset(x597_x13_1_reset),
    .io_a(x597_x13_1_io_a),
    .io_b(x597_x13_1_io_b),
    .io_flow(x597_x13_1_io_flow),
    .io_result(x597_x13_1_io_result)
  );
  x544_x13 x598_x14_1 ( // @[Math.scala 150:24:@47587.4]
    .clock(x598_x14_1_clock),
    .reset(x598_x14_1_reset),
    .io_a(x598_x14_1_io_a),
    .io_b(x598_x14_1_io_b),
    .io_flow(x598_x14_1_io_flow),
    .io_result(x598_x14_1_io_result)
  );
  x544_x13 x599_x13_1 ( // @[Math.scala 150:24:@47597.4]
    .clock(x599_x13_1_clock),
    .reset(x599_x13_1_reset),
    .io_a(x599_x13_1_io_a),
    .io_b(x599_x13_1_io_b),
    .io_flow(x599_x13_1_io_flow),
    .io_result(x599_x13_1_io_result)
  );
  x544_x13 x600_x14_1 ( // @[Math.scala 150:24:@47607.4]
    .clock(x600_x14_1_clock),
    .reset(x600_x14_1_reset),
    .io_a(x600_x14_1_io_a),
    .io_b(x600_x14_1_io_b),
    .io_flow(x600_x14_1_io_flow),
    .io_result(x600_x14_1_io_result)
  );
  x544_x13 x601_x13_1 ( // @[Math.scala 150:24:@47617.4]
    .clock(x601_x13_1_clock),
    .reset(x601_x13_1_reset),
    .io_a(x601_x13_1_io_a),
    .io_b(x601_x13_1_io_b),
    .io_flow(x601_x13_1_io_flow),
    .io_result(x601_x13_1_io_result)
  );
  RetimeWrapper_300 RetimeWrapper_116 ( // @[package.scala 93:22:@47627.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  x544_x13 x602_sum_1 ( // @[Math.scala 150:24:@47636.4]
    .clock(x602_sum_1_clock),
    .reset(x602_sum_1_reset),
    .io_a(x602_sum_1_io_a),
    .io_b(x602_sum_1_io_b),
    .io_flow(x602_sum_1_io_flow),
    .io_result(x602_sum_1_io_result)
  );
  x552 x603_1 ( // @[Math.scala 720:24:@47646.4]
    .io_b(x603_1_io_b),
    .io_result(x603_1_io_result)
  );
  x553_mul x604_mul_1 ( // @[Math.scala 262:24:@47657.4]
    .clock(x604_mul_1_clock),
    .io_a(x604_mul_1_io_a),
    .io_b(x604_mul_1_io_b),
    .io_flow(x604_mul_1_io_flow),
    .io_result(x604_mul_1_io_result)
  );
  x554 x605_1 ( // @[Math.scala 720:24:@47667.4]
    .io_b(x605_1_io_b),
    .io_result(x605_1_io_result)
  );
  RetimeWrapper_437 RetimeWrapper_117 ( // @[package.scala 93:22:@47676.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  x555_sub x606_sub_1 ( // @[Math.scala 191:24:@47687.4]
    .clock(x606_sub_1_clock),
    .reset(x606_sub_1_reset),
    .io_a(x606_sub_1_io_a),
    .io_b(x606_sub_1_io_b),
    .io_flow(x606_sub_1_io_flow),
    .io_result(x606_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_118 ( // @[package.scala 93:22:@47700.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  x555_sub x608_sub_1 ( // @[Math.scala 191:24:@47709.4]
    .clock(x608_sub_1_clock),
    .reset(x608_sub_1_reset),
    .io_a(x608_sub_1_io_a),
    .io_b(x608_sub_1_io_b),
    .io_flow(x608_sub_1_io_flow),
    .io_result(x608_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_119 ( // @[package.scala 93:22:@47722.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_120 ( // @[package.scala 93:22:@47734.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  x552 x612_1 ( // @[Math.scala 720:24:@47748.4]
    .io_b(x612_1_io_b),
    .io_result(x612_1_io_result)
  );
  x553_mul x613_mul_1 ( // @[Math.scala 262:24:@47759.4]
    .clock(x613_mul_1_clock),
    .io_a(x613_mul_1_io_a),
    .io_b(x613_mul_1_io_b),
    .io_flow(x613_mul_1_io_flow),
    .io_result(x613_mul_1_io_result)
  );
  x554 x614_1 ( // @[Math.scala 720:24:@47769.4]
    .io_b(x614_1_io_b),
    .io_result(x614_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_121 ( // @[package.scala 93:22:@47778.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  x544_x13 x615_sum_1 ( // @[Math.scala 150:24:@47787.4]
    .clock(x615_sum_1_clock),
    .reset(x615_sum_1_reset),
    .io_a(x615_sum_1_io_a),
    .io_b(x615_sum_1_io_b),
    .io_flow(x615_sum_1_io_flow),
    .io_result(x615_sum_1_io_result)
  );
  x544_x13 x620_x13_1 ( // @[Math.scala 150:24:@47817.4]
    .clock(x620_x13_1_clock),
    .reset(x620_x13_1_reset),
    .io_a(x620_x13_1_io_a),
    .io_b(x620_x13_1_io_b),
    .io_flow(x620_x13_1_io_flow),
    .io_result(x620_x13_1_io_result)
  );
  x544_x13 x621_x14_1 ( // @[Math.scala 150:24:@47827.4]
    .clock(x621_x14_1_clock),
    .reset(x621_x14_1_reset),
    .io_a(x621_x14_1_io_a),
    .io_b(x621_x14_1_io_b),
    .io_flow(x621_x14_1_io_flow),
    .io_result(x621_x14_1_io_result)
  );
  x544_x13 x622_x13_1 ( // @[Math.scala 150:24:@47837.4]
    .clock(x622_x13_1_clock),
    .reset(x622_x13_1_reset),
    .io_a(x622_x13_1_io_a),
    .io_b(x622_x13_1_io_b),
    .io_flow(x622_x13_1_io_flow),
    .io_result(x622_x13_1_io_result)
  );
  x544_x13 x623_x14_1 ( // @[Math.scala 150:24:@47847.4]
    .clock(x623_x14_1_clock),
    .reset(x623_x14_1_reset),
    .io_a(x623_x14_1_io_a),
    .io_b(x623_x14_1_io_b),
    .io_flow(x623_x14_1_io_flow),
    .io_result(x623_x14_1_io_result)
  );
  x544_x13 x624_x13_1 ( // @[Math.scala 150:24:@47857.4]
    .clock(x624_x13_1_clock),
    .reset(x624_x13_1_reset),
    .io_a(x624_x13_1_io_a),
    .io_b(x624_x13_1_io_b),
    .io_flow(x624_x13_1_io_flow),
    .io_result(x624_x13_1_io_result)
  );
  x544_x13 x625_x14_1 ( // @[Math.scala 150:24:@47867.4]
    .clock(x625_x14_1_clock),
    .reset(x625_x14_1_reset),
    .io_a(x625_x14_1_io_a),
    .io_b(x625_x14_1_io_b),
    .io_flow(x625_x14_1_io_flow),
    .io_result(x625_x14_1_io_result)
  );
  x544_x13 x626_x13_1 ( // @[Math.scala 150:24:@47877.4]
    .clock(x626_x13_1_clock),
    .reset(x626_x13_1_reset),
    .io_a(x626_x13_1_io_a),
    .io_b(x626_x13_1_io_b),
    .io_flow(x626_x13_1_io_flow),
    .io_result(x626_x13_1_io_result)
  );
  RetimeWrapper_300 RetimeWrapper_122 ( // @[package.scala 93:22:@47887.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  x544_x13 x627_sum_1 ( // @[Math.scala 150:24:@47896.4]
    .clock(x627_sum_1_clock),
    .reset(x627_sum_1_reset),
    .io_a(x627_sum_1_io_a),
    .io_b(x627_sum_1_io_b),
    .io_flow(x627_sum_1_io_flow),
    .io_result(x627_sum_1_io_result)
  );
  x552 x628_1 ( // @[Math.scala 720:24:@47906.4]
    .io_b(x628_1_io_b),
    .io_result(x628_1_io_result)
  );
  x553_mul x629_mul_1 ( // @[Math.scala 262:24:@47917.4]
    .clock(x629_mul_1_clock),
    .io_a(x629_mul_1_io_a),
    .io_b(x629_mul_1_io_b),
    .io_flow(x629_mul_1_io_flow),
    .io_result(x629_mul_1_io_result)
  );
  x554 x630_1 ( // @[Math.scala 720:24:@47927.4]
    .io_b(x630_1_io_b),
    .io_result(x630_1_io_result)
  );
  RetimeWrapper_437 RetimeWrapper_123 ( // @[package.scala 93:22:@47936.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  x555_sub x631_sub_1 ( // @[Math.scala 191:24:@47945.4]
    .clock(x631_sub_1_clock),
    .reset(x631_sub_1_reset),
    .io_a(x631_sub_1_io_a),
    .io_b(x631_sub_1_io_b),
    .io_flow(x631_sub_1_io_flow),
    .io_result(x631_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_124 ( // @[package.scala 93:22:@47958.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  x555_sub x633_sub_1 ( // @[Math.scala 191:24:@47967.4]
    .clock(x633_sub_1_clock),
    .reset(x633_sub_1_reset),
    .io_a(x633_sub_1_io_a),
    .io_b(x633_sub_1_io_b),
    .io_flow(x633_sub_1_io_flow),
    .io_result(x633_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_125 ( // @[package.scala 93:22:@47980.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_126 ( // @[package.scala 93:22:@47992.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  x552 x637_1 ( // @[Math.scala 720:24:@48006.4]
    .io_b(x637_1_io_b),
    .io_result(x637_1_io_result)
  );
  x553_mul x638_mul_1 ( // @[Math.scala 262:24:@48017.4]
    .clock(x638_mul_1_clock),
    .io_a(x638_mul_1_io_a),
    .io_b(x638_mul_1_io_b),
    .io_flow(x638_mul_1_io_flow),
    .io_result(x638_mul_1_io_result)
  );
  x554 x639_1 ( // @[Math.scala 720:24:@48027.4]
    .io_b(x639_1_io_b),
    .io_result(x639_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_127 ( // @[package.scala 93:22:@48036.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  x544_x13 x640_sum_1 ( // @[Math.scala 150:24:@48045.4]
    .clock(x640_sum_1_clock),
    .reset(x640_sum_1_reset),
    .io_a(x640_sum_1_io_a),
    .io_b(x640_sum_1_io_b),
    .io_flow(x640_sum_1_io_flow),
    .io_result(x640_sum_1_io_result)
  );
  RetimeWrapper_496 RetimeWrapper_128 ( // @[package.scala 93:22:@48065.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_129 ( // @[package.scala 93:22:@48074.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_130 ( // @[package.scala 93:22:@48083.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_131 ( // @[package.scala 93:22:@48092.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  assign b394 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 62:18:@44824.4]
  assign b395 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 63:18:@44825.4]
  assign _T_205 = b394 & b395; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 67:30:@44827.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 67:37:@44828.4]
  assign _T_210 = io_in_x353_TID == 8'h0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 69:76:@44833.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 69:62:@44834.4]
  assign _T_213 = io_in_x353_TDEST == 8'h0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 69:101:@44835.4]
  assign x729_x396_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@44844.4 package.scala 96:25:@44845.4]
  assign b392_number = __io_result; // @[Math.scala 723:22:@44809.4 Math.scala 724:14:@44810.4]
  assign _T_247 = $signed(b392_number); // @[Math.scala 406:49:@45009.4]
  assign _T_249 = $signed(_T_247) & $signed(32'sh3); // @[Math.scala 406:56:@45011.4]
  assign _T_250 = $signed(_T_249); // @[Math.scala 406:56:@45012.4]
  assign x709_number = $unsigned(_T_250); // @[implicits.scala 133:21:@45013.4]
  assign _T_260 = $signed(x709_number); // @[Math.scala 406:49:@45022.4]
  assign _T_262 = $signed(_T_260) & $signed(32'sh3); // @[Math.scala 406:56:@45024.4]
  assign _T_263 = $signed(_T_262); // @[Math.scala 406:56:@45025.4]
  assign _T_274 = x709_number[31]; // @[FixedPoint.scala 50:25:@45043.4]
  assign _T_278 = _T_274 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45045.4]
  assign _T_279 = x709_number[31:2]; // @[FixedPoint.scala 18:52:@45046.4]
  assign _T_285 = _T_279 == 30'h3fffffff; // @[Math.scala 451:55:@45048.4]
  assign _T_286 = x709_number[1:0]; // @[FixedPoint.scala 18:52:@45049.4]
  assign _T_292 = _T_286 != 2'h0; // @[Math.scala 451:110:@45051.4]
  assign _T_293 = _T_285 & _T_292; // @[Math.scala 451:94:@45052.4]
  assign _T_295 = {_T_278,_T_279}; // @[Cat.scala 30:58:@45054.4]
  assign x404_1_number = _T_293 ? 32'h0 : _T_295; // @[Math.scala 454:20:@45055.4]
  assign _GEN_0 = {{8'd0}, x404_1_number}; // @[Math.scala 461:32:@45060.4]
  assign _T_300 = _GEN_0 << 8; // @[Math.scala 461:32:@45060.4]
  assign _GEN_1 = {{6'd0}, x404_1_number}; // @[Math.scala 461:32:@45065.4]
  assign _T_303 = _GEN_1 << 6; // @[Math.scala 461:32:@45065.4]
  assign _T_339 = ~ io_sigsIn_break; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:101:@45163.4]
  assign _T_343 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@45171.4 package.scala 96:25:@45172.4]
  assign _T_345 = io_rr ? _T_343 : 1'h0; // @[implicits.scala 55:10:@45173.4]
  assign _T_346 = _T_339 & _T_345; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:118:@45174.4]
  assign _T_348 = _T_346 & _T_339; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:207:@45176.4]
  assign _T_349 = _T_348 & io_sigsIn_backpressure; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:226:@45177.4]
  assign x734_b394_D24 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@45142.4 package.scala 96:25:@45143.4]
  assign _T_350 = _T_349 & x734_b394_D24; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 117:252:@45178.4]
  assign x736_b395_D24 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@45160.4 package.scala 96:25:@45161.4]
  assign _T_394 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@45278.4 package.scala 96:25:@45279.4]
  assign _T_396 = io_rr ? _T_394 : 1'h0; // @[implicits.scala 55:10:@45280.4]
  assign _T_397 = _T_339 & _T_396; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:118:@45281.4]
  assign _T_399 = _T_397 & _T_339; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:207:@45283.4]
  assign _T_400 = _T_399 & io_sigsIn_backpressure; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:226:@45284.4]
  assign _T_401 = _T_400 & x734_b394_D24; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 140:252:@45285.4]
  assign _T_442 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@45376.4 package.scala 96:25:@45377.4]
  assign _T_444 = io_rr ? _T_442 : 1'h0; // @[implicits.scala 55:10:@45378.4]
  assign _T_445 = _T_339 & _T_444; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:118:@45379.4]
  assign _T_447 = _T_445 & _T_339; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:207:@45381.4]
  assign _T_448 = _T_447 & io_sigsIn_backpressure; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:226:@45382.4]
  assign _T_449 = _T_448 & x734_b394_D24; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 161:252:@45383.4]
  assign _T_490 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@45474.4 package.scala 96:25:@45475.4]
  assign _T_492 = io_rr ? _T_490 : 1'h0; // @[implicits.scala 55:10:@45476.4]
  assign _T_493 = _T_339 & _T_492; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:166:@45477.4]
  assign _T_495 = _T_493 & _T_339; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:255:@45479.4]
  assign _T_496 = _T_495 & io_sigsIn_backpressure; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:274:@45480.4]
  assign _T_497 = _T_496 & x734_b394_D24; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 188:300:@45481.4]
  assign x747_b392_D26_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@45495.4 package.scala 96:25:@45496.4]
  assign _T_509 = $signed(x747_b392_D26_number); // @[Math.scala 476:37:@45503.4]
  assign x748_x421_rdcol_D26_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@45520.4 package.scala 96:25:@45521.4]
  assign _T_522 = $signed(x748_x421_rdcol_D26_number); // @[Math.scala 476:37:@45526.4]
  assign x749_x428_D1 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@45543.4 package.scala 96:25:@45544.4]
  assign x429 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@45534.4 package.scala 96:25:@45535.4]
  assign x430 = x749_x428_D1 | x429; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 203:24:@45547.4]
  assign _T_563 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@45615.4 package.scala 96:25:@45616.4]
  assign _T_565 = io_rr ? _T_563 : 1'h0; // @[implicits.scala 55:10:@45617.4]
  assign _T_566 = _T_339 & _T_565; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 222:194:@45618.4]
  assign x754_x431_D20 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@45594.4 package.scala 96:25:@45595.4]
  assign _T_567 = _T_566 & x754_x431_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 222:283:@45619.4]
  assign x753_b394_D48 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@45585.4 package.scala 96:25:@45586.4]
  assign _T_568 = _T_567 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 222:291:@45620.4]
  assign x755_b395_D48 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@45603.4 package.scala 96:25:@45604.4]
  assign x756_x415_rdcol_D26_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@45636.4 package.scala 96:25:@45637.4]
  assign _T_579 = $signed(x756_x415_rdcol_D26_number); // @[Math.scala 476:37:@45642.4]
  assign x434 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@45650.4 package.scala 96:25:@45651.4]
  assign x435 = x749_x428_D1 | x434; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 230:24:@45654.4]
  assign _T_608 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@45695.4 package.scala 96:25:@45696.4]
  assign _T_610 = io_rr ? _T_608 : 1'h0; // @[implicits.scala 55:10:@45697.4]
  assign _T_611 = _T_339 & _T_610; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:194:@45698.4]
  assign x758_x436_D20 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@45674.4 package.scala 96:25:@45675.4]
  assign _T_612 = _T_611 & x758_x436_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:283:@45699.4]
  assign _T_613 = _T_612 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:291:@45700.4]
  assign x760_x409_rdcol_D26_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@45716.4 package.scala 96:25:@45717.4]
  assign _T_624 = $signed(x760_x409_rdcol_D26_number); // @[Math.scala 476:37:@45722.4]
  assign x439 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@45730.4 package.scala 96:25:@45731.4]
  assign x440 = x749_x428_D1 | x439; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 251:24:@45734.4]
  assign _T_653 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@45775.4 package.scala 96:25:@45776.4]
  assign _T_655 = io_rr ? _T_653 : 1'h0; // @[implicits.scala 55:10:@45777.4]
  assign _T_656 = _T_339 & _T_655; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:194:@45778.4]
  assign x763_x441_D20 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@45763.4 package.scala 96:25:@45764.4]
  assign _T_657 = _T_656 & x763_x441_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:283:@45779.4]
  assign _T_658 = _T_657 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:291:@45780.4]
  assign x764_b393_D26_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@45796.4 package.scala 96:25:@45797.4]
  assign _T_669 = $signed(x764_b393_D26_number); // @[Math.scala 476:37:@45802.4]
  assign x428 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@45511.4 package.scala 96:25:@45512.4]
  assign x444 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@45810.4 package.scala 96:25:@45811.4]
  assign x445 = x428 | x444; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 272:24:@45814.4]
  assign _T_698 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@45855.4 package.scala 96:25:@45856.4]
  assign _T_700 = io_rr ? _T_698 : 1'h0; // @[implicits.scala 55:10:@45857.4]
  assign _T_701 = _T_339 & _T_700; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:194:@45858.4]
  assign x767_x446_D21 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@45843.4 package.scala 96:25:@45844.4]
  assign _T_702 = _T_701 & x767_x446_D21; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:283:@45859.4]
  assign _T_703 = _T_702 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:291:@45860.4]
  assign x449_rdcol_number = x449_rdcol_1_io_result; // @[Math.scala 154:22:@45879.4 Math.scala 155:14:@45880.4]
  assign _T_718 = $signed(x449_rdcol_number); // @[Math.scala 476:37:@45885.4]
  assign x450 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@45893.4 package.scala 96:25:@45894.4]
  assign x451 = x749_x428_D1 | x450; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 293:24:@45897.4]
  assign _T_766 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@45974.4 package.scala 96:25:@45975.4]
  assign _T_768 = io_rr ? _T_766 : 1'h0; // @[implicits.scala 55:10:@45976.4]
  assign _T_769 = _T_339 & _T_768; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:194:@45977.4]
  assign x770_x452_D20 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@45962.4 package.scala 96:25:@45963.4]
  assign _T_770 = _T_769 & x770_x452_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:283:@45978.4]
  assign _T_771 = _T_770 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:291:@45979.4]
  assign x458_rdcol_number = x458_rdcol_1_io_result; // @[Math.scala 154:22:@45998.4 Math.scala 155:14:@45999.4]
  assign _T_786 = $signed(x458_rdcol_number); // @[Math.scala 476:37:@46004.4]
  assign x459 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@46012.4 package.scala 96:25:@46013.4]
  assign x460 = x749_x428_D1 | x459; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 328:59:@46016.4]
  assign _T_829 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@46082.4 package.scala 96:25:@46083.4]
  assign _T_831 = io_rr ? _T_829 : 1'h0; // @[implicits.scala 55:10:@46084.4]
  assign _T_832 = _T_339 & _T_831; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 345:194:@46085.4]
  assign x771_x461_D20 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@46061.4 package.scala 96:25:@46062.4]
  assign _T_833 = _T_832 & x771_x461_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 345:283:@46086.4]
  assign _T_834 = _T_833 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 345:291:@46087.4]
  assign x467_rdrow_number = x467_rdrow_1_io_result; // @[Math.scala 195:22:@46106.4 Math.scala 196:14:@46107.4]
  assign _T_851 = $signed(x467_rdrow_number); // @[Math.scala 406:49:@46113.4]
  assign _T_853 = $signed(_T_851) & $signed(32'sh3); // @[Math.scala 406:56:@46115.4]
  assign _T_854 = $signed(_T_853); // @[Math.scala 406:56:@46116.4]
  assign x714_number = $unsigned(_T_854); // @[implicits.scala 133:21:@46117.4]
  assign x469 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@46131.4 package.scala 96:25:@46132.4]
  assign x470 = x469 | x429; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 355:24:@46135.4]
  assign _T_877 = $signed(x714_number); // @[Math.scala 406:49:@46144.4]
  assign _T_879 = $signed(_T_877) & $signed(32'sh3); // @[Math.scala 406:56:@46146.4]
  assign _T_880 = $signed(_T_879); // @[Math.scala 406:56:@46147.4]
  assign _T_884 = $signed(RetimeWrapper_62_io_out); // @[package.scala 96:25:@46155.4]
  assign _T_888 = x714_number[31]; // @[FixedPoint.scala 50:25:@46162.4]
  assign _T_892 = _T_888 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@46164.4]
  assign _T_893 = x714_number[31:2]; // @[FixedPoint.scala 18:52:@46165.4]
  assign _T_899 = _T_893 == 30'h3fffffff; // @[Math.scala 451:55:@46167.4]
  assign _T_900 = x714_number[1:0]; // @[FixedPoint.scala 18:52:@46168.4]
  assign _T_906 = _T_900 != 2'h0; // @[Math.scala 451:110:@46170.4]
  assign _T_907 = _T_899 & _T_906; // @[Math.scala 451:94:@46171.4]
  assign _T_911 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@46179.4 package.scala 96:25:@46180.4]
  assign x473_1_number = _T_907 ? 32'h0 : _T_911; // @[Math.scala 454:20:@46181.4]
  assign _GEN_2 = {{8'd0}, x473_1_number}; // @[Math.scala 461:32:@46186.4]
  assign _T_916 = _GEN_2 << 8; // @[Math.scala 461:32:@46186.4]
  assign _GEN_3 = {{6'd0}, x473_1_number}; // @[Math.scala 461:32:@46191.4]
  assign _T_919 = _GEN_3 << 6; // @[Math.scala 461:32:@46191.4]
  assign _T_949 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@46259.4 package.scala 96:25:@46260.4]
  assign _T_951 = io_rr ? _T_949 : 1'h0; // @[implicits.scala 55:10:@46261.4]
  assign _T_952 = _T_339 & _T_951; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:194:@46262.4]
  assign x776_x471_D20 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@46247.4 package.scala 96:25:@46248.4]
  assign _T_953 = _T_952 & x776_x471_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:283:@46263.4]
  assign _T_954 = _T_953 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:291:@46264.4]
  assign x478 = x469 | x434; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 386:24:@46275.4]
  assign _T_981 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@46317.4 package.scala 96:25:@46318.4]
  assign _T_983 = io_rr ? _T_981 : 1'h0; // @[implicits.scala 55:10:@46319.4]
  assign _T_984 = _T_339 & _T_983; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:194:@46320.4]
  assign x778_x479_D20 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@46305.4 package.scala 96:25:@46306.4]
  assign _T_985 = _T_984 & x778_x479_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:283:@46321.4]
  assign _T_986 = _T_985 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:291:@46322.4]
  assign x483 = x469 | x439; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 403:24:@46333.4]
  assign _T_1013 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@46375.4 package.scala 96:25:@46376.4]
  assign _T_1015 = io_rr ? _T_1013 : 1'h0; // @[implicits.scala 55:10:@46377.4]
  assign _T_1016 = _T_339 & _T_1015; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:194:@46378.4]
  assign x780_x484_D20 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@46363.4 package.scala 96:25:@46364.4]
  assign _T_1017 = _T_1016 & x780_x484_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:283:@46379.4]
  assign _T_1018 = _T_1017 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:291:@46380.4]
  assign x781_x444_D1 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@46396.4 package.scala 96:25:@46397.4]
  assign x488 = x469 | x781_x444_D1; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 428:59:@46400.4]
  assign _T_1056 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@46462.4 package.scala 96:25:@46463.4]
  assign _T_1058 = io_rr ? _T_1056 : 1'h0; // @[implicits.scala 55:10:@46464.4]
  assign _T_1059 = _T_339 & _T_1058; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:194:@46465.4]
  assign x784_x489_D20 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@46441.4 package.scala 96:25:@46442.4]
  assign _T_1060 = _T_1059 & x784_x489_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:283:@46466.4]
  assign _T_1061 = _T_1060 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:291:@46467.4]
  assign x493 = x469 | x450; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 451:59:@46478.4]
  assign _T_1085 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@46511.4 package.scala 96:25:@46512.4]
  assign _T_1087 = io_rr ? _T_1085 : 1'h0; // @[implicits.scala 55:10:@46513.4]
  assign _T_1088 = _T_339 & _T_1087; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:194:@46514.4]
  assign x786_x494_D20 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@46499.4 package.scala 96:25:@46500.4]
  assign _T_1089 = _T_1088 & x786_x494_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:283:@46515.4]
  assign _T_1090 = _T_1089 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:291:@46516.4]
  assign x498 = x469 | x459; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 466:59:@46527.4]
  assign _T_1114 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@46560.4 package.scala 96:25:@46561.4]
  assign _T_1116 = io_rr ? _T_1114 : 1'h0; // @[implicits.scala 55:10:@46562.4]
  assign _T_1117 = _T_339 & _T_1116; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:194:@46563.4]
  assign x787_x499_D20 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@46548.4 package.scala 96:25:@46549.4]
  assign _T_1118 = _T_1117 & x787_x499_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:283:@46564.4]
  assign _T_1119 = _T_1118 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:291:@46565.4]
  assign x503_rdrow_number = x503_rdrow_1_io_result; // @[Math.scala 195:22:@46584.4 Math.scala 196:14:@46585.4]
  assign _T_1136 = $signed(x503_rdrow_number); // @[Math.scala 406:49:@46591.4]
  assign _T_1138 = $signed(_T_1136) & $signed(32'sh3); // @[Math.scala 406:56:@46593.4]
  assign _T_1139 = $signed(_T_1138); // @[Math.scala 406:56:@46594.4]
  assign x719_number = $unsigned(_T_1139); // @[implicits.scala 133:21:@46595.4]
  assign x505 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@46609.4 package.scala 96:25:@46610.4]
  assign x506 = x505 | x429; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 487:24:@46613.4]
  assign _T_1162 = $signed(x719_number); // @[Math.scala 406:49:@46622.4]
  assign _T_1164 = $signed(_T_1162) & $signed(32'sh3); // @[Math.scala 406:56:@46624.4]
  assign _T_1165 = $signed(_T_1164); // @[Math.scala 406:56:@46625.4]
  assign _T_1169 = $signed(RetimeWrapper_86_io_out); // @[package.scala 96:25:@46633.4]
  assign _T_1173 = x719_number[31]; // @[FixedPoint.scala 50:25:@46640.4]
  assign _T_1177 = _T_1173 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@46642.4]
  assign _T_1178 = x719_number[31:2]; // @[FixedPoint.scala 18:52:@46643.4]
  assign _T_1184 = _T_1178 == 30'h3fffffff; // @[Math.scala 451:55:@46645.4]
  assign _T_1185 = x719_number[1:0]; // @[FixedPoint.scala 18:52:@46646.4]
  assign _T_1191 = _T_1185 != 2'h0; // @[Math.scala 451:110:@46648.4]
  assign _T_1192 = _T_1184 & _T_1191; // @[Math.scala 451:94:@46649.4]
  assign _T_1196 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@46657.4 package.scala 96:25:@46658.4]
  assign x509_1_number = _T_1192 ? 32'h0 : _T_1196; // @[Math.scala 454:20:@46659.4]
  assign _GEN_4 = {{8'd0}, x509_1_number}; // @[Math.scala 461:32:@46664.4]
  assign _T_1201 = _GEN_4 << 8; // @[Math.scala 461:32:@46664.4]
  assign _GEN_5 = {{6'd0}, x509_1_number}; // @[Math.scala 461:32:@46669.4]
  assign _T_1204 = _GEN_5 << 6; // @[Math.scala 461:32:@46669.4]
  assign _T_1231 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@46728.4 package.scala 96:25:@46729.4]
  assign _T_1233 = io_rr ? _T_1231 : 1'h0; // @[implicits.scala 55:10:@46730.4]
  assign _T_1234 = _T_339 & _T_1233; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 512:194:@46731.4]
  assign x789_x507_D20 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@46707.4 package.scala 96:25:@46708.4]
  assign _T_1235 = _T_1234 & x789_x507_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 512:283:@46732.4]
  assign _T_1236 = _T_1235 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 512:291:@46733.4]
  assign x514 = x505 | x434; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 516:24:@46744.4]
  assign _T_1260 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@46777.4 package.scala 96:25:@46778.4]
  assign _T_1262 = io_rr ? _T_1260 : 1'h0; // @[implicits.scala 55:10:@46779.4]
  assign _T_1263 = _T_339 & _T_1262; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:194:@46780.4]
  assign x791_x515_D20 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@46765.4 package.scala 96:25:@46766.4]
  assign _T_1264 = _T_1263 & x791_x515_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:283:@46781.4]
  assign _T_1265 = _T_1264 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:291:@46782.4]
  assign x519 = x505 | x439; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 531:24:@46793.4]
  assign _T_1289 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@46826.4 package.scala 96:25:@46827.4]
  assign _T_1291 = io_rr ? _T_1289 : 1'h0; // @[implicits.scala 55:10:@46828.4]
  assign _T_1292 = _T_339 & _T_1291; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:194:@46829.4]
  assign x792_x520_D20 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@46814.4 package.scala 96:25:@46815.4]
  assign _T_1293 = _T_1292 & x792_x520_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:283:@46830.4]
  assign _T_1294 = _T_1293 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:326:@46831.4]
  assign x524 = x505 | x781_x444_D1; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 552:59:@46842.4]
  assign _T_1326 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@46895.4 package.scala 96:25:@46896.4]
  assign _T_1328 = io_rr ? _T_1326 : 1'h0; // @[implicits.scala 55:10:@46897.4]
  assign _T_1329 = _T_339 & _T_1328; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:194:@46898.4]
  assign x795_x525_D20 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@46883.4 package.scala 96:25:@46884.4]
  assign _T_1330 = _T_1329 & x795_x525_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:283:@46899.4]
  assign _T_1331 = _T_1330 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:291:@46900.4]
  assign x529 = x505 | x450; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 573:59:@46911.4]
  assign _T_1355 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@46944.4 package.scala 96:25:@46945.4]
  assign _T_1357 = io_rr ? _T_1355 : 1'h0; // @[implicits.scala 55:10:@46946.4]
  assign _T_1358 = _T_339 & _T_1357; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:194:@46947.4]
  assign x796_x530_D20 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@46932.4 package.scala 96:25:@46933.4]
  assign _T_1359 = _T_1358 & x796_x530_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:283:@46948.4]
  assign _T_1360 = _T_1359 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:291:@46949.4]
  assign x534 = x505 | x459; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 588:59:@46960.4]
  assign _T_1384 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@46993.4 package.scala 96:25:@46994.4]
  assign _T_1386 = io_rr ? _T_1384 : 1'h0; // @[implicits.scala 55:10:@46995.4]
  assign _T_1387 = _T_339 & _T_1386; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 599:194:@46996.4]
  assign x797_x535_D20 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@46981.4 package.scala 96:25:@46982.4]
  assign _T_1388 = _T_1387 & x797_x535_D20; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 599:283:@46997.4]
  assign _T_1389 = _T_1388 & x753_b394_D48; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 599:291:@46998.4]
  assign x437_rd_0_number = x398_lb_0_io_rPort_11_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 239:29:@45686.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 243:338:@45707.4]
  assign _GEN_6 = {{1'd0}, x437_rd_0_number}; // @[Math.scala 461:32:@47010.4]
  assign _T_1394 = _GEN_6 << 1; // @[Math.scala 461:32:@47010.4]
  assign x476_rd_0_number = x398_lb_0_io_rPort_6_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 378:29:@46250.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 382:408:@46271.4]
  assign _GEN_7 = {{1'd0}, x476_rd_0_number}; // @[Math.scala 461:32:@47015.4]
  assign _T_1397 = _GEN_7 << 1; // @[Math.scala 461:32:@47015.4]
  assign x481_rd_0_number = x398_lb_0_io_rPort_0_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 395:29:@46308.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 399:408:@46329.4]
  assign _GEN_8 = {{2'd0}, x481_rd_0_number}; // @[Math.scala 461:32:@47020.4]
  assign _T_1400 = _GEN_8 << 2; // @[Math.scala 461:32:@47020.4]
  assign x486_rd_0_number = x398_lb_0_io_rPort_15_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 412:29:@46366.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 416:408:@46387.4]
  assign _GEN_9 = {{1'd0}, x486_rd_0_number}; // @[Math.scala 461:32:@47025.4]
  assign _T_1403 = _GEN_9 << 1; // @[Math.scala 461:32:@47025.4]
  assign x517_rd_0_number = x398_lb_0_io_rPort_8_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 523:29:@46768.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 527:408:@46789.4]
  assign _GEN_10 = {{1'd0}, x517_rd_0_number}; // @[Math.scala 461:32:@47030.4]
  assign _T_1406 = _GEN_10 << 1; // @[Math.scala 461:32:@47030.4]
  assign x555_sub_number = x555_sub_1_io_result; // @[Math.scala 195:22:@47168.4 Math.scala 196:14:@47169.4]
  assign x557_sub_number = x557_sub_1_io_result; // @[Math.scala 195:22:@47190.4 Math.scala 196:14:@47191.4]
  assign x556 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@47180.4 package.scala 96:25:@47181.4]
  assign x558 = RetimeWrapper_107_io_out; // @[package.scala 96:25:@47202.4 package.scala 96:25:@47203.4]
  assign x559 = x556 | x558; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 647:24:@47206.4]
  assign x800_x555_sub_D1_number = RetimeWrapper_108_io_out; // @[package.scala 96:25:@47214.4 package.scala 96:25:@47215.4]
  assign x442_rd_0_number = x398_lb_0_io_rPort_13_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 260:29:@45766.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 264:338:@45787.4]
  assign _GEN_11 = {{1'd0}, x442_rd_0_number}; // @[Math.scala 461:32:@47275.4]
  assign _T_1506 = _GEN_11 << 1; // @[Math.scala 461:32:@47275.4]
  assign _GEN_12 = {{1'd0}, x481_rd_0_number}; // @[Math.scala 461:32:@47280.4]
  assign _T_1509 = _GEN_12 << 1; // @[Math.scala 461:32:@47280.4]
  assign _GEN_13 = {{2'd0}, x486_rd_0_number}; // @[Math.scala 461:32:@47285.4]
  assign _T_1512 = _GEN_13 << 2; // @[Math.scala 461:32:@47285.4]
  assign x491_rd_0_number = x398_lb_0_io_rPort_16_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 443:29:@46453.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 447:408:@46474.4]
  assign _GEN_14 = {{1'd0}, x491_rd_0_number}; // @[Math.scala 461:32:@47290.4]
  assign _T_1515 = _GEN_14 << 1; // @[Math.scala 461:32:@47290.4]
  assign x522_rd_0_number = x398_lb_0_io_rPort_3_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 544:29:@46817.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 548:443:@46838.4]
  assign _GEN_15 = {{1'd0}, x522_rd_0_number}; // @[Math.scala 461:32:@47295.4]
  assign _T_1518 = _GEN_15 << 1; // @[Math.scala 461:32:@47295.4]
  assign x581_sub_number = x581_sub_1_io_result; // @[Math.scala 195:22:@47433.4 Math.scala 196:14:@47434.4]
  assign x583_sub_number = x583_sub_1_io_result; // @[Math.scala 195:22:@47455.4 Math.scala 196:14:@47456.4]
  assign x582 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@47445.4 package.scala 96:25:@47446.4]
  assign x584 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@47467.4 package.scala 96:25:@47468.4]
  assign x585 = x582 | x584; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 715:24:@47471.4]
  assign x804_x581_sub_D1_number = RetimeWrapper_114_io_out; // @[package.scala 96:25:@47479.4 package.scala 96:25:@47480.4]
  assign x447_rd_0_number = x398_lb_0_io_rPort_9_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 281:29:@45846.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 285:338:@45867.4]
  assign _GEN_16 = {{1'd0}, x447_rd_0_number}; // @[Math.scala 461:32:@47538.4]
  assign _T_1616 = _GEN_16 << 1; // @[Math.scala 461:32:@47538.4]
  assign _GEN_17 = {{2'd0}, x491_rd_0_number}; // @[Math.scala 461:32:@47543.4]
  assign _T_1619 = _GEN_17 << 2; // @[Math.scala 461:32:@47543.4]
  assign x496_rd_0_number = x398_lb_0_io_rPort_17_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 458:29:@46502.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 462:408:@46523.4]
  assign _GEN_18 = {{1'd0}, x496_rd_0_number}; // @[Math.scala 461:32:@47548.4]
  assign _T_1622 = _GEN_18 << 1; // @[Math.scala 461:32:@47548.4]
  assign x527_rd_0_number = x398_lb_0_io_rPort_1_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 565:29:@46886.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 569:408:@46907.4]
  assign _GEN_19 = {{1'd0}, x527_rd_0_number}; // @[Math.scala 461:32:@47553.4]
  assign _T_1625 = _GEN_19 << 1; // @[Math.scala 461:32:@47553.4]
  assign x606_sub_number = x606_sub_1_io_result; // @[Math.scala 195:22:@47693.4 Math.scala 196:14:@47694.4]
  assign x608_sub_number = x608_sub_1_io_result; // @[Math.scala 195:22:@47715.4 Math.scala 196:14:@47716.4]
  assign x607 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@47705.4 package.scala 96:25:@47706.4]
  assign x609 = RetimeWrapper_119_io_out; // @[package.scala 96:25:@47727.4 package.scala 96:25:@47728.4]
  assign x610 = x607 | x609; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 781:24:@47731.4]
  assign x808_x606_sub_D1_number = RetimeWrapper_120_io_out; // @[package.scala 96:25:@47739.4 package.scala 96:25:@47740.4]
  assign x456_rd_0_number = x398_lb_0_io_rPort_4_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 316:29:@45965.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 320:408:@45986.4]
  assign _GEN_20 = {{1'd0}, x456_rd_0_number}; // @[Math.scala 461:32:@47798.4]
  assign _T_1725 = _GEN_20 << 1; // @[Math.scala 461:32:@47798.4]
  assign _GEN_21 = {{2'd0}, x496_rd_0_number}; // @[Math.scala 461:32:@47803.4]
  assign _T_1728 = _GEN_21 << 2; // @[Math.scala 461:32:@47803.4]
  assign x501_rd_0_number = x398_lb_0_io_rPort_14_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 473:29:@46551.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 477:408:@46572.4]
  assign _GEN_22 = {{1'd0}, x501_rd_0_number}; // @[Math.scala 461:32:@47808.4]
  assign _T_1731 = _GEN_22 << 1; // @[Math.scala 461:32:@47808.4]
  assign x532_rd_0_number = x398_lb_0_io_rPort_12_output_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 580:29:@46935.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 584:408:@46956.4]
  assign _GEN_23 = {{1'd0}, x532_rd_0_number}; // @[Math.scala 461:32:@47813.4]
  assign _T_1734 = _GEN_23 << 1; // @[Math.scala 461:32:@47813.4]
  assign x631_sub_number = x631_sub_1_io_result; // @[Math.scala 195:22:@47951.4 Math.scala 196:14:@47952.4]
  assign x633_sub_number = x633_sub_1_io_result; // @[Math.scala 195:22:@47973.4 Math.scala 196:14:@47974.4]
  assign x632 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@47963.4 package.scala 96:25:@47964.4]
  assign x634 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@47985.4 package.scala 96:25:@47986.4]
  assign x635 = x632 | x634; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 839:24:@47989.4]
  assign x812_x631_sub_D1_number = RetimeWrapper_126_io_out; // @[package.scala 96:25:@47997.4 package.scala 96:25:@47998.4]
  assign x615_sum_number = x615_sum_1_io_result; // @[Math.scala 154:22:@47793.4 Math.scala 155:14:@47794.4]
  assign x640_sum_number = x640_sum_1_io_result; // @[Math.scala 154:22:@48051.4 Math.scala 155:14:@48052.4]
  assign _T_1841 = {x615_sum_number,x640_sum_number}; // @[Cat.scala 30:58:@48060.4]
  assign x564_sum_number = x564_sum_1_io_result; // @[Math.scala 154:22:@47270.4 Math.scala 155:14:@47271.4]
  assign x590_sum_number = x590_sum_1_io_result; // @[Math.scala 154:22:@47533.4 Math.scala 155:14:@47534.4]
  assign _T_1842 = {x564_sum_number,x590_sum_number}; // @[Cat.scala 30:58:@48061.4]
  assign _T_1855 = RetimeWrapper_131_io_out; // @[package.scala 96:25:@48097.4 package.scala 96:25:@48098.4]
  assign _T_1857 = io_rr ? _T_1855 : 1'h0; // @[implicits.scala 55:10:@48099.4]
  assign x815_b394_D72 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@48088.4 package.scala 96:25:@48089.4]
  assign _T_1858 = _T_1857 & x815_b394_D72; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 863:117:@48100.4]
  assign x814_b395_D72 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@48079.4 package.scala 96:25:@48080.4]
  assign _T_1859 = _T_1858 & x814_b395_D72; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 863:123:@48101.4]
  assign x731_x407_sum_D3_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@45115.4 package.scala 96:25:@45116.4]
  assign x732_x710_D24_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@45124.4 package.scala 96:25:@45125.4]
  assign x733_x403_D8_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@45133.4 package.scala 96:25:@45134.4]
  assign x738_x411_D7_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@45249.4 package.scala 96:25:@45250.4]
  assign x739_x413_sum_D2_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@45258.4 package.scala 96:25:@45259.4]
  assign x741_x417_D7_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@45347.4 package.scala 96:25:@45348.4]
  assign x743_x419_sum_D2_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@45365.4 package.scala 96:25:@45366.4]
  assign x744_x425_sum_D2_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@45445.4 package.scala 96:25:@45446.4]
  assign x745_x423_D7_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@45454.4 package.scala 96:25:@45455.4]
  assign x750_x710_D48_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@45558.4 package.scala 96:25:@45559.4]
  assign x751_x425_sum_D26_number = RetimeWrapper_28_io_out; // @[package.scala 96:25:@45567.4 package.scala 96:25:@45568.4]
  assign x752_x423_D31_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@45576.4 package.scala 96:25:@45577.4]
  assign x757_x417_D31_number = RetimeWrapper_36_io_out; // @[package.scala 96:25:@45665.4 package.scala 96:25:@45666.4]
  assign x759_x419_sum_D26_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@45683.4 package.scala 96:25:@45684.4]
  assign x761_x411_D31_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@45745.4 package.scala 96:25:@45746.4]
  assign x762_x413_sum_D26_number = RetimeWrapper_43_io_out; // @[package.scala 96:25:@45754.4 package.scala 96:25:@45755.4]
  assign x765_x407_sum_D27_number = RetimeWrapper_48_io_out; // @[package.scala 96:25:@45825.4 package.scala 96:25:@45826.4]
  assign x766_x403_D32_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@45834.4 package.scala 96:25:@45835.4]
  assign x455_sum_number = x455_sum_1_io_result; // @[Math.scala 154:22:@45944.4 Math.scala 155:14:@45945.4]
  assign x769_x453_D5_number = RetimeWrapper_54_io_out; // @[package.scala 96:25:@45953.4 package.scala 96:25:@45954.4]
  assign x464_sum_number = x464_sum_1_io_result; // @[Math.scala 154:22:@46052.4 Math.scala 155:14:@46053.4]
  assign x772_x462_D5_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@46070.4 package.scala 96:25:@46071.4]
  assign x475_sum_number = x475_sum_1_io_result; // @[Math.scala 154:22:@46229.4 Math.scala 155:14:@46230.4]
  assign x775_x715_D20_number = RetimeWrapper_66_io_out; // @[package.scala 96:25:@46238.4 package.scala 96:25:@46239.4]
  assign x480_sum_number = x480_sum_1_io_result; // @[Math.scala 154:22:@46296.4 Math.scala 155:14:@46297.4]
  assign x485_sum_number = x485_sum_1_io_result; // @[Math.scala 154:22:@46354.4 Math.scala 155:14:@46355.4]
  assign x785_x490_sum_D1_number = RetimeWrapper_79_io_out; // @[package.scala 96:25:@46450.4 package.scala 96:25:@46451.4]
  assign x495_sum_number = x495_sum_1_io_result; // @[Math.scala 154:22:@46490.4 Math.scala 155:14:@46491.4]
  assign x500_sum_number = x500_sum_1_io_result; // @[Math.scala 154:22:@46539.4 Math.scala 155:14:@46540.4]
  assign x511_sum_number = x511_sum_1_io_result; // @[Math.scala 154:22:@46698.4 Math.scala 155:14:@46699.4]
  assign x790_x720_D20_number = RetimeWrapper_90_io_out; // @[package.scala 96:25:@46716.4 package.scala 96:25:@46717.4]
  assign x516_sum_number = x516_sum_1_io_result; // @[Math.scala 154:22:@46756.4 Math.scala 155:14:@46757.4]
  assign x521_sum_number = x521_sum_1_io_result; // @[Math.scala 154:22:@46805.4 Math.scala 155:14:@46806.4]
  assign x794_x526_sum_D1_number = RetimeWrapper_97_io_out; // @[package.scala 96:25:@46874.4 package.scala 96:25:@46875.4]
  assign x531_sum_number = x531_sum_1_io_result; // @[Math.scala 154:22:@46923.4 Math.scala 155:14:@46924.4]
  assign x536_sum_number = x536_sum_1_io_result; // @[Math.scala 154:22:@46972.4 Math.scala 155:14:@46973.4]
  assign io_in_x353_TREADY = _T_211 & _T_213; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 67:22:@44829.4 sm_x645_inr_Foreach_SAMPLER_BOX.scala 69:22:@44837.4]
  assign io_in_x354_TVALID = _T_1859 & io_sigsIn_backpressure; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 863:22:@48103.4]
  assign io_in_x354_TDATA = {{128'd0}, RetimeWrapper_128_io_out}; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 864:24:@48104.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@44807.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@44819.4]
  assign RetimeWrapper_clock = clock; // @[:@44840.4]
  assign RetimeWrapper_reset = reset; // @[:@44841.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44843.4]
  assign RetimeWrapper_io_in = io_in_x353_TDATA[127:0]; // @[package.scala 94:16:@44842.4]
  assign x398_lb_0_clock = clock; // @[:@44850.4]
  assign x398_lb_0_reset = reset; // @[:@44851.4]
  assign x398_lb_0_io_rPort_17_banks_1 = x769_x453_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@46519.4]
  assign x398_lb_0_io_rPort_17_banks_0 = x775_x715_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46518.4]
  assign x398_lb_0_io_rPort_17_ofs_0 = x495_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46520.4]
  assign x398_lb_0_io_rPort_17_en_0 = _T_1090 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46522.4]
  assign x398_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46521.4]
  assign x398_lb_0_io_rPort_16_banks_1 = x766_x403_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@46470.4]
  assign x398_lb_0_io_rPort_16_banks_0 = x775_x715_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46469.4]
  assign x398_lb_0_io_rPort_16_ofs_0 = x785_x490_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@46471.4]
  assign x398_lb_0_io_rPort_16_en_0 = _T_1061 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46473.4]
  assign x398_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46472.4]
  assign x398_lb_0_io_rPort_15_banks_1 = x761_x411_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@46383.4]
  assign x398_lb_0_io_rPort_15_banks_0 = x775_x715_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46382.4]
  assign x398_lb_0_io_rPort_15_ofs_0 = x485_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46384.4]
  assign x398_lb_0_io_rPort_15_en_0 = _T_1018 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46386.4]
  assign x398_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46385.4]
  assign x398_lb_0_io_rPort_14_banks_1 = x772_x462_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@46568.4]
  assign x398_lb_0_io_rPort_14_banks_0 = x775_x715_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46567.4]
  assign x398_lb_0_io_rPort_14_ofs_0 = x500_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46569.4]
  assign x398_lb_0_io_rPort_14_en_0 = _T_1119 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46571.4]
  assign x398_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46570.4]
  assign x398_lb_0_io_rPort_13_banks_1 = x761_x411_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45783.4]
  assign x398_lb_0_io_rPort_13_banks_0 = x750_x710_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@45782.4]
  assign x398_lb_0_io_rPort_13_ofs_0 = x762_x413_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@45784.4]
  assign x398_lb_0_io_rPort_13_en_0 = _T_658 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@45786.4]
  assign x398_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45785.4]
  assign x398_lb_0_io_rPort_12_banks_1 = x769_x453_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@46952.4]
  assign x398_lb_0_io_rPort_12_banks_0 = x790_x720_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46951.4]
  assign x398_lb_0_io_rPort_12_ofs_0 = x531_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46953.4]
  assign x398_lb_0_io_rPort_12_en_0 = _T_1360 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46955.4]
  assign x398_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46954.4]
  assign x398_lb_0_io_rPort_11_banks_1 = x757_x417_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45703.4]
  assign x398_lb_0_io_rPort_11_banks_0 = x750_x710_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@45702.4]
  assign x398_lb_0_io_rPort_11_ofs_0 = x759_x419_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@45704.4]
  assign x398_lb_0_io_rPort_11_en_0 = _T_613 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@45706.4]
  assign x398_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45705.4]
  assign x398_lb_0_io_rPort_10_banks_1 = x752_x423_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45623.4]
  assign x398_lb_0_io_rPort_10_banks_0 = x750_x710_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@45622.4]
  assign x398_lb_0_io_rPort_10_ofs_0 = x751_x425_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@45624.4]
  assign x398_lb_0_io_rPort_10_en_0 = _T_568 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@45626.4]
  assign x398_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45625.4]
  assign x398_lb_0_io_rPort_9_banks_1 = x766_x403_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@45863.4]
  assign x398_lb_0_io_rPort_9_banks_0 = x750_x710_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@45862.4]
  assign x398_lb_0_io_rPort_9_ofs_0 = x765_x407_sum_D27_number[8:0]; // @[MemInterfaceType.scala 107:54:@45864.4]
  assign x398_lb_0_io_rPort_9_en_0 = _T_703 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@45866.4]
  assign x398_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45865.4]
  assign x398_lb_0_io_rPort_8_banks_1 = x757_x417_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@46785.4]
  assign x398_lb_0_io_rPort_8_banks_0 = x790_x720_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46784.4]
  assign x398_lb_0_io_rPort_8_ofs_0 = x516_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46786.4]
  assign x398_lb_0_io_rPort_8_en_0 = _T_1265 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46788.4]
  assign x398_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46787.4]
  assign x398_lb_0_io_rPort_7_banks_1 = x772_x462_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@46090.4]
  assign x398_lb_0_io_rPort_7_banks_0 = x750_x710_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@46089.4]
  assign x398_lb_0_io_rPort_7_ofs_0 = x464_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46091.4]
  assign x398_lb_0_io_rPort_7_en_0 = _T_834 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46093.4]
  assign x398_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46092.4]
  assign x398_lb_0_io_rPort_6_banks_1 = x752_x423_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@46267.4]
  assign x398_lb_0_io_rPort_6_banks_0 = x775_x715_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46266.4]
  assign x398_lb_0_io_rPort_6_ofs_0 = x475_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46268.4]
  assign x398_lb_0_io_rPort_6_en_0 = _T_954 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46270.4]
  assign x398_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46269.4]
  assign x398_lb_0_io_rPort_5_banks_1 = x772_x462_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@47001.4]
  assign x398_lb_0_io_rPort_5_banks_0 = x790_x720_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@47000.4]
  assign x398_lb_0_io_rPort_5_ofs_0 = x536_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@47002.4]
  assign x398_lb_0_io_rPort_5_en_0 = _T_1389 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@47004.4]
  assign x398_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47003.4]
  assign x398_lb_0_io_rPort_4_banks_1 = x769_x453_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@45982.4]
  assign x398_lb_0_io_rPort_4_banks_0 = x750_x710_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@45981.4]
  assign x398_lb_0_io_rPort_4_ofs_0 = x455_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45983.4]
  assign x398_lb_0_io_rPort_4_en_0 = _T_771 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@45985.4]
  assign x398_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45984.4]
  assign x398_lb_0_io_rPort_3_banks_1 = x761_x411_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@46834.4]
  assign x398_lb_0_io_rPort_3_banks_0 = x790_x720_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46833.4]
  assign x398_lb_0_io_rPort_3_ofs_0 = x521_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46835.4]
  assign x398_lb_0_io_rPort_3_en_0 = _T_1294 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46837.4]
  assign x398_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46836.4]
  assign x398_lb_0_io_rPort_2_banks_1 = x752_x423_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@46736.4]
  assign x398_lb_0_io_rPort_2_banks_0 = x790_x720_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46735.4]
  assign x398_lb_0_io_rPort_2_ofs_0 = x511_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46737.4]
  assign x398_lb_0_io_rPort_2_en_0 = _T_1236 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46739.4]
  assign x398_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46738.4]
  assign x398_lb_0_io_rPort_1_banks_1 = x766_x403_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@46903.4]
  assign x398_lb_0_io_rPort_1_banks_0 = x790_x720_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46902.4]
  assign x398_lb_0_io_rPort_1_ofs_0 = x794_x526_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@46904.4]
  assign x398_lb_0_io_rPort_1_en_0 = _T_1331 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46906.4]
  assign x398_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46905.4]
  assign x398_lb_0_io_rPort_0_banks_1 = x757_x417_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@46325.4]
  assign x398_lb_0_io_rPort_0_banks_0 = x775_x715_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@46324.4]
  assign x398_lb_0_io_rPort_0_ofs_0 = x480_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@46326.4]
  assign x398_lb_0_io_rPort_0_en_0 = _T_986 & x755_b395_D48; // @[MemInterfaceType.scala 110:79:@46328.4]
  assign x398_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46327.4]
  assign x398_lb_0_io_wPort_3_banks_1 = x745_x423_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@45484.4]
  assign x398_lb_0_io_wPort_3_banks_0 = x732_x710_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@45483.4]
  assign x398_lb_0_io_wPort_3_ofs_0 = x744_x425_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@45485.4]
  assign x398_lb_0_io_wPort_3_data_0 = RetimeWrapper_20_io_out; // @[MemInterfaceType.scala 90:56:@45486.4]
  assign x398_lb_0_io_wPort_3_en_0 = _T_497 & x736_b395_D24; // @[MemInterfaceType.scala 93:57:@45488.4]
  assign x398_lb_0_io_wPort_2_banks_1 = x741_x417_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@45386.4]
  assign x398_lb_0_io_wPort_2_banks_0 = x732_x710_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@45385.4]
  assign x398_lb_0_io_wPort_2_ofs_0 = x743_x419_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@45387.4]
  assign x398_lb_0_io_wPort_2_data_0 = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 90:56:@45388.4]
  assign x398_lb_0_io_wPort_2_en_0 = _T_449 & x736_b395_D24; // @[MemInterfaceType.scala 93:57:@45390.4]
  assign x398_lb_0_io_wPort_1_banks_1 = x738_x411_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@45288.4]
  assign x398_lb_0_io_wPort_1_banks_0 = x732_x710_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@45287.4]
  assign x398_lb_0_io_wPort_1_ofs_0 = x739_x413_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@45289.4]
  assign x398_lb_0_io_wPort_1_data_0 = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 90:56:@45290.4]
  assign x398_lb_0_io_wPort_1_en_0 = _T_401 & x736_b395_D24; // @[MemInterfaceType.scala 93:57:@45292.4]
  assign x398_lb_0_io_wPort_0_banks_1 = x733_x403_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@45181.4]
  assign x398_lb_0_io_wPort_0_banks_0 = x732_x710_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@45180.4]
  assign x398_lb_0_io_wPort_0_ofs_0 = x731_x407_sum_D3_number[8:0]; // @[MemInterfaceType.scala 89:54:@45182.4]
  assign x398_lb_0_io_wPort_0_data_0 = RetimeWrapper_6_io_out; // @[MemInterfaceType.scala 90:56:@45183.4]
  assign x398_lb_0_io_wPort_0_en_0 = _T_350 & x736_b395_D24; // @[MemInterfaceType.scala 93:57:@45185.4]
  assign x403_1_clock = clock; // @[:@45033.4]
  assign x403_1_io_a = __1_io_result; // @[Math.scala 367:17:@45035.4]
  assign x403_1_io_flow = io_in_x354_TREADY; // @[Math.scala 369:20:@45037.4]
  assign x713_sum_1_clock = clock; // @[:@45070.4]
  assign x713_sum_1_reset = reset; // @[:@45071.4]
  assign x713_sum_1_io_a = _T_300[31:0]; // @[Math.scala 151:17:@45072.4]
  assign x713_sum_1_io_b = _T_303[31:0]; // @[Math.scala 152:17:@45073.4]
  assign x713_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45074.4]
  assign x406_div_1_clock = clock; // @[:@45082.4]
  assign x406_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@45084.4]
  assign x406_div_1_io_flow = io_in_x354_TREADY; // @[Math.scala 330:20:@45086.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45092.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45093.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45095.4]
  assign RetimeWrapper_1_io_in = x713_sum_1_io_result; // @[package.scala 94:16:@45094.4]
  assign x407_sum_1_clock = clock; // @[:@45101.4]
  assign x407_sum_1_reset = reset; // @[:@45102.4]
  assign x407_sum_1_io_a = RetimeWrapper_1_io_out; // @[Math.scala 151:17:@45103.4]
  assign x407_sum_1_io_b = x406_div_1_io_result; // @[Math.scala 152:17:@45104.4]
  assign x407_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45105.4]
  assign RetimeWrapper_2_clock = clock; // @[:@45111.4]
  assign RetimeWrapper_2_reset = reset; // @[:@45112.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45114.4]
  assign RetimeWrapper_2_io_in = x407_sum_1_io_result; // @[package.scala 94:16:@45113.4]
  assign RetimeWrapper_3_clock = clock; // @[:@45120.4]
  assign RetimeWrapper_3_reset = reset; // @[:@45121.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45123.4]
  assign RetimeWrapper_3_io_in = $unsigned(_T_263); // @[package.scala 94:16:@45122.4]
  assign RetimeWrapper_4_clock = clock; // @[:@45129.4]
  assign RetimeWrapper_4_reset = reset; // @[:@45130.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45132.4]
  assign RetimeWrapper_4_io_in = x403_1_io_result; // @[package.scala 94:16:@45131.4]
  assign RetimeWrapper_5_clock = clock; // @[:@45138.4]
  assign RetimeWrapper_5_reset = reset; // @[:@45139.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45141.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@45140.4]
  assign RetimeWrapper_6_clock = clock; // @[:@45147.4]
  assign RetimeWrapper_6_reset = reset; // @[:@45148.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45150.4]
  assign RetimeWrapper_6_io_in = x729_x396_D1_0_number[31:0]; // @[package.scala 94:16:@45149.4]
  assign RetimeWrapper_7_clock = clock; // @[:@45156.4]
  assign RetimeWrapper_7_reset = reset; // @[:@45157.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45159.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@45158.4]
  assign RetimeWrapper_8_clock = clock; // @[:@45167.4]
  assign RetimeWrapper_8_reset = reset; // @[:@45168.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45170.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45169.4]
  assign x409_rdcol_1_clock = clock; // @[:@45190.4]
  assign x409_rdcol_1_reset = reset; // @[:@45191.4]
  assign x409_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@45192.4]
  assign x409_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@45193.4]
  assign x409_rdcol_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45194.4]
  assign x411_1_clock = clock; // @[:@45204.4]
  assign x411_1_io_a = x409_rdcol_1_io_result; // @[Math.scala 367:17:@45206.4]
  assign x411_1_io_flow = io_in_x354_TREADY; // @[Math.scala 369:20:@45208.4]
  assign x412_div_1_clock = clock; // @[:@45216.4]
  assign x412_div_1_io_a = x409_rdcol_1_io_result; // @[Math.scala 328:17:@45218.4]
  assign x412_div_1_io_flow = io_in_x354_TREADY; // @[Math.scala 330:20:@45220.4]
  assign RetimeWrapper_9_clock = clock; // @[:@45226.4]
  assign RetimeWrapper_9_reset = reset; // @[:@45227.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45229.4]
  assign RetimeWrapper_9_io_in = x713_sum_1_io_result; // @[package.scala 94:16:@45228.4]
  assign x413_sum_1_clock = clock; // @[:@45235.4]
  assign x413_sum_1_reset = reset; // @[:@45236.4]
  assign x413_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@45237.4]
  assign x413_sum_1_io_b = x412_div_1_io_result; // @[Math.scala 152:17:@45238.4]
  assign x413_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45239.4]
  assign RetimeWrapper_10_clock = clock; // @[:@45245.4]
  assign RetimeWrapper_10_reset = reset; // @[:@45246.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45248.4]
  assign RetimeWrapper_10_io_in = x411_1_io_result; // @[package.scala 94:16:@45247.4]
  assign RetimeWrapper_11_clock = clock; // @[:@45254.4]
  assign RetimeWrapper_11_reset = reset; // @[:@45255.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45257.4]
  assign RetimeWrapper_11_io_in = x413_sum_1_io_result; // @[package.scala 94:16:@45256.4]
  assign RetimeWrapper_12_clock = clock; // @[:@45263.4]
  assign RetimeWrapper_12_reset = reset; // @[:@45264.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45266.4]
  assign RetimeWrapper_12_io_in = x729_x396_D1_0_number[63:32]; // @[package.scala 94:16:@45265.4]
  assign RetimeWrapper_13_clock = clock; // @[:@45274.4]
  assign RetimeWrapper_13_reset = reset; // @[:@45275.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45277.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45276.4]
  assign x415_rdcol_1_clock = clock; // @[:@45297.4]
  assign x415_rdcol_1_reset = reset; // @[:@45298.4]
  assign x415_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@45299.4]
  assign x415_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@45300.4]
  assign x415_rdcol_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45301.4]
  assign x417_1_clock = clock; // @[:@45311.4]
  assign x417_1_io_a = x415_rdcol_1_io_result; // @[Math.scala 367:17:@45313.4]
  assign x417_1_io_flow = io_in_x354_TREADY; // @[Math.scala 369:20:@45315.4]
  assign x418_div_1_clock = clock; // @[:@45323.4]
  assign x418_div_1_io_a = x415_rdcol_1_io_result; // @[Math.scala 328:17:@45325.4]
  assign x418_div_1_io_flow = io_in_x354_TREADY; // @[Math.scala 330:20:@45327.4]
  assign x419_sum_1_clock = clock; // @[:@45333.4]
  assign x419_sum_1_reset = reset; // @[:@45334.4]
  assign x419_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@45335.4]
  assign x419_sum_1_io_b = x418_div_1_io_result; // @[Math.scala 152:17:@45336.4]
  assign x419_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45337.4]
  assign RetimeWrapper_14_clock = clock; // @[:@45343.4]
  assign RetimeWrapper_14_reset = reset; // @[:@45344.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45346.4]
  assign RetimeWrapper_14_io_in = x417_1_io_result; // @[package.scala 94:16:@45345.4]
  assign RetimeWrapper_15_clock = clock; // @[:@45352.4]
  assign RetimeWrapper_15_reset = reset; // @[:@45353.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45355.4]
  assign RetimeWrapper_15_io_in = x729_x396_D1_0_number[95:64]; // @[package.scala 94:16:@45354.4]
  assign RetimeWrapper_16_clock = clock; // @[:@45361.4]
  assign RetimeWrapper_16_reset = reset; // @[:@45362.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45364.4]
  assign RetimeWrapper_16_io_in = x419_sum_1_io_result; // @[package.scala 94:16:@45363.4]
  assign RetimeWrapper_17_clock = clock; // @[:@45372.4]
  assign RetimeWrapper_17_reset = reset; // @[:@45373.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45375.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45374.4]
  assign x421_rdcol_1_clock = clock; // @[:@45395.4]
  assign x421_rdcol_1_reset = reset; // @[:@45396.4]
  assign x421_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@45397.4]
  assign x421_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@45398.4]
  assign x421_rdcol_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45399.4]
  assign x423_1_clock = clock; // @[:@45409.4]
  assign x423_1_io_a = x421_rdcol_1_io_result; // @[Math.scala 367:17:@45411.4]
  assign x423_1_io_flow = io_in_x354_TREADY; // @[Math.scala 369:20:@45413.4]
  assign x424_div_1_clock = clock; // @[:@45421.4]
  assign x424_div_1_io_a = x421_rdcol_1_io_result; // @[Math.scala 328:17:@45423.4]
  assign x424_div_1_io_flow = io_in_x354_TREADY; // @[Math.scala 330:20:@45425.4]
  assign x425_sum_1_clock = clock; // @[:@45431.4]
  assign x425_sum_1_reset = reset; // @[:@45432.4]
  assign x425_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@45433.4]
  assign x425_sum_1_io_b = x424_div_1_io_result; // @[Math.scala 152:17:@45434.4]
  assign x425_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45435.4]
  assign RetimeWrapper_18_clock = clock; // @[:@45441.4]
  assign RetimeWrapper_18_reset = reset; // @[:@45442.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45444.4]
  assign RetimeWrapper_18_io_in = x425_sum_1_io_result; // @[package.scala 94:16:@45443.4]
  assign RetimeWrapper_19_clock = clock; // @[:@45450.4]
  assign RetimeWrapper_19_reset = reset; // @[:@45451.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45453.4]
  assign RetimeWrapper_19_io_in = x423_1_io_result; // @[package.scala 94:16:@45452.4]
  assign RetimeWrapper_20_clock = clock; // @[:@45459.4]
  assign RetimeWrapper_20_reset = reset; // @[:@45460.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45462.4]
  assign RetimeWrapper_20_io_in = x729_x396_D1_0_number[127:96]; // @[package.scala 94:16:@45461.4]
  assign RetimeWrapper_21_clock = clock; // @[:@45470.4]
  assign RetimeWrapper_21_reset = reset; // @[:@45471.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45473.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45472.4]
  assign RetimeWrapper_22_clock = clock; // @[:@45491.4]
  assign RetimeWrapper_22_reset = reset; // @[:@45492.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45494.4]
  assign RetimeWrapper_22_io_in = __io_result; // @[package.scala 94:16:@45493.4]
  assign RetimeWrapper_23_clock = clock; // @[:@45507.4]
  assign RetimeWrapper_23_reset = reset; // @[:@45508.4]
  assign RetimeWrapper_23_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@45510.4]
  assign RetimeWrapper_23_io_in = $signed(_T_509) < $signed(32'sh0); // @[package.scala 94:16:@45509.4]
  assign RetimeWrapper_24_clock = clock; // @[:@45516.4]
  assign RetimeWrapper_24_reset = reset; // @[:@45517.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45519.4]
  assign RetimeWrapper_24_io_in = x421_rdcol_1_io_result; // @[package.scala 94:16:@45518.4]
  assign RetimeWrapper_25_clock = clock; // @[:@45530.4]
  assign RetimeWrapper_25_reset = reset; // @[:@45531.4]
  assign RetimeWrapper_25_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@45533.4]
  assign RetimeWrapper_25_io_in = $signed(_T_522) < $signed(32'sh0); // @[package.scala 94:16:@45532.4]
  assign RetimeWrapper_26_clock = clock; // @[:@45539.4]
  assign RetimeWrapper_26_reset = reset; // @[:@45540.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45542.4]
  assign RetimeWrapper_26_io_in = RetimeWrapper_23_io_out; // @[package.scala 94:16:@45541.4]
  assign RetimeWrapper_27_clock = clock; // @[:@45554.4]
  assign RetimeWrapper_27_reset = reset; // @[:@45555.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45557.4]
  assign RetimeWrapper_27_io_in = $unsigned(_T_263); // @[package.scala 94:16:@45556.4]
  assign RetimeWrapper_28_clock = clock; // @[:@45563.4]
  assign RetimeWrapper_28_reset = reset; // @[:@45564.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45566.4]
  assign RetimeWrapper_28_io_in = x425_sum_1_io_result; // @[package.scala 94:16:@45565.4]
  assign RetimeWrapper_29_clock = clock; // @[:@45572.4]
  assign RetimeWrapper_29_reset = reset; // @[:@45573.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45575.4]
  assign RetimeWrapper_29_io_in = x423_1_io_result; // @[package.scala 94:16:@45574.4]
  assign RetimeWrapper_30_clock = clock; // @[:@45581.4]
  assign RetimeWrapper_30_reset = reset; // @[:@45582.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45584.4]
  assign RetimeWrapper_30_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@45583.4]
  assign RetimeWrapper_31_clock = clock; // @[:@45590.4]
  assign RetimeWrapper_31_reset = reset; // @[:@45591.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45593.4]
  assign RetimeWrapper_31_io_in = ~ x430; // @[package.scala 94:16:@45592.4]
  assign RetimeWrapper_32_clock = clock; // @[:@45599.4]
  assign RetimeWrapper_32_reset = reset; // @[:@45600.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45602.4]
  assign RetimeWrapper_32_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@45601.4]
  assign RetimeWrapper_33_clock = clock; // @[:@45611.4]
  assign RetimeWrapper_33_reset = reset; // @[:@45612.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45614.4]
  assign RetimeWrapper_33_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45613.4]
  assign RetimeWrapper_34_clock = clock; // @[:@45632.4]
  assign RetimeWrapper_34_reset = reset; // @[:@45633.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45635.4]
  assign RetimeWrapper_34_io_in = x415_rdcol_1_io_result; // @[package.scala 94:16:@45634.4]
  assign RetimeWrapper_35_clock = clock; // @[:@45646.4]
  assign RetimeWrapper_35_reset = reset; // @[:@45647.4]
  assign RetimeWrapper_35_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@45649.4]
  assign RetimeWrapper_35_io_in = $signed(_T_579) < $signed(32'sh0); // @[package.scala 94:16:@45648.4]
  assign RetimeWrapper_36_clock = clock; // @[:@45661.4]
  assign RetimeWrapper_36_reset = reset; // @[:@45662.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45664.4]
  assign RetimeWrapper_36_io_in = x417_1_io_result; // @[package.scala 94:16:@45663.4]
  assign RetimeWrapper_37_clock = clock; // @[:@45670.4]
  assign RetimeWrapper_37_reset = reset; // @[:@45671.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45673.4]
  assign RetimeWrapper_37_io_in = ~ x435; // @[package.scala 94:16:@45672.4]
  assign RetimeWrapper_38_clock = clock; // @[:@45679.4]
  assign RetimeWrapper_38_reset = reset; // @[:@45680.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45682.4]
  assign RetimeWrapper_38_io_in = x419_sum_1_io_result; // @[package.scala 94:16:@45681.4]
  assign RetimeWrapper_39_clock = clock; // @[:@45691.4]
  assign RetimeWrapper_39_reset = reset; // @[:@45692.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45694.4]
  assign RetimeWrapper_39_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45693.4]
  assign RetimeWrapper_40_clock = clock; // @[:@45712.4]
  assign RetimeWrapper_40_reset = reset; // @[:@45713.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45715.4]
  assign RetimeWrapper_40_io_in = x409_rdcol_1_io_result; // @[package.scala 94:16:@45714.4]
  assign RetimeWrapper_41_clock = clock; // @[:@45726.4]
  assign RetimeWrapper_41_reset = reset; // @[:@45727.4]
  assign RetimeWrapper_41_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@45729.4]
  assign RetimeWrapper_41_io_in = $signed(_T_624) < $signed(32'sh0); // @[package.scala 94:16:@45728.4]
  assign RetimeWrapper_42_clock = clock; // @[:@45741.4]
  assign RetimeWrapper_42_reset = reset; // @[:@45742.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45744.4]
  assign RetimeWrapper_42_io_in = x411_1_io_result; // @[package.scala 94:16:@45743.4]
  assign RetimeWrapper_43_clock = clock; // @[:@45750.4]
  assign RetimeWrapper_43_reset = reset; // @[:@45751.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45753.4]
  assign RetimeWrapper_43_io_in = x413_sum_1_io_result; // @[package.scala 94:16:@45752.4]
  assign RetimeWrapper_44_clock = clock; // @[:@45759.4]
  assign RetimeWrapper_44_reset = reset; // @[:@45760.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45762.4]
  assign RetimeWrapper_44_io_in = ~ x440; // @[package.scala 94:16:@45761.4]
  assign RetimeWrapper_45_clock = clock; // @[:@45771.4]
  assign RetimeWrapper_45_reset = reset; // @[:@45772.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45774.4]
  assign RetimeWrapper_45_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45773.4]
  assign RetimeWrapper_46_clock = clock; // @[:@45792.4]
  assign RetimeWrapper_46_reset = reset; // @[:@45793.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45795.4]
  assign RetimeWrapper_46_io_in = __1_io_result; // @[package.scala 94:16:@45794.4]
  assign RetimeWrapper_47_clock = clock; // @[:@45806.4]
  assign RetimeWrapper_47_reset = reset; // @[:@45807.4]
  assign RetimeWrapper_47_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@45809.4]
  assign RetimeWrapper_47_io_in = $signed(_T_669) < $signed(32'sh0); // @[package.scala 94:16:@45808.4]
  assign RetimeWrapper_48_clock = clock; // @[:@45821.4]
  assign RetimeWrapper_48_reset = reset; // @[:@45822.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45824.4]
  assign RetimeWrapper_48_io_in = x407_sum_1_io_result; // @[package.scala 94:16:@45823.4]
  assign RetimeWrapper_49_clock = clock; // @[:@45830.4]
  assign RetimeWrapper_49_reset = reset; // @[:@45831.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45833.4]
  assign RetimeWrapper_49_io_in = x403_1_io_result; // @[package.scala 94:16:@45832.4]
  assign RetimeWrapper_50_clock = clock; // @[:@45839.4]
  assign RetimeWrapper_50_reset = reset; // @[:@45840.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45842.4]
  assign RetimeWrapper_50_io_in = ~ x445; // @[package.scala 94:16:@45841.4]
  assign RetimeWrapper_51_clock = clock; // @[:@45851.4]
  assign RetimeWrapper_51_reset = reset; // @[:@45852.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45854.4]
  assign RetimeWrapper_51_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45853.4]
  assign x449_rdcol_1_clock = clock; // @[:@45874.4]
  assign x449_rdcol_1_reset = reset; // @[:@45875.4]
  assign x449_rdcol_1_io_a = RetimeWrapper_46_io_out; // @[Math.scala 151:17:@45876.4]
  assign x449_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@45877.4]
  assign x449_rdcol_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45878.4]
  assign RetimeWrapper_52_clock = clock; // @[:@45889.4]
  assign RetimeWrapper_52_reset = reset; // @[:@45890.4]
  assign RetimeWrapper_52_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@45892.4]
  assign RetimeWrapper_52_io_in = $signed(_T_718) < $signed(32'sh0); // @[package.scala 94:16:@45891.4]
  assign x453_1_clock = clock; // @[:@45908.4]
  assign x453_1_io_a = x449_rdcol_1_io_result; // @[Math.scala 367:17:@45910.4]
  assign x453_1_io_flow = io_in_x354_TREADY; // @[Math.scala 369:20:@45912.4]
  assign x454_div_1_clock = clock; // @[:@45920.4]
  assign x454_div_1_io_a = x449_rdcol_1_io_result; // @[Math.scala 328:17:@45922.4]
  assign x454_div_1_io_flow = io_in_x354_TREADY; // @[Math.scala 330:20:@45924.4]
  assign RetimeWrapper_53_clock = clock; // @[:@45930.4]
  assign RetimeWrapper_53_reset = reset; // @[:@45931.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45933.4]
  assign RetimeWrapper_53_io_in = x713_sum_1_io_result; // @[package.scala 94:16:@45932.4]
  assign x455_sum_1_clock = clock; // @[:@45939.4]
  assign x455_sum_1_reset = reset; // @[:@45940.4]
  assign x455_sum_1_io_a = RetimeWrapper_53_io_out; // @[Math.scala 151:17:@45941.4]
  assign x455_sum_1_io_b = x454_div_1_io_result; // @[Math.scala 152:17:@45942.4]
  assign x455_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45943.4]
  assign RetimeWrapper_54_clock = clock; // @[:@45949.4]
  assign RetimeWrapper_54_reset = reset; // @[:@45950.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45952.4]
  assign RetimeWrapper_54_io_in = x453_1_io_result; // @[package.scala 94:16:@45951.4]
  assign RetimeWrapper_55_clock = clock; // @[:@45958.4]
  assign RetimeWrapper_55_reset = reset; // @[:@45959.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45961.4]
  assign RetimeWrapper_55_io_in = ~ x451; // @[package.scala 94:16:@45960.4]
  assign RetimeWrapper_56_clock = clock; // @[:@45970.4]
  assign RetimeWrapper_56_reset = reset; // @[:@45971.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45973.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45972.4]
  assign x458_rdcol_1_clock = clock; // @[:@45993.4]
  assign x458_rdcol_1_reset = reset; // @[:@45994.4]
  assign x458_rdcol_1_io_a = RetimeWrapper_46_io_out; // @[Math.scala 151:17:@45995.4]
  assign x458_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@45996.4]
  assign x458_rdcol_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@45997.4]
  assign RetimeWrapper_57_clock = clock; // @[:@46008.4]
  assign RetimeWrapper_57_reset = reset; // @[:@46009.4]
  assign RetimeWrapper_57_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@46011.4]
  assign RetimeWrapper_57_io_in = $signed(_T_786) < $signed(32'sh0); // @[package.scala 94:16:@46010.4]
  assign x462_1_clock = clock; // @[:@46025.4]
  assign x462_1_io_a = x458_rdcol_1_io_result; // @[Math.scala 367:17:@46027.4]
  assign x462_1_io_flow = io_in_x354_TREADY; // @[Math.scala 369:20:@46029.4]
  assign x463_div_1_clock = clock; // @[:@46037.4]
  assign x463_div_1_io_a = x458_rdcol_1_io_result; // @[Math.scala 328:17:@46039.4]
  assign x463_div_1_io_flow = io_in_x354_TREADY; // @[Math.scala 330:20:@46041.4]
  assign x464_sum_1_clock = clock; // @[:@46047.4]
  assign x464_sum_1_reset = reset; // @[:@46048.4]
  assign x464_sum_1_io_a = RetimeWrapper_53_io_out; // @[Math.scala 151:17:@46049.4]
  assign x464_sum_1_io_b = x463_div_1_io_result; // @[Math.scala 152:17:@46050.4]
  assign x464_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46051.4]
  assign RetimeWrapper_58_clock = clock; // @[:@46057.4]
  assign RetimeWrapper_58_reset = reset; // @[:@46058.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46060.4]
  assign RetimeWrapper_58_io_in = ~ x460; // @[package.scala 94:16:@46059.4]
  assign RetimeWrapper_59_clock = clock; // @[:@46066.4]
  assign RetimeWrapper_59_reset = reset; // @[:@46067.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46069.4]
  assign RetimeWrapper_59_io_in = x462_1_io_result; // @[package.scala 94:16:@46068.4]
  assign RetimeWrapper_60_clock = clock; // @[:@46078.4]
  assign RetimeWrapper_60_reset = reset; // @[:@46079.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46081.4]
  assign RetimeWrapper_60_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46080.4]
  assign x467_rdrow_1_clock = clock; // @[:@46101.4]
  assign x467_rdrow_1_reset = reset; // @[:@46102.4]
  assign x467_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@46103.4]
  assign x467_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@46104.4]
  assign x467_rdrow_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@46105.4]
  assign RetimeWrapper_61_clock = clock; // @[:@46127.4]
  assign RetimeWrapper_61_reset = reset; // @[:@46128.4]
  assign RetimeWrapper_61_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@46130.4]
  assign RetimeWrapper_61_io_in = $signed(_T_851) < $signed(32'sh0); // @[package.scala 94:16:@46129.4]
  assign RetimeWrapper_62_clock = clock; // @[:@46149.4]
  assign RetimeWrapper_62_reset = reset; // @[:@46150.4]
  assign RetimeWrapper_62_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@46153.4]
  assign RetimeWrapper_62_io_in = $unsigned(_T_880); // @[package.scala 94:16:@46152.4]
  assign RetimeWrapper_63_clock = clock; // @[:@46175.4]
  assign RetimeWrapper_63_reset = reset; // @[:@46176.4]
  assign RetimeWrapper_63_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@46178.4]
  assign RetimeWrapper_63_io_in = {_T_892,_T_893}; // @[package.scala 94:16:@46177.4]
  assign x718_sum_1_clock = clock; // @[:@46196.4]
  assign x718_sum_1_reset = reset; // @[:@46197.4]
  assign x718_sum_1_io_a = _T_916[31:0]; // @[Math.scala 151:17:@46198.4]
  assign x718_sum_1_io_b = _T_919[31:0]; // @[Math.scala 152:17:@46199.4]
  assign x718_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46200.4]
  assign RetimeWrapper_64_clock = clock; // @[:@46206.4]
  assign RetimeWrapper_64_reset = reset; // @[:@46207.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46209.4]
  assign RetimeWrapper_64_io_in = x718_sum_1_io_result; // @[package.scala 94:16:@46208.4]
  assign RetimeWrapper_65_clock = clock; // @[:@46215.4]
  assign RetimeWrapper_65_reset = reset; // @[:@46216.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46218.4]
  assign RetimeWrapper_65_io_in = x424_div_1_io_result; // @[package.scala 94:16:@46217.4]
  assign x475_sum_1_clock = clock; // @[:@46224.4]
  assign x475_sum_1_reset = reset; // @[:@46225.4]
  assign x475_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@46226.4]
  assign x475_sum_1_io_b = RetimeWrapper_65_io_out; // @[Math.scala 152:17:@46227.4]
  assign x475_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46228.4]
  assign RetimeWrapper_66_clock = clock; // @[:@46234.4]
  assign RetimeWrapper_66_reset = reset; // @[:@46235.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46237.4]
  assign RetimeWrapper_66_io_in = $unsigned(_T_884); // @[package.scala 94:16:@46236.4]
  assign RetimeWrapper_67_clock = clock; // @[:@46243.4]
  assign RetimeWrapper_67_reset = reset; // @[:@46244.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46246.4]
  assign RetimeWrapper_67_io_in = ~ x470; // @[package.scala 94:16:@46245.4]
  assign RetimeWrapper_68_clock = clock; // @[:@46255.4]
  assign RetimeWrapper_68_reset = reset; // @[:@46256.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46258.4]
  assign RetimeWrapper_68_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46257.4]
  assign RetimeWrapper_69_clock = clock; // @[:@46282.4]
  assign RetimeWrapper_69_reset = reset; // @[:@46283.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46285.4]
  assign RetimeWrapper_69_io_in = x418_div_1_io_result; // @[package.scala 94:16:@46284.4]
  assign x480_sum_1_clock = clock; // @[:@46291.4]
  assign x480_sum_1_reset = reset; // @[:@46292.4]
  assign x480_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@46293.4]
  assign x480_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@46294.4]
  assign x480_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46295.4]
  assign RetimeWrapper_70_clock = clock; // @[:@46301.4]
  assign RetimeWrapper_70_reset = reset; // @[:@46302.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46304.4]
  assign RetimeWrapper_70_io_in = ~ x478; // @[package.scala 94:16:@46303.4]
  assign RetimeWrapper_71_clock = clock; // @[:@46313.4]
  assign RetimeWrapper_71_reset = reset; // @[:@46314.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46316.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46315.4]
  assign RetimeWrapper_72_clock = clock; // @[:@46340.4]
  assign RetimeWrapper_72_reset = reset; // @[:@46341.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46343.4]
  assign RetimeWrapper_72_io_in = x412_div_1_io_result; // @[package.scala 94:16:@46342.4]
  assign x485_sum_1_clock = clock; // @[:@46349.4]
  assign x485_sum_1_reset = reset; // @[:@46350.4]
  assign x485_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@46351.4]
  assign x485_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@46352.4]
  assign x485_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46353.4]
  assign RetimeWrapper_73_clock = clock; // @[:@46359.4]
  assign RetimeWrapper_73_reset = reset; // @[:@46360.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46362.4]
  assign RetimeWrapper_73_io_in = ~ x483; // @[package.scala 94:16:@46361.4]
  assign RetimeWrapper_74_clock = clock; // @[:@46371.4]
  assign RetimeWrapper_74_reset = reset; // @[:@46372.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46374.4]
  assign RetimeWrapper_74_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46373.4]
  assign RetimeWrapper_75_clock = clock; // @[:@46392.4]
  assign RetimeWrapper_75_reset = reset; // @[:@46393.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46395.4]
  assign RetimeWrapper_75_io_in = RetimeWrapper_47_io_out; // @[package.scala 94:16:@46394.4]
  assign RetimeWrapper_76_clock = clock; // @[:@46407.4]
  assign RetimeWrapper_76_reset = reset; // @[:@46408.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46410.4]
  assign RetimeWrapper_76_io_in = x406_div_1_io_result; // @[package.scala 94:16:@46409.4]
  assign RetimeWrapper_77_clock = clock; // @[:@46416.4]
  assign RetimeWrapper_77_reset = reset; // @[:@46417.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46419.4]
  assign RetimeWrapper_77_io_in = x718_sum_1_io_result; // @[package.scala 94:16:@46418.4]
  assign x490_sum_1_clock = clock; // @[:@46427.4]
  assign x490_sum_1_reset = reset; // @[:@46428.4]
  assign x490_sum_1_io_a = RetimeWrapper_77_io_out; // @[Math.scala 151:17:@46429.4]
  assign x490_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@46430.4]
  assign x490_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46431.4]
  assign RetimeWrapper_78_clock = clock; // @[:@46437.4]
  assign RetimeWrapper_78_reset = reset; // @[:@46438.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46440.4]
  assign RetimeWrapper_78_io_in = ~ x488; // @[package.scala 94:16:@46439.4]
  assign RetimeWrapper_79_clock = clock; // @[:@46446.4]
  assign RetimeWrapper_79_reset = reset; // @[:@46447.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46449.4]
  assign RetimeWrapper_79_io_in = x490_sum_1_io_result; // @[package.scala 94:16:@46448.4]
  assign RetimeWrapper_80_clock = clock; // @[:@46458.4]
  assign RetimeWrapper_80_reset = reset; // @[:@46459.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46461.4]
  assign RetimeWrapper_80_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46460.4]
  assign x495_sum_1_clock = clock; // @[:@46485.4]
  assign x495_sum_1_reset = reset; // @[:@46486.4]
  assign x495_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@46487.4]
  assign x495_sum_1_io_b = x454_div_1_io_result; // @[Math.scala 152:17:@46488.4]
  assign x495_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46489.4]
  assign RetimeWrapper_81_clock = clock; // @[:@46495.4]
  assign RetimeWrapper_81_reset = reset; // @[:@46496.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46498.4]
  assign RetimeWrapper_81_io_in = ~ x493; // @[package.scala 94:16:@46497.4]
  assign RetimeWrapper_82_clock = clock; // @[:@46507.4]
  assign RetimeWrapper_82_reset = reset; // @[:@46508.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46510.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46509.4]
  assign x500_sum_1_clock = clock; // @[:@46534.4]
  assign x500_sum_1_reset = reset; // @[:@46535.4]
  assign x500_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@46536.4]
  assign x500_sum_1_io_b = x463_div_1_io_result; // @[Math.scala 152:17:@46537.4]
  assign x500_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46538.4]
  assign RetimeWrapper_83_clock = clock; // @[:@46544.4]
  assign RetimeWrapper_83_reset = reset; // @[:@46545.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46547.4]
  assign RetimeWrapper_83_io_in = ~ x498; // @[package.scala 94:16:@46546.4]
  assign RetimeWrapper_84_clock = clock; // @[:@46556.4]
  assign RetimeWrapper_84_reset = reset; // @[:@46557.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46559.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46558.4]
  assign x503_rdrow_1_clock = clock; // @[:@46579.4]
  assign x503_rdrow_1_reset = reset; // @[:@46580.4]
  assign x503_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@46581.4]
  assign x503_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@46582.4]
  assign x503_rdrow_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@46583.4]
  assign RetimeWrapper_85_clock = clock; // @[:@46605.4]
  assign RetimeWrapper_85_reset = reset; // @[:@46606.4]
  assign RetimeWrapper_85_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@46608.4]
  assign RetimeWrapper_85_io_in = $signed(_T_1136) < $signed(32'sh0); // @[package.scala 94:16:@46607.4]
  assign RetimeWrapper_86_clock = clock; // @[:@46627.4]
  assign RetimeWrapper_86_reset = reset; // @[:@46628.4]
  assign RetimeWrapper_86_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@46631.4]
  assign RetimeWrapper_86_io_in = $unsigned(_T_1165); // @[package.scala 94:16:@46630.4]
  assign RetimeWrapper_87_clock = clock; // @[:@46653.4]
  assign RetimeWrapper_87_reset = reset; // @[:@46654.4]
  assign RetimeWrapper_87_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@46656.4]
  assign RetimeWrapper_87_io_in = {_T_1177,_T_1178}; // @[package.scala 94:16:@46655.4]
  assign x723_sum_1_clock = clock; // @[:@46674.4]
  assign x723_sum_1_reset = reset; // @[:@46675.4]
  assign x723_sum_1_io_a = _T_1201[31:0]; // @[Math.scala 151:17:@46676.4]
  assign x723_sum_1_io_b = _T_1204[31:0]; // @[Math.scala 152:17:@46677.4]
  assign x723_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46678.4]
  assign RetimeWrapper_88_clock = clock; // @[:@46684.4]
  assign RetimeWrapper_88_reset = reset; // @[:@46685.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46687.4]
  assign RetimeWrapper_88_io_in = x723_sum_1_io_result; // @[package.scala 94:16:@46686.4]
  assign x511_sum_1_clock = clock; // @[:@46693.4]
  assign x511_sum_1_reset = reset; // @[:@46694.4]
  assign x511_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@46695.4]
  assign x511_sum_1_io_b = RetimeWrapper_65_io_out; // @[Math.scala 152:17:@46696.4]
  assign x511_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46697.4]
  assign RetimeWrapper_89_clock = clock; // @[:@46703.4]
  assign RetimeWrapper_89_reset = reset; // @[:@46704.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46706.4]
  assign RetimeWrapper_89_io_in = ~ x506; // @[package.scala 94:16:@46705.4]
  assign RetimeWrapper_90_clock = clock; // @[:@46712.4]
  assign RetimeWrapper_90_reset = reset; // @[:@46713.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46715.4]
  assign RetimeWrapper_90_io_in = $unsigned(_T_1169); // @[package.scala 94:16:@46714.4]
  assign RetimeWrapper_91_clock = clock; // @[:@46724.4]
  assign RetimeWrapper_91_reset = reset; // @[:@46725.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46727.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46726.4]
  assign x516_sum_1_clock = clock; // @[:@46751.4]
  assign x516_sum_1_reset = reset; // @[:@46752.4]
  assign x516_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@46753.4]
  assign x516_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@46754.4]
  assign x516_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46755.4]
  assign RetimeWrapper_92_clock = clock; // @[:@46761.4]
  assign RetimeWrapper_92_reset = reset; // @[:@46762.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46764.4]
  assign RetimeWrapper_92_io_in = ~ x514; // @[package.scala 94:16:@46763.4]
  assign RetimeWrapper_93_clock = clock; // @[:@46773.4]
  assign RetimeWrapper_93_reset = reset; // @[:@46774.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46776.4]
  assign RetimeWrapper_93_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46775.4]
  assign x521_sum_1_clock = clock; // @[:@46800.4]
  assign x521_sum_1_reset = reset; // @[:@46801.4]
  assign x521_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@46802.4]
  assign x521_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@46803.4]
  assign x521_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46804.4]
  assign RetimeWrapper_94_clock = clock; // @[:@46810.4]
  assign RetimeWrapper_94_reset = reset; // @[:@46811.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46813.4]
  assign RetimeWrapper_94_io_in = ~ x519; // @[package.scala 94:16:@46812.4]
  assign RetimeWrapper_95_clock = clock; // @[:@46822.4]
  assign RetimeWrapper_95_reset = reset; // @[:@46823.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46825.4]
  assign RetimeWrapper_95_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46824.4]
  assign RetimeWrapper_96_clock = clock; // @[:@46849.4]
  assign RetimeWrapper_96_reset = reset; // @[:@46850.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46852.4]
  assign RetimeWrapper_96_io_in = x723_sum_1_io_result; // @[package.scala 94:16:@46851.4]
  assign x526_sum_1_clock = clock; // @[:@46860.4]
  assign x526_sum_1_reset = reset; // @[:@46861.4]
  assign x526_sum_1_io_a = RetimeWrapper_96_io_out; // @[Math.scala 151:17:@46862.4]
  assign x526_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@46863.4]
  assign x526_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46864.4]
  assign RetimeWrapper_97_clock = clock; // @[:@46870.4]
  assign RetimeWrapper_97_reset = reset; // @[:@46871.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46873.4]
  assign RetimeWrapper_97_io_in = x526_sum_1_io_result; // @[package.scala 94:16:@46872.4]
  assign RetimeWrapper_98_clock = clock; // @[:@46879.4]
  assign RetimeWrapper_98_reset = reset; // @[:@46880.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46882.4]
  assign RetimeWrapper_98_io_in = ~ x524; // @[package.scala 94:16:@46881.4]
  assign RetimeWrapper_99_clock = clock; // @[:@46891.4]
  assign RetimeWrapper_99_reset = reset; // @[:@46892.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46894.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46893.4]
  assign x531_sum_1_clock = clock; // @[:@46918.4]
  assign x531_sum_1_reset = reset; // @[:@46919.4]
  assign x531_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@46920.4]
  assign x531_sum_1_io_b = x454_div_1_io_result; // @[Math.scala 152:17:@46921.4]
  assign x531_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46922.4]
  assign RetimeWrapper_100_clock = clock; // @[:@46928.4]
  assign RetimeWrapper_100_reset = reset; // @[:@46929.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46931.4]
  assign RetimeWrapper_100_io_in = ~ x529; // @[package.scala 94:16:@46930.4]
  assign RetimeWrapper_101_clock = clock; // @[:@46940.4]
  assign RetimeWrapper_101_reset = reset; // @[:@46941.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46943.4]
  assign RetimeWrapper_101_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46942.4]
  assign x536_sum_1_clock = clock; // @[:@46967.4]
  assign x536_sum_1_reset = reset; // @[:@46968.4]
  assign x536_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@46969.4]
  assign x536_sum_1_io_b = x463_div_1_io_result; // @[Math.scala 152:17:@46970.4]
  assign x536_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@46971.4]
  assign RetimeWrapper_102_clock = clock; // @[:@46977.4]
  assign RetimeWrapper_102_reset = reset; // @[:@46978.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46980.4]
  assign RetimeWrapper_102_io_in = ~ x534; // @[package.scala 94:16:@46979.4]
  assign RetimeWrapper_103_clock = clock; // @[:@46989.4]
  assign RetimeWrapper_103_reset = reset; // @[:@46990.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46992.4]
  assign RetimeWrapper_103_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46991.4]
  assign x544_x13_1_clock = clock; // @[:@47035.4]
  assign x544_x13_1_reset = reset; // @[:@47036.4]
  assign x544_x13_1_io_a = x398_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@47037.4]
  assign x544_x13_1_io_b = _T_1394[31:0]; // @[Math.scala 152:17:@47038.4]
  assign x544_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47039.4]
  assign x545_x14_1_clock = clock; // @[:@47045.4]
  assign x545_x14_1_reset = reset; // @[:@47046.4]
  assign x545_x14_1_io_a = x398_lb_0_io_rPort_13_output_0; // @[Math.scala 151:17:@47047.4]
  assign x545_x14_1_io_b = _T_1397[31:0]; // @[Math.scala 152:17:@47048.4]
  assign x545_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47049.4]
  assign x546_x13_1_clock = clock; // @[:@47055.4]
  assign x546_x13_1_reset = reset; // @[:@47056.4]
  assign x546_x13_1_io_a = _T_1400[31:0]; // @[Math.scala 151:17:@47057.4]
  assign x546_x13_1_io_b = _T_1403[31:0]; // @[Math.scala 152:17:@47058.4]
  assign x546_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47059.4]
  assign x547_x14_1_clock = clock; // @[:@47065.4]
  assign x547_x14_1_reset = reset; // @[:@47066.4]
  assign x547_x14_1_io_a = x398_lb_0_io_rPort_2_output_0; // @[Math.scala 151:17:@47067.4]
  assign x547_x14_1_io_b = _T_1406[31:0]; // @[Math.scala 152:17:@47068.4]
  assign x547_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47069.4]
  assign x548_x13_1_clock = clock; // @[:@47075.4]
  assign x548_x13_1_reset = reset; // @[:@47076.4]
  assign x548_x13_1_io_a = x544_x13_1_io_result; // @[Math.scala 151:17:@47077.4]
  assign x548_x13_1_io_b = x545_x14_1_io_result; // @[Math.scala 152:17:@47078.4]
  assign x548_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47079.4]
  assign x549_x14_1_clock = clock; // @[:@47085.4]
  assign x549_x14_1_reset = reset; // @[:@47086.4]
  assign x549_x14_1_io_a = x546_x13_1_io_result; // @[Math.scala 151:17:@47087.4]
  assign x549_x14_1_io_b = x547_x14_1_io_result; // @[Math.scala 152:17:@47088.4]
  assign x549_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47089.4]
  assign x550_x13_1_clock = clock; // @[:@47095.4]
  assign x550_x13_1_reset = reset; // @[:@47096.4]
  assign x550_x13_1_io_a = x548_x13_1_io_result; // @[Math.scala 151:17:@47097.4]
  assign x550_x13_1_io_b = x549_x14_1_io_result; // @[Math.scala 152:17:@47098.4]
  assign x550_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47099.4]
  assign RetimeWrapper_104_clock = clock; // @[:@47105.4]
  assign RetimeWrapper_104_reset = reset; // @[:@47106.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47108.4]
  assign RetimeWrapper_104_io_in = x398_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@47107.4]
  assign x551_sum_1_clock = clock; // @[:@47114.4]
  assign x551_sum_1_reset = reset; // @[:@47115.4]
  assign x551_sum_1_io_a = x550_x13_1_io_result; // @[Math.scala 151:17:@47116.4]
  assign x551_sum_1_io_b = RetimeWrapper_104_io_out; // @[Math.scala 152:17:@47117.4]
  assign x551_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47118.4]
  assign x552_1_io_b = x551_sum_1_io_result; // @[Math.scala 721:17:@47126.4]
  assign x553_mul_1_clock = clock; // @[:@47135.4]
  assign x553_mul_1_io_a = x552_1_io_result; // @[Math.scala 263:17:@47137.4]
  assign x553_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@47138.4]
  assign x553_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@47139.4]
  assign x554_1_io_b = x553_mul_1_io_result; // @[Math.scala 721:17:@47147.4]
  assign RetimeWrapper_105_clock = clock; // @[:@47154.4]
  assign RetimeWrapper_105_reset = reset; // @[:@47155.4]
  assign RetimeWrapper_105_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47157.4]
  assign RetimeWrapper_105_io_in = x398_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@47156.4]
  assign x555_sub_1_clock = clock; // @[:@47163.4]
  assign x555_sub_1_reset = reset; // @[:@47164.4]
  assign x555_sub_1_io_a = RetimeWrapper_105_io_out; // @[Math.scala 192:17:@47165.4]
  assign x555_sub_1_io_b = x554_1_io_result; // @[Math.scala 193:17:@47166.4]
  assign x555_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47167.4]
  assign RetimeWrapper_106_clock = clock; // @[:@47176.4]
  assign RetimeWrapper_106_reset = reset; // @[:@47177.4]
  assign RetimeWrapper_106_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47179.4]
  assign RetimeWrapper_106_io_in = 32'hf < x555_sub_number; // @[package.scala 94:16:@47178.4]
  assign x557_sub_1_clock = clock; // @[:@47185.4]
  assign x557_sub_1_reset = reset; // @[:@47186.4]
  assign x557_sub_1_io_a = x554_1_io_result; // @[Math.scala 192:17:@47187.4]
  assign x557_sub_1_io_b = RetimeWrapper_105_io_out; // @[Math.scala 193:17:@47188.4]
  assign x557_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47189.4]
  assign RetimeWrapper_107_clock = clock; // @[:@47198.4]
  assign RetimeWrapper_107_reset = reset; // @[:@47199.4]
  assign RetimeWrapper_107_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47201.4]
  assign RetimeWrapper_107_io_in = 32'hf < x557_sub_number; // @[package.scala 94:16:@47200.4]
  assign RetimeWrapper_108_clock = clock; // @[:@47210.4]
  assign RetimeWrapper_108_reset = reset; // @[:@47211.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47213.4]
  assign RetimeWrapper_108_io_in = x555_sub_1_io_result; // @[package.scala 94:16:@47212.4]
  assign x561_1_io_b = x559 ? x800_x555_sub_D1_number : 32'h0; // @[Math.scala 721:17:@47226.4]
  assign x562_mul_1_clock = clock; // @[:@47235.4]
  assign x562_mul_1_io_a = x561_1_io_result; // @[Math.scala 263:17:@47237.4]
  assign x562_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@47238.4]
  assign x562_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@47239.4]
  assign x563_1_io_b = x562_mul_1_io_result; // @[Math.scala 721:17:@47249.4]
  assign RetimeWrapper_109_clock = clock; // @[:@47256.4]
  assign RetimeWrapper_109_reset = reset; // @[:@47257.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47259.4]
  assign RetimeWrapper_109_io_in = x398_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@47258.4]
  assign x564_sum_1_clock = clock; // @[:@47265.4]
  assign x564_sum_1_reset = reset; // @[:@47266.4]
  assign x564_sum_1_io_a = RetimeWrapper_109_io_out; // @[Math.scala 151:17:@47267.4]
  assign x564_sum_1_io_b = x563_1_io_result; // @[Math.scala 152:17:@47268.4]
  assign x564_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47269.4]
  assign x570_x13_1_clock = clock; // @[:@47300.4]
  assign x570_x13_1_reset = reset; // @[:@47301.4]
  assign x570_x13_1_io_a = x398_lb_0_io_rPort_11_output_0; // @[Math.scala 151:17:@47302.4]
  assign x570_x13_1_io_b = _T_1506[31:0]; // @[Math.scala 152:17:@47303.4]
  assign x570_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47304.4]
  assign x571_x14_1_clock = clock; // @[:@47310.4]
  assign x571_x14_1_reset = reset; // @[:@47311.4]
  assign x571_x14_1_io_a = x398_lb_0_io_rPort_9_output_0; // @[Math.scala 151:17:@47312.4]
  assign x571_x14_1_io_b = _T_1509[31:0]; // @[Math.scala 152:17:@47313.4]
  assign x571_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47314.4]
  assign x572_x13_1_clock = clock; // @[:@47320.4]
  assign x572_x13_1_reset = reset; // @[:@47321.4]
  assign x572_x13_1_io_a = _T_1512[31:0]; // @[Math.scala 151:17:@47322.4]
  assign x572_x13_1_io_b = _T_1515[31:0]; // @[Math.scala 152:17:@47323.4]
  assign x572_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47324.4]
  assign x573_x14_1_clock = clock; // @[:@47330.4]
  assign x573_x14_1_reset = reset; // @[:@47331.4]
  assign x573_x14_1_io_a = x398_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@47332.4]
  assign x573_x14_1_io_b = _T_1518[31:0]; // @[Math.scala 152:17:@47333.4]
  assign x573_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47334.4]
  assign x574_x13_1_clock = clock; // @[:@47340.4]
  assign x574_x13_1_reset = reset; // @[:@47341.4]
  assign x574_x13_1_io_a = x570_x13_1_io_result; // @[Math.scala 151:17:@47342.4]
  assign x574_x13_1_io_b = x571_x14_1_io_result; // @[Math.scala 152:17:@47343.4]
  assign x574_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47344.4]
  assign x575_x14_1_clock = clock; // @[:@47350.4]
  assign x575_x14_1_reset = reset; // @[:@47351.4]
  assign x575_x14_1_io_a = x572_x13_1_io_result; // @[Math.scala 151:17:@47352.4]
  assign x575_x14_1_io_b = x573_x14_1_io_result; // @[Math.scala 152:17:@47353.4]
  assign x575_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47354.4]
  assign x576_x13_1_clock = clock; // @[:@47360.4]
  assign x576_x13_1_reset = reset; // @[:@47361.4]
  assign x576_x13_1_io_a = x574_x13_1_io_result; // @[Math.scala 151:17:@47362.4]
  assign x576_x13_1_io_b = x575_x14_1_io_result; // @[Math.scala 152:17:@47363.4]
  assign x576_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47364.4]
  assign RetimeWrapper_110_clock = clock; // @[:@47370.4]
  assign RetimeWrapper_110_reset = reset; // @[:@47371.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47373.4]
  assign RetimeWrapper_110_io_in = x398_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@47372.4]
  assign x577_sum_1_clock = clock; // @[:@47379.4]
  assign x577_sum_1_reset = reset; // @[:@47380.4]
  assign x577_sum_1_io_a = x576_x13_1_io_result; // @[Math.scala 151:17:@47381.4]
  assign x577_sum_1_io_b = RetimeWrapper_110_io_out; // @[Math.scala 152:17:@47382.4]
  assign x577_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47383.4]
  assign x578_1_io_b = x577_sum_1_io_result; // @[Math.scala 721:17:@47391.4]
  assign x579_mul_1_clock = clock; // @[:@47400.4]
  assign x579_mul_1_io_a = x578_1_io_result; // @[Math.scala 263:17:@47402.4]
  assign x579_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@47403.4]
  assign x579_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@47404.4]
  assign x580_1_io_b = x579_mul_1_io_result; // @[Math.scala 721:17:@47412.4]
  assign RetimeWrapper_111_clock = clock; // @[:@47419.4]
  assign RetimeWrapper_111_reset = reset; // @[:@47420.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47422.4]
  assign RetimeWrapper_111_io_in = x398_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@47421.4]
  assign x581_sub_1_clock = clock; // @[:@47428.4]
  assign x581_sub_1_reset = reset; // @[:@47429.4]
  assign x581_sub_1_io_a = RetimeWrapper_111_io_out; // @[Math.scala 192:17:@47430.4]
  assign x581_sub_1_io_b = x580_1_io_result; // @[Math.scala 193:17:@47431.4]
  assign x581_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47432.4]
  assign RetimeWrapper_112_clock = clock; // @[:@47441.4]
  assign RetimeWrapper_112_reset = reset; // @[:@47442.4]
  assign RetimeWrapper_112_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47444.4]
  assign RetimeWrapper_112_io_in = 32'hf < x581_sub_number; // @[package.scala 94:16:@47443.4]
  assign x583_sub_1_clock = clock; // @[:@47450.4]
  assign x583_sub_1_reset = reset; // @[:@47451.4]
  assign x583_sub_1_io_a = x580_1_io_result; // @[Math.scala 192:17:@47452.4]
  assign x583_sub_1_io_b = RetimeWrapper_111_io_out; // @[Math.scala 193:17:@47453.4]
  assign x583_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47454.4]
  assign RetimeWrapper_113_clock = clock; // @[:@47463.4]
  assign RetimeWrapper_113_reset = reset; // @[:@47464.4]
  assign RetimeWrapper_113_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47466.4]
  assign RetimeWrapper_113_io_in = 32'hf < x583_sub_number; // @[package.scala 94:16:@47465.4]
  assign RetimeWrapper_114_clock = clock; // @[:@47475.4]
  assign RetimeWrapper_114_reset = reset; // @[:@47476.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47478.4]
  assign RetimeWrapper_114_io_in = x581_sub_1_io_result; // @[package.scala 94:16:@47477.4]
  assign x587_1_io_b = x585 ? x804_x581_sub_D1_number : 32'h0; // @[Math.scala 721:17:@47491.4]
  assign x588_mul_1_clock = clock; // @[:@47500.4]
  assign x588_mul_1_io_a = x587_1_io_result; // @[Math.scala 263:17:@47502.4]
  assign x588_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@47503.4]
  assign x588_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@47504.4]
  assign x589_1_io_b = x588_mul_1_io_result; // @[Math.scala 721:17:@47512.4]
  assign RetimeWrapper_115_clock = clock; // @[:@47519.4]
  assign RetimeWrapper_115_reset = reset; // @[:@47520.4]
  assign RetimeWrapper_115_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47522.4]
  assign RetimeWrapper_115_io_in = x398_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@47521.4]
  assign x590_sum_1_clock = clock; // @[:@47528.4]
  assign x590_sum_1_reset = reset; // @[:@47529.4]
  assign x590_sum_1_io_a = RetimeWrapper_115_io_out; // @[Math.scala 151:17:@47530.4]
  assign x590_sum_1_io_b = x589_1_io_result; // @[Math.scala 152:17:@47531.4]
  assign x590_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47532.4]
  assign x595_x13_1_clock = clock; // @[:@47558.4]
  assign x595_x13_1_reset = reset; // @[:@47559.4]
  assign x595_x13_1_io_a = x398_lb_0_io_rPort_13_output_0; // @[Math.scala 151:17:@47560.4]
  assign x595_x13_1_io_b = _T_1616[31:0]; // @[Math.scala 152:17:@47561.4]
  assign x595_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47562.4]
  assign x596_x14_1_clock = clock; // @[:@47568.4]
  assign x596_x14_1_reset = reset; // @[:@47569.4]
  assign x596_x14_1_io_a = x398_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@47570.4]
  assign x596_x14_1_io_b = _T_1403[31:0]; // @[Math.scala 152:17:@47571.4]
  assign x596_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47572.4]
  assign x597_x13_1_clock = clock; // @[:@47578.4]
  assign x597_x13_1_reset = reset; // @[:@47579.4]
  assign x597_x13_1_io_a = _T_1619[31:0]; // @[Math.scala 151:17:@47580.4]
  assign x597_x13_1_io_b = _T_1622[31:0]; // @[Math.scala 152:17:@47581.4]
  assign x597_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47582.4]
  assign x598_x14_1_clock = clock; // @[:@47588.4]
  assign x598_x14_1_reset = reset; // @[:@47589.4]
  assign x598_x14_1_io_a = x398_lb_0_io_rPort_3_output_0; // @[Math.scala 151:17:@47590.4]
  assign x598_x14_1_io_b = _T_1625[31:0]; // @[Math.scala 152:17:@47591.4]
  assign x598_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47592.4]
  assign x599_x13_1_clock = clock; // @[:@47598.4]
  assign x599_x13_1_reset = reset; // @[:@47599.4]
  assign x599_x13_1_io_a = x595_x13_1_io_result; // @[Math.scala 151:17:@47600.4]
  assign x599_x13_1_io_b = x596_x14_1_io_result; // @[Math.scala 152:17:@47601.4]
  assign x599_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47602.4]
  assign x600_x14_1_clock = clock; // @[:@47608.4]
  assign x600_x14_1_reset = reset; // @[:@47609.4]
  assign x600_x14_1_io_a = x597_x13_1_io_result; // @[Math.scala 151:17:@47610.4]
  assign x600_x14_1_io_b = x598_x14_1_io_result; // @[Math.scala 152:17:@47611.4]
  assign x600_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47612.4]
  assign x601_x13_1_clock = clock; // @[:@47618.4]
  assign x601_x13_1_reset = reset; // @[:@47619.4]
  assign x601_x13_1_io_a = x599_x13_1_io_result; // @[Math.scala 151:17:@47620.4]
  assign x601_x13_1_io_b = x600_x14_1_io_result; // @[Math.scala 152:17:@47621.4]
  assign x601_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47622.4]
  assign RetimeWrapper_116_clock = clock; // @[:@47628.4]
  assign RetimeWrapper_116_reset = reset; // @[:@47629.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47631.4]
  assign RetimeWrapper_116_io_in = x398_lb_0_io_rPort_12_output_0; // @[package.scala 94:16:@47630.4]
  assign x602_sum_1_clock = clock; // @[:@47637.4]
  assign x602_sum_1_reset = reset; // @[:@47638.4]
  assign x602_sum_1_io_a = x601_x13_1_io_result; // @[Math.scala 151:17:@47639.4]
  assign x602_sum_1_io_b = RetimeWrapper_116_io_out; // @[Math.scala 152:17:@47640.4]
  assign x602_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47641.4]
  assign x603_1_io_b = x602_sum_1_io_result; // @[Math.scala 721:17:@47649.4]
  assign x604_mul_1_clock = clock; // @[:@47658.4]
  assign x604_mul_1_io_a = x603_1_io_result; // @[Math.scala 263:17:@47660.4]
  assign x604_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@47661.4]
  assign x604_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@47662.4]
  assign x605_1_io_b = x604_mul_1_io_result; // @[Math.scala 721:17:@47670.4]
  assign RetimeWrapper_117_clock = clock; // @[:@47677.4]
  assign RetimeWrapper_117_reset = reset; // @[:@47678.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47680.4]
  assign RetimeWrapper_117_io_in = x398_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@47679.4]
  assign x606_sub_1_clock = clock; // @[:@47688.4]
  assign x606_sub_1_reset = reset; // @[:@47689.4]
  assign x606_sub_1_io_a = RetimeWrapper_117_io_out; // @[Math.scala 192:17:@47690.4]
  assign x606_sub_1_io_b = x605_1_io_result; // @[Math.scala 193:17:@47691.4]
  assign x606_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47692.4]
  assign RetimeWrapper_118_clock = clock; // @[:@47701.4]
  assign RetimeWrapper_118_reset = reset; // @[:@47702.4]
  assign RetimeWrapper_118_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47704.4]
  assign RetimeWrapper_118_io_in = 32'hf < x606_sub_number; // @[package.scala 94:16:@47703.4]
  assign x608_sub_1_clock = clock; // @[:@47710.4]
  assign x608_sub_1_reset = reset; // @[:@47711.4]
  assign x608_sub_1_io_a = x605_1_io_result; // @[Math.scala 192:17:@47712.4]
  assign x608_sub_1_io_b = RetimeWrapper_117_io_out; // @[Math.scala 193:17:@47713.4]
  assign x608_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47714.4]
  assign RetimeWrapper_119_clock = clock; // @[:@47723.4]
  assign RetimeWrapper_119_reset = reset; // @[:@47724.4]
  assign RetimeWrapper_119_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47726.4]
  assign RetimeWrapper_119_io_in = 32'hf < x608_sub_number; // @[package.scala 94:16:@47725.4]
  assign RetimeWrapper_120_clock = clock; // @[:@47735.4]
  assign RetimeWrapper_120_reset = reset; // @[:@47736.4]
  assign RetimeWrapper_120_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47738.4]
  assign RetimeWrapper_120_io_in = x606_sub_1_io_result; // @[package.scala 94:16:@47737.4]
  assign x612_1_io_b = x610 ? x808_x606_sub_D1_number : 32'h0; // @[Math.scala 721:17:@47751.4]
  assign x613_mul_1_clock = clock; // @[:@47760.4]
  assign x613_mul_1_io_a = x612_1_io_result; // @[Math.scala 263:17:@47762.4]
  assign x613_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@47763.4]
  assign x613_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@47764.4]
  assign x614_1_io_b = x613_mul_1_io_result; // @[Math.scala 721:17:@47772.4]
  assign RetimeWrapper_121_clock = clock; // @[:@47779.4]
  assign RetimeWrapper_121_reset = reset; // @[:@47780.4]
  assign RetimeWrapper_121_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47782.4]
  assign RetimeWrapper_121_io_in = x398_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@47781.4]
  assign x615_sum_1_clock = clock; // @[:@47788.4]
  assign x615_sum_1_reset = reset; // @[:@47789.4]
  assign x615_sum_1_io_a = RetimeWrapper_121_io_out; // @[Math.scala 151:17:@47790.4]
  assign x615_sum_1_io_b = x614_1_io_result; // @[Math.scala 152:17:@47791.4]
  assign x615_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47792.4]
  assign x620_x13_1_clock = clock; // @[:@47818.4]
  assign x620_x13_1_reset = reset; // @[:@47819.4]
  assign x620_x13_1_io_a = x398_lb_0_io_rPort_9_output_0; // @[Math.scala 151:17:@47820.4]
  assign x620_x13_1_io_b = _T_1725[31:0]; // @[Math.scala 152:17:@47821.4]
  assign x620_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47822.4]
  assign x621_x14_1_clock = clock; // @[:@47828.4]
  assign x621_x14_1_reset = reset; // @[:@47829.4]
  assign x621_x14_1_io_a = x398_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@47830.4]
  assign x621_x14_1_io_b = _T_1515[31:0]; // @[Math.scala 152:17:@47831.4]
  assign x621_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47832.4]
  assign x622_x13_1_clock = clock; // @[:@47838.4]
  assign x622_x13_1_reset = reset; // @[:@47839.4]
  assign x622_x13_1_io_a = _T_1728[31:0]; // @[Math.scala 151:17:@47840.4]
  assign x622_x13_1_io_b = _T_1731[31:0]; // @[Math.scala 152:17:@47841.4]
  assign x622_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47842.4]
  assign x623_x14_1_clock = clock; // @[:@47848.4]
  assign x623_x14_1_reset = reset; // @[:@47849.4]
  assign x623_x14_1_io_a = x398_lb_0_io_rPort_1_output_0; // @[Math.scala 151:17:@47850.4]
  assign x623_x14_1_io_b = _T_1734[31:0]; // @[Math.scala 152:17:@47851.4]
  assign x623_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47852.4]
  assign x624_x13_1_clock = clock; // @[:@47858.4]
  assign x624_x13_1_reset = reset; // @[:@47859.4]
  assign x624_x13_1_io_a = x620_x13_1_io_result; // @[Math.scala 151:17:@47860.4]
  assign x624_x13_1_io_b = x621_x14_1_io_result; // @[Math.scala 152:17:@47861.4]
  assign x624_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47862.4]
  assign x625_x14_1_clock = clock; // @[:@47868.4]
  assign x625_x14_1_reset = reset; // @[:@47869.4]
  assign x625_x14_1_io_a = x622_x13_1_io_result; // @[Math.scala 151:17:@47870.4]
  assign x625_x14_1_io_b = x623_x14_1_io_result; // @[Math.scala 152:17:@47871.4]
  assign x625_x14_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47872.4]
  assign x626_x13_1_clock = clock; // @[:@47878.4]
  assign x626_x13_1_reset = reset; // @[:@47879.4]
  assign x626_x13_1_io_a = x624_x13_1_io_result; // @[Math.scala 151:17:@47880.4]
  assign x626_x13_1_io_b = x625_x14_1_io_result; // @[Math.scala 152:17:@47881.4]
  assign x626_x13_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47882.4]
  assign RetimeWrapper_122_clock = clock; // @[:@47888.4]
  assign RetimeWrapper_122_reset = reset; // @[:@47889.4]
  assign RetimeWrapper_122_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47891.4]
  assign RetimeWrapper_122_io_in = x398_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@47890.4]
  assign x627_sum_1_clock = clock; // @[:@47897.4]
  assign x627_sum_1_reset = reset; // @[:@47898.4]
  assign x627_sum_1_io_a = x626_x13_1_io_result; // @[Math.scala 151:17:@47899.4]
  assign x627_sum_1_io_b = RetimeWrapper_122_io_out; // @[Math.scala 152:17:@47900.4]
  assign x627_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@47901.4]
  assign x628_1_io_b = x627_sum_1_io_result; // @[Math.scala 721:17:@47909.4]
  assign x629_mul_1_clock = clock; // @[:@47918.4]
  assign x629_mul_1_io_a = x628_1_io_result; // @[Math.scala 263:17:@47920.4]
  assign x629_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@47921.4]
  assign x629_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@47922.4]
  assign x630_1_io_b = x629_mul_1_io_result; // @[Math.scala 721:17:@47930.4]
  assign RetimeWrapper_123_clock = clock; // @[:@47937.4]
  assign RetimeWrapper_123_reset = reset; // @[:@47938.4]
  assign RetimeWrapper_123_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47940.4]
  assign RetimeWrapper_123_io_in = x398_lb_0_io_rPort_9_output_0; // @[package.scala 94:16:@47939.4]
  assign x631_sub_1_clock = clock; // @[:@47946.4]
  assign x631_sub_1_reset = reset; // @[:@47947.4]
  assign x631_sub_1_io_a = RetimeWrapper_123_io_out; // @[Math.scala 192:17:@47948.4]
  assign x631_sub_1_io_b = x630_1_io_result; // @[Math.scala 193:17:@47949.4]
  assign x631_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47950.4]
  assign RetimeWrapper_124_clock = clock; // @[:@47959.4]
  assign RetimeWrapper_124_reset = reset; // @[:@47960.4]
  assign RetimeWrapper_124_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47962.4]
  assign RetimeWrapper_124_io_in = 32'hf < x631_sub_number; // @[package.scala 94:16:@47961.4]
  assign x633_sub_1_clock = clock; // @[:@47968.4]
  assign x633_sub_1_reset = reset; // @[:@47969.4]
  assign x633_sub_1_io_a = x630_1_io_result; // @[Math.scala 192:17:@47970.4]
  assign x633_sub_1_io_b = RetimeWrapper_123_io_out; // @[Math.scala 193:17:@47971.4]
  assign x633_sub_1_io_flow = io_in_x354_TREADY; // @[Math.scala 194:20:@47972.4]
  assign RetimeWrapper_125_clock = clock; // @[:@47981.4]
  assign RetimeWrapper_125_reset = reset; // @[:@47982.4]
  assign RetimeWrapper_125_io_flow = io_in_x354_TREADY; // @[package.scala 95:18:@47984.4]
  assign RetimeWrapper_125_io_in = 32'hf < x633_sub_number; // @[package.scala 94:16:@47983.4]
  assign RetimeWrapper_126_clock = clock; // @[:@47993.4]
  assign RetimeWrapper_126_reset = reset; // @[:@47994.4]
  assign RetimeWrapper_126_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47996.4]
  assign RetimeWrapper_126_io_in = x631_sub_1_io_result; // @[package.scala 94:16:@47995.4]
  assign x637_1_io_b = x635 ? x812_x631_sub_D1_number : 32'h0; // @[Math.scala 721:17:@48009.4]
  assign x638_mul_1_clock = clock; // @[:@48018.4]
  assign x638_mul_1_io_a = x637_1_io_result; // @[Math.scala 263:17:@48020.4]
  assign x638_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@48021.4]
  assign x638_mul_1_io_flow = io_in_x354_TREADY; // @[Math.scala 265:20:@48022.4]
  assign x639_1_io_b = x638_mul_1_io_result; // @[Math.scala 721:17:@48030.4]
  assign RetimeWrapper_127_clock = clock; // @[:@48037.4]
  assign RetimeWrapper_127_reset = reset; // @[:@48038.4]
  assign RetimeWrapper_127_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48040.4]
  assign RetimeWrapper_127_io_in = x398_lb_0_io_rPort_9_output_0; // @[package.scala 94:16:@48039.4]
  assign x640_sum_1_clock = clock; // @[:@48046.4]
  assign x640_sum_1_reset = reset; // @[:@48047.4]
  assign x640_sum_1_io_a = RetimeWrapper_127_io_out; // @[Math.scala 151:17:@48048.4]
  assign x640_sum_1_io_b = x639_1_io_result; // @[Math.scala 152:17:@48049.4]
  assign x640_sum_1_io_flow = io_in_x354_TREADY; // @[Math.scala 153:20:@48050.4]
  assign RetimeWrapper_128_clock = clock; // @[:@48066.4]
  assign RetimeWrapper_128_reset = reset; // @[:@48067.4]
  assign RetimeWrapper_128_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48069.4]
  assign RetimeWrapper_128_io_in = {_T_1842,_T_1841}; // @[package.scala 94:16:@48068.4]
  assign RetimeWrapper_129_clock = clock; // @[:@48075.4]
  assign RetimeWrapper_129_reset = reset; // @[:@48076.4]
  assign RetimeWrapper_129_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48078.4]
  assign RetimeWrapper_129_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@48077.4]
  assign RetimeWrapper_130_clock = clock; // @[:@48084.4]
  assign RetimeWrapper_130_reset = reset; // @[:@48085.4]
  assign RetimeWrapper_130_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48087.4]
  assign RetimeWrapper_130_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@48086.4]
  assign RetimeWrapper_131_clock = clock; // @[:@48093.4]
  assign RetimeWrapper_131_reset = reset; // @[:@48094.4]
  assign RetimeWrapper_131_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48096.4]
  assign RetimeWrapper_131_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@48095.4]
endmodule
module x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1( // @[:@48114.2]
  input          clock, // @[:@48115.4]
  input          reset, // @[:@48116.4]
  input          io_in_x353_TVALID, // @[:@48117.4]
  output         io_in_x353_TREADY, // @[:@48117.4]
  input  [255:0] io_in_x353_TDATA, // @[:@48117.4]
  input  [7:0]   io_in_x353_TID, // @[:@48117.4]
  input  [7:0]   io_in_x353_TDEST, // @[:@48117.4]
  output         io_in_x354_TVALID, // @[:@48117.4]
  input          io_in_x354_TREADY, // @[:@48117.4]
  output [255:0] io_in_x354_TDATA, // @[:@48117.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@48117.4]
  input          io_sigsIn_smChildAcks_0, // @[:@48117.4]
  output         io_sigsOut_smDoneIn_0, // @[:@48117.4]
  input          io_rr // @[:@48117.4]
);
  wire  x391_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire  x391_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire  x391_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire  x391_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire [12:0] x391_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire [12:0] x391_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire  x391_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire  x391_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire  x391_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@48151.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48239.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48239.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48239.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@48239.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@48239.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48281.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48281.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48281.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48281.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48281.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@48289.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@48289.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@48289.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@48289.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@48289.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TREADY; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire [255:0] x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TDATA; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire [7:0] x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TID; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire [7:0] x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TDEST; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TVALID; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TREADY; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire [255:0] x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TDATA; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire [31:0] x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire [31:0] x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
  wire  _T_240; // @[package.scala 96:25:@48244.4 package.scala 96:25:@48245.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x646_outr_UnitPipe.scala 69:66:@48250.4]
  wire  _T_253; // @[package.scala 96:25:@48286.4 package.scala 96:25:@48287.4]
  wire  _T_259; // @[package.scala 96:25:@48294.4 package.scala 96:25:@48295.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@48297.4]
  wire  x645_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@48298.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@48306.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@48307.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@48319.4]
  x361_ctrchain x391_ctrchain ( // @[SpatialBlocks.scala 37:22:@48151.4]
    .clock(x391_ctrchain_clock),
    .reset(x391_ctrchain_reset),
    .io_input_reset(x391_ctrchain_io_input_reset),
    .io_input_enable(x391_ctrchain_io_input_enable),
    .io_output_counts_1(x391_ctrchain_io_output_counts_1),
    .io_output_counts_0(x391_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x391_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x391_ctrchain_io_output_oobs_1),
    .io_output_done(x391_ctrchain_io_output_done)
  );
  x645_inr_Foreach_SAMPLER_BOX_sm x645_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 32:18:@48211.4]
    .clock(x645_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x645_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x645_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x645_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x645_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x645_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x645_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x645_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x645_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@48239.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@48281.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@48289.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1 x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 876:24:@48323.4]
    .clock(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x353_TREADY(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TREADY),
    .io_in_x353_TDATA(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TDATA),
    .io_in_x353_TID(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TID),
    .io_in_x353_TDEST(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TDEST),
    .io_in_x354_TVALID(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TVALID),
    .io_in_x354_TREADY(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TREADY),
    .io_in_x354_TDATA(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TDATA),
    .io_sigsIn_backpressure(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@48244.4 package.scala 96:25:@48245.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x353_TVALID | x645_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x646_outr_UnitPipe.scala 69:66:@48250.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@48286.4 package.scala 96:25:@48287.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@48294.4 package.scala 96:25:@48295.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@48297.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@48298.4]
  assign _T_264 = x645_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@48306.4]
  assign _T_265 = ~ x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@48307.4]
  assign _T_272 = x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@48319.4]
  assign io_in_x353_TREADY = x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TREADY; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 48:23:@48381.4]
  assign io_in_x354_TVALID = x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TVALID; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 49:23:@48391.4]
  assign io_in_x354_TDATA = x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TDATA; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 49:23:@48389.4]
  assign io_sigsOut_smDoneIn_0 = x645_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@48304.4]
  assign x391_ctrchain_clock = clock; // @[:@48152.4]
  assign x391_ctrchain_reset = reset; // @[:@48153.4]
  assign x391_ctrchain_io_input_reset = x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@48322.4]
  assign x391_ctrchain_io_input_enable = _T_272 & x645_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@48274.4 SpatialBlocks.scala 159:42:@48321.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@48212.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@48213.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sm_io_enable = x645_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x645_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@48301.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x646_outr_UnitPipe.scala 67:50:@48247.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@48303.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x354_TREADY | x645_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@48275.4]
  assign x645_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x646_outr_UnitPipe.scala 71:48:@48253.4]
  assign RetimeWrapper_clock = clock; // @[:@48240.4]
  assign RetimeWrapper_reset = reset; // @[:@48241.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48243.4]
  assign RetimeWrapper_io_in = x391_ctrchain_io_output_done; // @[package.scala 94:16:@48242.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48282.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48283.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48285.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@48284.4]
  assign RetimeWrapper_2_clock = clock; // @[:@48290.4]
  assign RetimeWrapper_2_reset = reset; // @[:@48291.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@48293.4]
  assign RetimeWrapper_2_io_in = x645_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@48292.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@48324.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@48325.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TDATA = io_in_x353_TDATA; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 48:23:@48380.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TID = io_in_x353_TID; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 48:23:@48376.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x353_TDEST = io_in_x353_TDEST; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 48:23:@48375.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x354_TREADY = io_in_x354_TREADY; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 49:23:@48390.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x354_TREADY | x645_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 881:22:@48408.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 881:22:@48406.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x645_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 881:22:@48404.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x391_ctrchain_io_output_counts_1[12]}},x391_ctrchain_io_output_counts_1}; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 881:22:@48399.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x391_ctrchain_io_output_counts_0[12]}},x391_ctrchain_io_output_counts_0}; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 881:22:@48398.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x391_ctrchain_io_output_oobs_0; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 881:22:@48396.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x391_ctrchain_io_output_oobs_1; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 881:22:@48397.4]
  assign x645_inr_Foreach_SAMPLER_BOX_kernelx645_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x645_inr_Foreach_SAMPLER_BOX.scala 880:18:@48392.4]
endmodule
module x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1( // @[:@48422.2]
  input          clock, // @[:@48423.4]
  input          reset, // @[:@48424.4]
  input          io_in_x353_TVALID, // @[:@48425.4]
  output         io_in_x353_TREADY, // @[:@48425.4]
  input  [255:0] io_in_x353_TDATA, // @[:@48425.4]
  input  [7:0]   io_in_x353_TID, // @[:@48425.4]
  input  [7:0]   io_in_x353_TDEST, // @[:@48425.4]
  output         io_in_x354_TVALID, // @[:@48425.4]
  input          io_in_x354_TREADY, // @[:@48425.4]
  output [255:0] io_in_x354_TDATA, // @[:@48425.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@48425.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@48425.4]
  input          io_sigsIn_smChildAcks_0, // @[:@48425.4]
  input          io_sigsIn_smChildAcks_1, // @[:@48425.4]
  output         io_sigsOut_smDoneIn_0, // @[:@48425.4]
  output         io_sigsOut_smDoneIn_1, // @[:@48425.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@48425.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@48425.4]
  input          io_rr // @[:@48425.4]
);
  wire  x356_fifoinraw_0_clock; // @[m_x356_fifoinraw_0.scala 27:17:@48439.4]
  wire  x356_fifoinraw_0_reset; // @[m_x356_fifoinraw_0.scala 27:17:@48439.4]
  wire  x357_fifoinpacked_0_clock; // @[m_x357_fifoinpacked_0.scala 27:17:@48463.4]
  wire  x357_fifoinpacked_0_reset; // @[m_x357_fifoinpacked_0.scala 27:17:@48463.4]
  wire  x357_fifoinpacked_0_io_wPort_0_en_0; // @[m_x357_fifoinpacked_0.scala 27:17:@48463.4]
  wire  x357_fifoinpacked_0_io_full; // @[m_x357_fifoinpacked_0.scala 27:17:@48463.4]
  wire  x357_fifoinpacked_0_io_active_0_in; // @[m_x357_fifoinpacked_0.scala 27:17:@48463.4]
  wire  x357_fifoinpacked_0_io_active_0_out; // @[m_x357_fifoinpacked_0.scala 27:17:@48463.4]
  wire  x358_fifooutraw_0_clock; // @[m_x358_fifooutraw_0.scala 27:17:@48487.4]
  wire  x358_fifooutraw_0_reset; // @[m_x358_fifooutraw_0.scala 27:17:@48487.4]
  wire  x361_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire  x361_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire  x361_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire  x361_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire [12:0] x361_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire [12:0] x361_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire  x361_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire  x361_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire  x361_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@48511.4]
  wire  x387_inr_Foreach_sm_clock; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_reset; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_enable; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_done; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_doneLatch; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_ctrDone; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_datapathEn; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_ctrInc; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_ctrRst; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_parentAck; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_backpressure; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  x387_inr_Foreach_sm_io_break; // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48599.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48599.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48599.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@48599.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@48599.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48645.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48645.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48645.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48645.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48645.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@48653.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@48653.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@48653.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@48653.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@48653.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_clock; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_reset; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_wPort_0_en_0; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_full; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_active_0_in; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_active_0_out; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire [31:0] x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire [31:0] x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_rr; // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
  wire  x646_outr_UnitPipe_sm_clock; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_reset; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_enable; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_done; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_rst; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_ctrDone; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_ctrInc; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_parentAck; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  x646_outr_UnitPipe_sm_io_childAck_0; // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@48885.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@48885.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@48885.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@48885.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@48885.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_clock; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_reset; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TVALID; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TREADY; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire [255:0] x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TDATA; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire [7:0] x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TID; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire [7:0] x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TDEST; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TVALID; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TREADY; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire [255:0] x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TDATA; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_rr; // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
  wire  _T_254; // @[package.scala 96:25:@48604.4 package.scala 96:25:@48605.4]
  wire  _T_260; // @[implicits.scala 47:10:@48608.4]
  wire  _T_261; // @[sm_x647_outr_UnitPipe.scala 70:41:@48609.4]
  wire  _T_262; // @[sm_x647_outr_UnitPipe.scala 70:78:@48610.4]
  wire  _T_263; // @[sm_x647_outr_UnitPipe.scala 70:76:@48611.4]
  wire  _T_275; // @[package.scala 96:25:@48650.4 package.scala 96:25:@48651.4]
  wire  _T_281; // @[package.scala 96:25:@48658.4 package.scala 96:25:@48659.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@48661.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@48670.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@48671.4]
  wire  _T_354; // @[package.scala 100:49:@48848.4]
  reg  _T_357; // @[package.scala 48:56:@48849.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@48882.4 package.scala 96:25:@48883.4]
  wire  _T_377; // @[package.scala 96:25:@48890.4 package.scala 96:25:@48891.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@48893.4]
  x356_fifoinraw_0 x356_fifoinraw_0 ( // @[m_x356_fifoinraw_0.scala 27:17:@48439.4]
    .clock(x356_fifoinraw_0_clock),
    .reset(x356_fifoinraw_0_reset)
  );
  x357_fifoinpacked_0 x357_fifoinpacked_0 ( // @[m_x357_fifoinpacked_0.scala 27:17:@48463.4]
    .clock(x357_fifoinpacked_0_clock),
    .reset(x357_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x357_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x357_fifoinpacked_0_io_full),
    .io_active_0_in(x357_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x357_fifoinpacked_0_io_active_0_out)
  );
  x356_fifoinraw_0 x358_fifooutraw_0 ( // @[m_x358_fifooutraw_0.scala 27:17:@48487.4]
    .clock(x358_fifooutraw_0_clock),
    .reset(x358_fifooutraw_0_reset)
  );
  x361_ctrchain x361_ctrchain ( // @[SpatialBlocks.scala 37:22:@48511.4]
    .clock(x361_ctrchain_clock),
    .reset(x361_ctrchain_reset),
    .io_input_reset(x361_ctrchain_io_input_reset),
    .io_input_enable(x361_ctrchain_io_input_enable),
    .io_output_counts_1(x361_ctrchain_io_output_counts_1),
    .io_output_counts_0(x361_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x361_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x361_ctrchain_io_output_oobs_1),
    .io_output_done(x361_ctrchain_io_output_done)
  );
  x387_inr_Foreach_sm x387_inr_Foreach_sm ( // @[sm_x387_inr_Foreach.scala 32:18:@48571.4]
    .clock(x387_inr_Foreach_sm_clock),
    .reset(x387_inr_Foreach_sm_reset),
    .io_enable(x387_inr_Foreach_sm_io_enable),
    .io_done(x387_inr_Foreach_sm_io_done),
    .io_doneLatch(x387_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x387_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x387_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x387_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x387_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x387_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x387_inr_Foreach_sm_io_backpressure),
    .io_break(x387_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@48599.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@48645.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@48653.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x387_inr_Foreach_kernelx387_inr_Foreach_concrete1 x387_inr_Foreach_kernelx387_inr_Foreach_concrete1 ( // @[sm_x387_inr_Foreach.scala 126:24:@48688.4]
    .clock(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_clock),
    .reset(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_reset),
    .io_in_x357_fifoinpacked_0_wPort_0_en_0(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_wPort_0_en_0),
    .io_in_x357_fifoinpacked_0_full(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_full),
    .io_in_x357_fifoinpacked_0_active_0_in(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_active_0_in),
    .io_in_x357_fifoinpacked_0_active_0_out(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x646_outr_UnitPipe_sm ( // @[sm_x646_outr_UnitPipe.scala 32:18:@48820.4]
    .clock(x646_outr_UnitPipe_sm_clock),
    .reset(x646_outr_UnitPipe_sm_reset),
    .io_enable(x646_outr_UnitPipe_sm_io_enable),
    .io_done(x646_outr_UnitPipe_sm_io_done),
    .io_rst(x646_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x646_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x646_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x646_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x646_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x646_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x646_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@48877.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@48885.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1 x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1 ( // @[sm_x646_outr_UnitPipe.scala 76:24:@48915.4]
    .clock(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_clock),
    .reset(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_reset),
    .io_in_x353_TVALID(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TVALID),
    .io_in_x353_TREADY(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TREADY),
    .io_in_x353_TDATA(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TDATA),
    .io_in_x353_TID(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TID),
    .io_in_x353_TDEST(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TDEST),
    .io_in_x354_TVALID(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TVALID),
    .io_in_x354_TREADY(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TREADY),
    .io_in_x354_TDATA(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TDATA),
    .io_sigsIn_smEnableOuts_0(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@48604.4 package.scala 96:25:@48605.4]
  assign _T_260 = x357_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@48608.4]
  assign _T_261 = ~ _T_260; // @[sm_x647_outr_UnitPipe.scala 70:41:@48609.4]
  assign _T_262 = ~ x357_fifoinpacked_0_io_active_0_out; // @[sm_x647_outr_UnitPipe.scala 70:78:@48610.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x647_outr_UnitPipe.scala 70:76:@48611.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@48650.4 package.scala 96:25:@48651.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@48658.4 package.scala 96:25:@48659.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@48661.4]
  assign _T_286 = x387_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@48670.4]
  assign _T_287 = ~ x387_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@48671.4]
  assign _T_354 = x646_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@48848.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@48882.4 package.scala 96:25:@48883.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@48890.4 package.scala 96:25:@48891.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@48893.4]
  assign io_in_x353_TREADY = x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TREADY; // @[sm_x646_outr_UnitPipe.scala 48:23:@48971.4]
  assign io_in_x354_TVALID = x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TVALID; // @[sm_x646_outr_UnitPipe.scala 49:23:@48981.4]
  assign io_in_x354_TDATA = x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TDATA; // @[sm_x646_outr_UnitPipe.scala 49:23:@48979.4]
  assign io_sigsOut_smDoneIn_0 = x387_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@48668.4]
  assign io_sigsOut_smDoneIn_1 = x646_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@48900.4]
  assign io_sigsOut_smCtrCopyDone_0 = x387_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@48687.4]
  assign io_sigsOut_smCtrCopyDone_1 = x646_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@48914.4]
  assign x356_fifoinraw_0_clock = clock; // @[:@48440.4]
  assign x356_fifoinraw_0_reset = reset; // @[:@48441.4]
  assign x357_fifoinpacked_0_clock = clock; // @[:@48464.4]
  assign x357_fifoinpacked_0_reset = reset; // @[:@48465.4]
  assign x357_fifoinpacked_0_io_wPort_0_en_0 = x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@48748.4]
  assign x357_fifoinpacked_0_io_active_0_in = x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@48747.4]
  assign x358_fifooutraw_0_clock = clock; // @[:@48488.4]
  assign x358_fifooutraw_0_reset = reset; // @[:@48489.4]
  assign x361_ctrchain_clock = clock; // @[:@48512.4]
  assign x361_ctrchain_reset = reset; // @[:@48513.4]
  assign x361_ctrchain_io_input_reset = x387_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@48686.4]
  assign x361_ctrchain_io_input_enable = x387_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@48638.4 SpatialBlocks.scala 159:42:@48685.4]
  assign x387_inr_Foreach_sm_clock = clock; // @[:@48572.4]
  assign x387_inr_Foreach_sm_reset = reset; // @[:@48573.4]
  assign x387_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@48665.4]
  assign x387_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x647_outr_UnitPipe.scala 69:38:@48607.4]
  assign x387_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@48667.4]
  assign x387_inr_Foreach_sm_io_backpressure = _T_263 | x387_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@48639.4]
  assign x387_inr_Foreach_sm_io_break = 1'h0; // @[sm_x647_outr_UnitPipe.scala 73:36:@48617.4]
  assign RetimeWrapper_clock = clock; // @[:@48600.4]
  assign RetimeWrapper_reset = reset; // @[:@48601.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48603.4]
  assign RetimeWrapper_io_in = x361_ctrchain_io_output_done; // @[package.scala 94:16:@48602.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48646.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48647.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48649.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@48648.4]
  assign RetimeWrapper_2_clock = clock; // @[:@48654.4]
  assign RetimeWrapper_2_reset = reset; // @[:@48655.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@48657.4]
  assign RetimeWrapper_2_io_in = x387_inr_Foreach_sm_io_done; // @[package.scala 94:16:@48656.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_clock = clock; // @[:@48689.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_reset = reset; // @[:@48690.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_full = x357_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@48742.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_in_x357_fifoinpacked_0_active_0_out = x357_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@48741.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x387_inr_Foreach_sm_io_doneLatch; // @[sm_x387_inr_Foreach.scala 131:22:@48771.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x387_inr_Foreach.scala 131:22:@48769.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_break = x387_inr_Foreach_sm_io_break; // @[sm_x387_inr_Foreach.scala 131:22:@48767.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x361_ctrchain_io_output_counts_1[12]}},x361_ctrchain_io_output_counts_1}; // @[sm_x387_inr_Foreach.scala 131:22:@48762.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x361_ctrchain_io_output_counts_0[12]}},x361_ctrchain_io_output_counts_0}; // @[sm_x387_inr_Foreach.scala 131:22:@48761.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x361_ctrchain_io_output_oobs_0; // @[sm_x387_inr_Foreach.scala 131:22:@48759.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x361_ctrchain_io_output_oobs_1; // @[sm_x387_inr_Foreach.scala 131:22:@48760.4]
  assign x387_inr_Foreach_kernelx387_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x387_inr_Foreach.scala 130:18:@48755.4]
  assign x646_outr_UnitPipe_sm_clock = clock; // @[:@48821.4]
  assign x646_outr_UnitPipe_sm_reset = reset; // @[:@48822.4]
  assign x646_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@48897.4]
  assign x646_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@48872.4]
  assign x646_outr_UnitPipe_sm_io_ctrDone = x646_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x647_outr_UnitPipe.scala 78:40:@48852.4]
  assign x646_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@48899.4]
  assign x646_outr_UnitPipe_sm_io_doneIn_0 = x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@48869.4]
  assign RetimeWrapper_3_clock = clock; // @[:@48878.4]
  assign RetimeWrapper_3_reset = reset; // @[:@48879.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@48881.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@48880.4]
  assign RetimeWrapper_4_clock = clock; // @[:@48886.4]
  assign RetimeWrapper_4_reset = reset; // @[:@48887.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@48889.4]
  assign RetimeWrapper_4_io_in = x646_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@48888.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_clock = clock; // @[:@48916.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_reset = reset; // @[:@48917.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TVALID = io_in_x353_TVALID; // @[sm_x646_outr_UnitPipe.scala 48:23:@48972.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TDATA = io_in_x353_TDATA; // @[sm_x646_outr_UnitPipe.scala 48:23:@48970.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TID = io_in_x353_TID; // @[sm_x646_outr_UnitPipe.scala 48:23:@48966.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x353_TDEST = io_in_x353_TDEST; // @[sm_x646_outr_UnitPipe.scala 48:23:@48965.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_in_x354_TREADY = io_in_x354_TREADY; // @[sm_x646_outr_UnitPipe.scala 49:23:@48980.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x646_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x646_outr_UnitPipe.scala 81:22:@48990.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x646_outr_UnitPipe_sm_io_childAck_0; // @[sm_x646_outr_UnitPipe.scala 81:22:@48988.4]
  assign x646_outr_UnitPipe_kernelx646_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x646_outr_UnitPipe.scala 80:18:@48982.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x669_outr_UnitPipe_sm( // @[:@49479.2]
  input   clock, // @[:@49480.4]
  input   reset, // @[:@49481.4]
  input   io_enable, // @[:@49482.4]
  output  io_done, // @[:@49482.4]
  input   io_parentAck, // @[:@49482.4]
  input   io_doneIn_0, // @[:@49482.4]
  input   io_doneIn_1, // @[:@49482.4]
  input   io_doneIn_2, // @[:@49482.4]
  output  io_enableOut_0, // @[:@49482.4]
  output  io_enableOut_1, // @[:@49482.4]
  output  io_enableOut_2, // @[:@49482.4]
  output  io_childAck_0, // @[:@49482.4]
  output  io_childAck_1, // @[:@49482.4]
  output  io_childAck_2, // @[:@49482.4]
  input   io_ctrCopyDone_0, // @[:@49482.4]
  input   io_ctrCopyDone_1, // @[:@49482.4]
  input   io_ctrCopyDone_2 // @[:@49482.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@49485.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@49485.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@49485.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@49485.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@49485.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@49485.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@49488.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@49488.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@49488.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@49488.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@49488.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@49488.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@49491.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@49491.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@49491.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@49491.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@49491.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@49491.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@49494.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@49494.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@49494.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@49494.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@49494.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@49494.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@49497.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@49497.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@49497.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@49497.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@49497.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@49497.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@49500.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@49500.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@49500.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@49500.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@49500.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@49500.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@49541.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@49541.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@49541.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@49541.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@49541.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@49541.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@49544.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@49544.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@49544.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@49544.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@49544.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@49544.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@49547.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@49547.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@49547.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@49547.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@49547.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@49547.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49598.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49598.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49598.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@49598.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@49598.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@49612.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@49612.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@49612.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@49612.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@49612.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@49630.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@49630.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@49630.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@49630.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@49630.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@49667.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@49667.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@49667.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@49667.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@49667.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@49681.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@49681.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@49681.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@49681.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@49681.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@49699.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@49699.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@49699.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@49699.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@49699.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@49736.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@49736.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@49736.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@49736.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@49736.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@49750.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@49750.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@49750.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@49750.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@49750.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@49768.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@49768.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@49768.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@49768.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@49768.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@49825.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@49825.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@49825.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@49825.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@49825.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@49842.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@49842.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@49842.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@49842.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@49842.4]
  wire  _T_77; // @[Controllers.scala 80:47:@49503.4]
  wire  allDone; // @[Controllers.scala 80:47:@49504.4]
  wire  _T_151; // @[Controllers.scala 165:35:@49582.4]
  wire  _T_153; // @[Controllers.scala 165:60:@49583.4]
  wire  _T_154; // @[Controllers.scala 165:58:@49584.4]
  wire  _T_156; // @[Controllers.scala 165:76:@49585.4]
  wire  _T_157; // @[Controllers.scala 165:74:@49586.4]
  wire  _T_161; // @[Controllers.scala 165:109:@49589.4]
  wire  _T_164; // @[Controllers.scala 165:141:@49591.4]
  wire  _T_172; // @[package.scala 96:25:@49603.4 package.scala 96:25:@49604.4]
  wire  _T_176; // @[Controllers.scala 167:54:@49606.4]
  wire  _T_177; // @[Controllers.scala 167:52:@49607.4]
  wire  _T_184; // @[package.scala 96:25:@49617.4 package.scala 96:25:@49618.4]
  wire  _T_202; // @[package.scala 96:25:@49635.4 package.scala 96:25:@49636.4]
  wire  _T_206; // @[Controllers.scala 169:67:@49638.4]
  wire  _T_207; // @[Controllers.scala 169:86:@49639.4]
  wire  _T_219; // @[Controllers.scala 165:35:@49651.4]
  wire  _T_221; // @[Controllers.scala 165:60:@49652.4]
  wire  _T_222; // @[Controllers.scala 165:58:@49653.4]
  wire  _T_224; // @[Controllers.scala 165:76:@49654.4]
  wire  _T_225; // @[Controllers.scala 165:74:@49655.4]
  wire  _T_229; // @[Controllers.scala 165:109:@49658.4]
  wire  _T_232; // @[Controllers.scala 165:141:@49660.4]
  wire  _T_240; // @[package.scala 96:25:@49672.4 package.scala 96:25:@49673.4]
  wire  _T_244; // @[Controllers.scala 167:54:@49675.4]
  wire  _T_245; // @[Controllers.scala 167:52:@49676.4]
  wire  _T_252; // @[package.scala 96:25:@49686.4 package.scala 96:25:@49687.4]
  wire  _T_270; // @[package.scala 96:25:@49704.4 package.scala 96:25:@49705.4]
  wire  _T_274; // @[Controllers.scala 169:67:@49707.4]
  wire  _T_275; // @[Controllers.scala 169:86:@49708.4]
  wire  _T_287; // @[Controllers.scala 165:35:@49720.4]
  wire  _T_289; // @[Controllers.scala 165:60:@49721.4]
  wire  _T_290; // @[Controllers.scala 165:58:@49722.4]
  wire  _T_292; // @[Controllers.scala 165:76:@49723.4]
  wire  _T_293; // @[Controllers.scala 165:74:@49724.4]
  wire  _T_297; // @[Controllers.scala 165:109:@49727.4]
  wire  _T_300; // @[Controllers.scala 165:141:@49729.4]
  wire  _T_308; // @[package.scala 96:25:@49741.4 package.scala 96:25:@49742.4]
  wire  _T_312; // @[Controllers.scala 167:54:@49744.4]
  wire  _T_313; // @[Controllers.scala 167:52:@49745.4]
  wire  _T_320; // @[package.scala 96:25:@49755.4 package.scala 96:25:@49756.4]
  wire  _T_338; // @[package.scala 96:25:@49773.4 package.scala 96:25:@49774.4]
  wire  _T_342; // @[Controllers.scala 169:67:@49776.4]
  wire  _T_343; // @[Controllers.scala 169:86:@49777.4]
  wire  _T_358; // @[Controllers.scala 213:68:@49795.4]
  wire  _T_360; // @[Controllers.scala 213:90:@49797.4]
  wire  _T_362; // @[Controllers.scala 213:132:@49799.4]
  wire  _T_366; // @[Controllers.scala 213:68:@49804.4]
  wire  _T_368; // @[Controllers.scala 213:90:@49806.4]
  wire  _T_374; // @[Controllers.scala 213:68:@49812.4]
  wire  _T_376; // @[Controllers.scala 213:90:@49814.4]
  wire  _T_383; // @[package.scala 100:49:@49820.4]
  reg  _T_386; // @[package.scala 48:56:@49821.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@49823.4]
  reg  _T_400; // @[package.scala 48:56:@49839.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@49485.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@49488.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@49491.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@49494.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@49497.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@49500.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@49541.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@49544.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@49547.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@49598.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@49612.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@49630.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@49667.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@49681.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@49699.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@49736.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@49750.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@49768.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@49825.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@49842.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@49503.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@49504.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@49582.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@49583.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@49584.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@49585.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@49586.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@49589.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@49591.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@49603.4 package.scala 96:25:@49604.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@49606.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@49607.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@49617.4 package.scala 96:25:@49618.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@49635.4 package.scala 96:25:@49636.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@49638.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@49639.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@49651.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@49652.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@49653.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@49654.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@49655.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@49658.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@49660.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@49672.4 package.scala 96:25:@49673.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@49675.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@49676.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@49686.4 package.scala 96:25:@49687.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@49704.4 package.scala 96:25:@49705.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@49707.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@49708.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@49720.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@49721.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@49722.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@49723.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@49724.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@49727.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@49729.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@49741.4 package.scala 96:25:@49742.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@49744.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@49745.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@49755.4 package.scala 96:25:@49756.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@49773.4 package.scala 96:25:@49774.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@49776.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@49777.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@49795.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@49797.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@49799.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@49804.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@49806.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@49812.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@49814.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@49820.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@49823.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@49849.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@49803.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@49811.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@49819.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@49790.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@49792.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@49794.4]
  assign active_0_clock = clock; // @[:@49486.4]
  assign active_0_reset = reset; // @[:@49487.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@49593.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@49597.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@49507.4]
  assign active_1_clock = clock; // @[:@49489.4]
  assign active_1_reset = reset; // @[:@49490.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@49662.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@49666.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@49508.4]
  assign active_2_clock = clock; // @[:@49492.4]
  assign active_2_reset = reset; // @[:@49493.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@49731.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@49735.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@49509.4]
  assign done_0_clock = clock; // @[:@49495.4]
  assign done_0_reset = reset; // @[:@49496.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@49643.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@49521.4 Controllers.scala 170:32:@49650.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@49510.4]
  assign done_1_clock = clock; // @[:@49498.4]
  assign done_1_reset = reset; // @[:@49499.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@49712.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@49530.4 Controllers.scala 170:32:@49719.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@49511.4]
  assign done_2_clock = clock; // @[:@49501.4]
  assign done_2_reset = reset; // @[:@49502.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@49781.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@49539.4 Controllers.scala 170:32:@49788.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@49512.4]
  assign iterDone_0_clock = clock; // @[:@49542.4]
  assign iterDone_0_reset = reset; // @[:@49543.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@49611.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@49561.4 Controllers.scala 168:36:@49627.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@49550.4]
  assign iterDone_1_clock = clock; // @[:@49545.4]
  assign iterDone_1_reset = reset; // @[:@49546.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@49680.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@49570.4 Controllers.scala 168:36:@49696.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@49551.4]
  assign iterDone_2_clock = clock; // @[:@49548.4]
  assign iterDone_2_reset = reset; // @[:@49549.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@49749.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@49579.4 Controllers.scala 168:36:@49765.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@49552.4]
  assign RetimeWrapper_clock = clock; // @[:@49599.4]
  assign RetimeWrapper_reset = reset; // @[:@49600.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@49602.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@49601.4]
  assign RetimeWrapper_1_clock = clock; // @[:@49613.4]
  assign RetimeWrapper_1_reset = reset; // @[:@49614.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@49616.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@49615.4]
  assign RetimeWrapper_2_clock = clock; // @[:@49631.4]
  assign RetimeWrapper_2_reset = reset; // @[:@49632.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@49634.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@49633.4]
  assign RetimeWrapper_3_clock = clock; // @[:@49668.4]
  assign RetimeWrapper_3_reset = reset; // @[:@49669.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@49671.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@49670.4]
  assign RetimeWrapper_4_clock = clock; // @[:@49682.4]
  assign RetimeWrapper_4_reset = reset; // @[:@49683.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@49685.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@49684.4]
  assign RetimeWrapper_5_clock = clock; // @[:@49700.4]
  assign RetimeWrapper_5_reset = reset; // @[:@49701.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@49703.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@49702.4]
  assign RetimeWrapper_6_clock = clock; // @[:@49737.4]
  assign RetimeWrapper_6_reset = reset; // @[:@49738.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@49740.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@49739.4]
  assign RetimeWrapper_7_clock = clock; // @[:@49751.4]
  assign RetimeWrapper_7_reset = reset; // @[:@49752.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@49754.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@49753.4]
  assign RetimeWrapper_8_clock = clock; // @[:@49769.4]
  assign RetimeWrapper_8_reset = reset; // @[:@49770.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@49772.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@49771.4]
  assign RetimeWrapper_9_clock = clock; // @[:@49826.4]
  assign RetimeWrapper_9_reset = reset; // @[:@49827.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@49829.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@49828.4]
  assign RetimeWrapper_10_clock = clock; // @[:@49843.4]
  assign RetimeWrapper_10_reset = reset; // @[:@49844.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@49846.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@49845.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x655_inr_UnitPipe_sm( // @[:@50022.2]
  input   clock, // @[:@50023.4]
  input   reset, // @[:@50024.4]
  input   io_enable, // @[:@50025.4]
  output  io_done, // @[:@50025.4]
  output  io_doneLatch, // @[:@50025.4]
  input   io_ctrDone, // @[:@50025.4]
  output  io_datapathEn, // @[:@50025.4]
  output  io_ctrInc, // @[:@50025.4]
  input   io_parentAck, // @[:@50025.4]
  input   io_backpressure // @[:@50025.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@50027.4]
  wire  active_reset; // @[Controllers.scala 261:22:@50027.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@50027.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@50027.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@50027.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@50027.4]
  wire  done_clock; // @[Controllers.scala 262:20:@50030.4]
  wire  done_reset; // @[Controllers.scala 262:20:@50030.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@50030.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@50030.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@50030.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@50030.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50084.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50084.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50084.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50084.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50084.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50092.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50092.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50092.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50092.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50092.4]
  wire  _T_80; // @[Controllers.scala 264:48:@50035.4]
  wire  _T_81; // @[Controllers.scala 264:46:@50036.4]
  wire  _T_82; // @[Controllers.scala 264:62:@50037.4]
  wire  _T_83; // @[Controllers.scala 264:60:@50038.4]
  wire  _T_100; // @[package.scala 100:49:@50055.4]
  reg  _T_103; // @[package.scala 48:56:@50056.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@50064.4]
  wire  _T_116; // @[Controllers.scala 283:41:@50072.4]
  wire  _T_117; // @[Controllers.scala 283:59:@50073.4]
  wire  _T_119; // @[Controllers.scala 284:37:@50076.4]
  reg  _T_125; // @[package.scala 48:56:@50080.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@50102.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@50105.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@50107.4]
  wire  _T_152; // @[Controllers.scala 292:61:@50108.4]
  wire  _T_153; // @[Controllers.scala 292:24:@50109.4]
  SRFF active ( // @[Controllers.scala 261:22:@50027.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@50030.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50084.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@50092.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@50035.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@50036.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@50037.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@50038.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@50055.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@50064.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@50072.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@50073.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@50076.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@50107.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@50108.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@50109.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@50083.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@50111.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@50075.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@50078.4]
  assign active_clock = clock; // @[:@50028.4]
  assign active_reset = reset; // @[:@50029.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@50040.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@50044.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@50045.4]
  assign done_clock = clock; // @[:@50031.4]
  assign done_reset = reset; // @[:@50032.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@50060.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@50053.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@50054.4]
  assign RetimeWrapper_clock = clock; // @[:@50085.4]
  assign RetimeWrapper_reset = reset; // @[:@50086.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50088.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@50087.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50093.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50094.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@50096.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@50095.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1( // @[:@50186.2]
  output        io_in_x648_valid, // @[:@50189.4]
  output [63:0] io_in_x648_bits_addr, // @[:@50189.4]
  output [31:0] io_in_x648_bits_size, // @[:@50189.4]
  input  [63:0] io_in_x351_outdram_number, // @[:@50189.4]
  input         io_sigsIn_backpressure, // @[:@50189.4]
  input         io_sigsIn_datapathEn, // @[:@50189.4]
  input         io_rr // @[:@50189.4]
);
  wire [96:0] x652_tuple; // @[Cat.scala 30:58:@50203.4]
  wire  _T_135; // @[implicits.scala 55:10:@50206.4]
  assign x652_tuple = {33'h7e9000,io_in_x351_outdram_number}; // @[Cat.scala 30:58:@50203.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@50206.4]
  assign io_in_x648_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x655_inr_UnitPipe.scala 65:18:@50209.4]
  assign io_in_x648_bits_addr = x652_tuple[63:0]; // @[sm_x655_inr_UnitPipe.scala 66:22:@50211.4]
  assign io_in_x648_bits_size = x652_tuple[95:64]; // @[sm_x655_inr_UnitPipe.scala 67:22:@50213.4]
endmodule
module FF_13( // @[:@50215.2]
  input         clock, // @[:@50216.4]
  input         reset, // @[:@50217.4]
  output [22:0] io_rPort_0_output_0, // @[:@50218.4]
  input  [22:0] io_wPort_0_data_0, // @[:@50218.4]
  input         io_wPort_0_reset, // @[:@50218.4]
  input         io_wPort_0_en_0 // @[:@50218.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@50233.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@50235.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@50236.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@50235.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@50236.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@50238.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@50253.2]
  input         clock, // @[:@50254.4]
  input         reset, // @[:@50255.4]
  input         io_input_reset, // @[:@50256.4]
  input         io_input_enable, // @[:@50256.4]
  output [22:0] io_output_count_0, // @[:@50256.4]
  output        io_output_oobs_0, // @[:@50256.4]
  output        io_output_done // @[:@50256.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@50269.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@50269.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@50269.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@50269.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@50269.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@50269.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@50285.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@50285.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@50285.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@50285.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@50285.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@50285.4]
  wire  _T_36; // @[Counter.scala 264:45:@50288.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@50313.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@50314.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@50315.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@50316.4]
  wire  _T_57; // @[Counter.scala 293:18:@50318.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@50326.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@50329.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@50330.4]
  wire  _T_75; // @[Counter.scala 322:102:@50334.4]
  wire  _T_77; // @[Counter.scala 322:130:@50335.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@50269.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@50285.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@50288.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@50313.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@50314.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@50315.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@50316.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@50318.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@50326.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@50329.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@50330.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@50334.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@50335.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@50333.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@50337.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@50339.4]
  assign bases_0_clock = clock; // @[:@50270.4]
  assign bases_0_reset = reset; // @[:@50271.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@50332.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@50311.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@50312.4]
  assign SRFF_clock = clock; // @[:@50286.4]
  assign SRFF_reset = reset; // @[:@50287.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@50290.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@50292.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@50293.4]
endmodule
module x657_ctrchain( // @[:@50344.2]
  input         clock, // @[:@50345.4]
  input         reset, // @[:@50346.4]
  input         io_input_reset, // @[:@50347.4]
  input         io_input_enable, // @[:@50347.4]
  output [22:0] io_output_counts_0, // @[:@50347.4]
  output        io_output_oobs_0, // @[:@50347.4]
  output        io_output_done // @[:@50347.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@50349.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@50349.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@50349.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@50349.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@50349.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@50349.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@50349.4]
  reg  wasDone; // @[Counter.scala 542:24:@50358.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@50364.4]
  wire  _T_47; // @[Counter.scala 546:80:@50365.4]
  reg  doneLatch; // @[Counter.scala 550:26:@50370.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@50371.4]
  wire  _T_55; // @[Counter.scala 551:19:@50372.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@50349.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@50364.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@50365.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@50371.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@50372.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@50374.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@50376.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@50367.4]
  assign ctrs_0_clock = clock; // @[:@50350.4]
  assign ctrs_0_reset = reset; // @[:@50351.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@50355.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@50356.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x664_inr_Foreach_sm( // @[:@50564.2]
  input   clock, // @[:@50565.4]
  input   reset, // @[:@50566.4]
  input   io_enable, // @[:@50567.4]
  output  io_done, // @[:@50567.4]
  output  io_doneLatch, // @[:@50567.4]
  input   io_ctrDone, // @[:@50567.4]
  output  io_datapathEn, // @[:@50567.4]
  output  io_ctrInc, // @[:@50567.4]
  output  io_ctrRst, // @[:@50567.4]
  input   io_parentAck, // @[:@50567.4]
  input   io_backpressure, // @[:@50567.4]
  input   io_break // @[:@50567.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@50569.4]
  wire  active_reset; // @[Controllers.scala 261:22:@50569.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@50569.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@50569.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@50569.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@50569.4]
  wire  done_clock; // @[Controllers.scala 262:20:@50572.4]
  wire  done_reset; // @[Controllers.scala 262:20:@50572.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@50572.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@50572.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@50572.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@50572.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50606.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50606.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50606.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50606.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50606.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50628.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50628.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50628.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50628.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50628.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@50640.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@50640.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@50640.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@50640.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@50640.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@50648.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@50648.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@50648.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@50648.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@50648.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@50664.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@50664.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@50664.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@50664.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@50664.4]
  wire  _T_80; // @[Controllers.scala 264:48:@50577.4]
  wire  _T_81; // @[Controllers.scala 264:46:@50578.4]
  wire  _T_82; // @[Controllers.scala 264:62:@50579.4]
  wire  _T_83; // @[Controllers.scala 264:60:@50580.4]
  wire  _T_100; // @[package.scala 100:49:@50597.4]
  reg  _T_103; // @[package.scala 48:56:@50598.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@50611.4 package.scala 96:25:@50612.4]
  wire  _T_110; // @[package.scala 100:49:@50613.4]
  reg  _T_113; // @[package.scala 48:56:@50614.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@50616.4]
  wire  _T_118; // @[Controllers.scala 283:41:@50621.4]
  wire  _T_119; // @[Controllers.scala 283:59:@50622.4]
  wire  _T_121; // @[Controllers.scala 284:37:@50625.4]
  wire  _T_124; // @[package.scala 96:25:@50633.4 package.scala 96:25:@50634.4]
  wire  _T_126; // @[package.scala 100:49:@50635.4]
  reg  _T_129; // @[package.scala 48:56:@50636.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@50658.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@50660.4]
  reg  _T_153; // @[package.scala 48:56:@50661.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@50669.4 package.scala 96:25:@50670.4]
  wire  _T_158; // @[Controllers.scala 292:61:@50671.4]
  wire  _T_159; // @[Controllers.scala 292:24:@50672.4]
  SRFF active ( // @[Controllers.scala 261:22:@50569.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@50572.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@50606.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@50628.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@50640.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@50648.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@50664.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@50577.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@50578.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@50579.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@50580.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@50597.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@50611.4 package.scala 96:25:@50612.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@50613.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@50616.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@50621.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@50622.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@50625.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@50633.4 package.scala 96:25:@50634.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@50635.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@50660.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@50669.4 package.scala 96:25:@50670.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@50671.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@50672.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@50639.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@50674.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@50624.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@50627.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@50619.4]
  assign active_clock = clock; // @[:@50570.4]
  assign active_reset = reset; // @[:@50571.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@50582.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@50586.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@50587.4]
  assign done_clock = clock; // @[:@50573.4]
  assign done_reset = reset; // @[:@50574.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@50602.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@50595.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@50596.4]
  assign RetimeWrapper_clock = clock; // @[:@50607.4]
  assign RetimeWrapper_reset = reset; // @[:@50608.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@50610.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@50609.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50629.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50630.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@50632.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@50631.4]
  assign RetimeWrapper_2_clock = clock; // @[:@50641.4]
  assign RetimeWrapper_2_reset = reset; // @[:@50642.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@50644.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@50643.4]
  assign RetimeWrapper_3_clock = clock; // @[:@50649.4]
  assign RetimeWrapper_3_reset = reset; // @[:@50650.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@50652.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@50651.4]
  assign RetimeWrapper_4_clock = clock; // @[:@50665.4]
  assign RetimeWrapper_4_reset = reset; // @[:@50666.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@50668.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@50667.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x664_inr_Foreach_kernelx664_inr_Foreach_concrete1( // @[:@50881.2]
  input         clock, // @[:@50882.4]
  input         reset, // @[:@50883.4]
  output        io_in_x649_valid, // @[:@50884.4]
  output [31:0] io_in_x649_bits_wdata_0, // @[:@50884.4]
  output        io_in_x649_bits_wstrb, // @[:@50884.4]
  output [20:0] io_in_x355_outbuf_0_rPort_0_ofs_0, // @[:@50884.4]
  output        io_in_x355_outbuf_0_rPort_0_en_0, // @[:@50884.4]
  output        io_in_x355_outbuf_0_rPort_0_backpressure, // @[:@50884.4]
  input  [31:0] io_in_x355_outbuf_0_rPort_0_output_0, // @[:@50884.4]
  input         io_sigsIn_backpressure, // @[:@50884.4]
  input         io_sigsIn_datapathEn, // @[:@50884.4]
  input         io_sigsIn_break, // @[:@50884.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@50884.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@50884.4]
  input         io_rr // @[:@50884.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@50911.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@50911.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50940.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50940.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50940.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50940.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50940.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50949.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50949.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50949.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50949.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50949.4]
  wire  b659; // @[sm_x664_inr_Foreach.scala 62:18:@50919.4]
  wire  _T_274; // @[sm_x664_inr_Foreach.scala 67:129:@50923.4]
  wire  _T_278; // @[implicits.scala 55:10:@50926.4]
  wire  _T_279; // @[sm_x664_inr_Foreach.scala 67:146:@50927.4]
  wire [32:0] x662_tuple; // @[Cat.scala 30:58:@50937.4]
  wire  _T_290; // @[package.scala 96:25:@50954.4 package.scala 96:25:@50955.4]
  wire  _T_292; // @[implicits.scala 55:10:@50956.4]
  wire  x816_b659_D2; // @[package.scala 96:25:@50945.4 package.scala 96:25:@50946.4]
  wire  _T_293; // @[sm_x664_inr_Foreach.scala 74:112:@50957.4]
  wire [31:0] b658_number; // @[Math.scala 723:22:@50916.4 Math.scala 724:14:@50917.4]
  _ _ ( // @[Math.scala 720:24:@50911.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@50940.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@50949.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b659 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x664_inr_Foreach.scala 62:18:@50919.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x664_inr_Foreach.scala 67:129:@50923.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@50926.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x664_inr_Foreach.scala 67:146:@50927.4]
  assign x662_tuple = {1'h1,io_in_x355_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@50937.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@50954.4 package.scala 96:25:@50955.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@50956.4]
  assign x816_b659_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@50945.4 package.scala 96:25:@50946.4]
  assign _T_293 = _T_292 & x816_b659_D2; // @[sm_x664_inr_Foreach.scala 74:112:@50957.4]
  assign b658_number = __io_result; // @[Math.scala 723:22:@50916.4 Math.scala 724:14:@50917.4]
  assign io_in_x649_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x664_inr_Foreach.scala 74:18:@50959.4]
  assign io_in_x649_bits_wdata_0 = x662_tuple[31:0]; // @[sm_x664_inr_Foreach.scala 75:26:@50961.4]
  assign io_in_x649_bits_wstrb = x662_tuple[32]; // @[sm_x664_inr_Foreach.scala 76:23:@50963.4]
  assign io_in_x355_outbuf_0_rPort_0_ofs_0 = b658_number[20:0]; // @[MemInterfaceType.scala 107:54:@50930.4]
  assign io_in_x355_outbuf_0_rPort_0_en_0 = _T_279 & b659; // @[MemInterfaceType.scala 110:79:@50932.4]
  assign io_in_x355_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@50931.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@50914.4]
  assign RetimeWrapper_clock = clock; // @[:@50941.4]
  assign RetimeWrapper_reset = reset; // @[:@50942.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@50944.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@50943.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50950.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50951.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@50953.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@50952.4]
endmodule
module x668_inr_UnitPipe_sm( // @[:@51119.2]
  input   clock, // @[:@51120.4]
  input   reset, // @[:@51121.4]
  input   io_enable, // @[:@51122.4]
  output  io_done, // @[:@51122.4]
  output  io_doneLatch, // @[:@51122.4]
  input   io_ctrDone, // @[:@51122.4]
  output  io_datapathEn, // @[:@51122.4]
  output  io_ctrInc, // @[:@51122.4]
  input   io_parentAck // @[:@51122.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@51124.4]
  wire  active_reset; // @[Controllers.scala 261:22:@51124.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@51124.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@51124.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@51124.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@51124.4]
  wire  done_clock; // @[Controllers.scala 262:20:@51127.4]
  wire  done_reset; // @[Controllers.scala 262:20:@51127.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@51127.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@51127.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@51127.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@51127.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@51161.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@51161.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@51161.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@51161.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@51161.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@51183.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@51183.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@51183.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@51183.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@51183.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@51195.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@51195.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@51195.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@51195.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@51195.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@51203.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@51203.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@51203.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@51203.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@51203.4]
  wire  _T_80; // @[Controllers.scala 264:48:@51132.4]
  wire  _T_81; // @[Controllers.scala 264:46:@51133.4]
  wire  _T_82; // @[Controllers.scala 264:62:@51134.4]
  wire  _T_100; // @[package.scala 100:49:@51152.4]
  reg  _T_103; // @[package.scala 48:56:@51153.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@51176.4]
  wire  _T_124; // @[package.scala 96:25:@51188.4 package.scala 96:25:@51189.4]
  wire  _T_126; // @[package.scala 100:49:@51190.4]
  reg  _T_129; // @[package.scala 48:56:@51191.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@51213.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@51215.4]
  reg  _T_153; // @[package.scala 48:56:@51216.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@51218.4]
  wire  _T_156; // @[Controllers.scala 292:61:@51219.4]
  wire  _T_157; // @[Controllers.scala 292:24:@51220.4]
  SRFF active ( // @[Controllers.scala 261:22:@51124.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@51127.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@51161.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@51183.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@51195.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@51203.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@51132.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@51133.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@51134.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@51152.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@51176.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@51188.4 package.scala 96:25:@51189.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@51190.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@51215.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@51218.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@51219.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@51220.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@51194.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@51222.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@51179.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@51182.4]
  assign active_clock = clock; // @[:@51125.4]
  assign active_reset = reset; // @[:@51126.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@51137.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@51141.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@51142.4]
  assign done_clock = clock; // @[:@51128.4]
  assign done_reset = reset; // @[:@51129.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@51157.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@51150.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@51151.4]
  assign RetimeWrapper_clock = clock; // @[:@51162.4]
  assign RetimeWrapper_reset = reset; // @[:@51163.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@51165.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@51164.4]
  assign RetimeWrapper_1_clock = clock; // @[:@51184.4]
  assign RetimeWrapper_1_reset = reset; // @[:@51185.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@51187.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@51186.4]
  assign RetimeWrapper_2_clock = clock; // @[:@51196.4]
  assign RetimeWrapper_2_reset = reset; // @[:@51197.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@51199.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@51198.4]
  assign RetimeWrapper_3_clock = clock; // @[:@51204.4]
  assign RetimeWrapper_3_reset = reset; // @[:@51205.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@51207.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@51206.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1( // @[:@51297.2]
  output  io_in_x650_ready, // @[:@51300.4]
  input   io_sigsIn_datapathEn // @[:@51300.4]
);
  assign io_in_x650_ready = io_sigsIn_datapathEn; // @[sm_x668_inr_UnitPipe.scala 57:18:@51312.4]
endmodule
module x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1( // @[:@51315.2]
  input         clock, // @[:@51316.4]
  input         reset, // @[:@51317.4]
  output        io_in_x650_ready, // @[:@51318.4]
  input         io_in_x650_valid, // @[:@51318.4]
  input         io_in_x649_ready, // @[:@51318.4]
  output        io_in_x649_valid, // @[:@51318.4]
  output [31:0] io_in_x649_bits_wdata_0, // @[:@51318.4]
  output        io_in_x649_bits_wstrb, // @[:@51318.4]
  input         io_in_x648_ready, // @[:@51318.4]
  output        io_in_x648_valid, // @[:@51318.4]
  output [63:0] io_in_x648_bits_addr, // @[:@51318.4]
  output [31:0] io_in_x648_bits_size, // @[:@51318.4]
  output [20:0] io_in_x355_outbuf_0_rPort_0_ofs_0, // @[:@51318.4]
  output        io_in_x355_outbuf_0_rPort_0_en_0, // @[:@51318.4]
  output        io_in_x355_outbuf_0_rPort_0_backpressure, // @[:@51318.4]
  input  [31:0] io_in_x355_outbuf_0_rPort_0_output_0, // @[:@51318.4]
  input  [63:0] io_in_x351_outdram_number, // @[:@51318.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@51318.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@51318.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@51318.4]
  input         io_sigsIn_smChildAcks_0, // @[:@51318.4]
  input         io_sigsIn_smChildAcks_1, // @[:@51318.4]
  input         io_sigsIn_smChildAcks_2, // @[:@51318.4]
  output        io_sigsOut_smDoneIn_0, // @[:@51318.4]
  output        io_sigsOut_smDoneIn_1, // @[:@51318.4]
  output        io_sigsOut_smDoneIn_2, // @[:@51318.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@51318.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@51318.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@51318.4]
  input         io_rr // @[:@51318.4]
);
  wire  x655_inr_UnitPipe_sm_clock; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_reset; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_enable; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_done; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_doneLatch; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_ctrDone; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_datapathEn; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_ctrInc; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_parentAck; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  x655_inr_UnitPipe_sm_io_backpressure; // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@51442.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@51442.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@51442.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@51442.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@51442.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@51450.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@51450.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@51450.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@51450.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@51450.4]
  wire  x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_valid; // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
  wire [63:0] x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_bits_addr; // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
  wire [31:0] x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_bits_size; // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
  wire [63:0] x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x351_outdram_number; // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
  wire  x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
  wire  x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
  wire  x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_rr; // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
  wire  x657_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@51548.4]
  wire  x657_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@51548.4]
  wire  x657_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@51548.4]
  wire  x657_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@51548.4]
  wire [22:0] x657_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@51548.4]
  wire  x657_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@51548.4]
  wire  x657_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@51548.4]
  wire  x664_inr_Foreach_sm_clock; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_reset; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_enable; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_done; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_doneLatch; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_ctrDone; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_datapathEn; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_ctrInc; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_ctrRst; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_parentAck; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_backpressure; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  x664_inr_Foreach_sm_io_break; // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@51629.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@51629.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@51629.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@51629.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@51629.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@51669.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@51669.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@51669.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@51669.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@51669.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@51677.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@51677.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@51677.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@51677.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@51677.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_clock; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_reset; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_valid; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire [31:0] x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_bits_wdata_0; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_bits_wstrb; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire [20:0] x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_en_0; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire [31:0] x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_output_0; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire [31:0] x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_rr; // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
  wire  x668_inr_UnitPipe_sm_clock; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_reset; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_io_enable; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_io_done; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_io_doneLatch; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_io_ctrDone; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_io_datapathEn; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_io_ctrInc; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  x668_inr_UnitPipe_sm_io_parentAck; // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@51889.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@51889.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@51889.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@51889.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@51889.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@51897.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@51897.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@51897.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@51897.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@51897.4]
  wire  x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1_io_in_x650_ready; // @[sm_x668_inr_UnitPipe.scala 60:24:@51927.4]
  wire  x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x668_inr_UnitPipe.scala 60:24:@51927.4]
  wire  _T_359; // @[package.scala 100:49:@51413.4]
  reg  _T_362; // @[package.scala 48:56:@51414.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@51447.4 package.scala 96:25:@51448.4]
  wire  _T_381; // @[package.scala 96:25:@51455.4 package.scala 96:25:@51456.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@51458.4]
  wire  _T_454; // @[package.scala 96:25:@51634.4 package.scala 96:25:@51635.4]
  wire  _T_468; // @[package.scala 96:25:@51674.4 package.scala 96:25:@51675.4]
  wire  _T_474; // @[package.scala 96:25:@51682.4 package.scala 96:25:@51683.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@51685.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@51694.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@51695.4]
  wire  _T_547; // @[package.scala 100:49:@51860.4]
  reg  _T_550; // @[package.scala 48:56:@51861.4]
  reg [31:0] _RAND_1;
  wire  x668_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x669_outr_UnitPipe.scala 101:55:@51867.4]
  wire  _T_563; // @[package.scala 96:25:@51894.4 package.scala 96:25:@51895.4]
  wire  _T_569; // @[package.scala 96:25:@51902.4 package.scala 96:25:@51903.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@51905.4]
  wire  x668_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@51906.4]
  x655_inr_UnitPipe_sm x655_inr_UnitPipe_sm ( // @[sm_x655_inr_UnitPipe.scala 33:18:@51385.4]
    .clock(x655_inr_UnitPipe_sm_clock),
    .reset(x655_inr_UnitPipe_sm_reset),
    .io_enable(x655_inr_UnitPipe_sm_io_enable),
    .io_done(x655_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x655_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x655_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x655_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x655_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x655_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x655_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@51442.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@51450.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1 x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1 ( // @[sm_x655_inr_UnitPipe.scala 69:24:@51480.4]
    .io_in_x648_valid(x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_valid),
    .io_in_x648_bits_addr(x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_bits_addr),
    .io_in_x648_bits_size(x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_bits_size),
    .io_in_x351_outdram_number(x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x351_outdram_number),
    .io_sigsIn_backpressure(x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_rr)
  );
  x657_ctrchain x657_ctrchain ( // @[SpatialBlocks.scala 37:22:@51548.4]
    .clock(x657_ctrchain_clock),
    .reset(x657_ctrchain_reset),
    .io_input_reset(x657_ctrchain_io_input_reset),
    .io_input_enable(x657_ctrchain_io_input_enable),
    .io_output_counts_0(x657_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x657_ctrchain_io_output_oobs_0),
    .io_output_done(x657_ctrchain_io_output_done)
  );
  x664_inr_Foreach_sm x664_inr_Foreach_sm ( // @[sm_x664_inr_Foreach.scala 33:18:@51601.4]
    .clock(x664_inr_Foreach_sm_clock),
    .reset(x664_inr_Foreach_sm_reset),
    .io_enable(x664_inr_Foreach_sm_io_enable),
    .io_done(x664_inr_Foreach_sm_io_done),
    .io_doneLatch(x664_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x664_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x664_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x664_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x664_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x664_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x664_inr_Foreach_sm_io_backpressure),
    .io_break(x664_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@51629.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@51669.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@51677.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x664_inr_Foreach_kernelx664_inr_Foreach_concrete1 x664_inr_Foreach_kernelx664_inr_Foreach_concrete1 ( // @[sm_x664_inr_Foreach.scala 78:24:@51712.4]
    .clock(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_clock),
    .reset(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_reset),
    .io_in_x649_valid(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_valid),
    .io_in_x649_bits_wdata_0(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_bits_wdata_0),
    .io_in_x649_bits_wstrb(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_bits_wstrb),
    .io_in_x355_outbuf_0_rPort_0_ofs_0(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0),
    .io_in_x355_outbuf_0_rPort_0_en_0(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_en_0),
    .io_in_x355_outbuf_0_rPort_0_backpressure(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure),
    .io_in_x355_outbuf_0_rPort_0_output_0(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_output_0),
    .io_sigsIn_backpressure(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_rr)
  );
  x668_inr_UnitPipe_sm x668_inr_UnitPipe_sm ( // @[sm_x668_inr_UnitPipe.scala 32:18:@51832.4]
    .clock(x668_inr_UnitPipe_sm_clock),
    .reset(x668_inr_UnitPipe_sm_reset),
    .io_enable(x668_inr_UnitPipe_sm_io_enable),
    .io_done(x668_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x668_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x668_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x668_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x668_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x668_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@51889.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@51897.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1 x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1 ( // @[sm_x668_inr_UnitPipe.scala 60:24:@51927.4]
    .io_in_x650_ready(x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1_io_in_x650_ready),
    .io_sigsIn_datapathEn(x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x655_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@51413.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@51447.4 package.scala 96:25:@51448.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@51455.4 package.scala 96:25:@51456.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@51458.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@51634.4 package.scala 96:25:@51635.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@51674.4 package.scala 96:25:@51675.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@51682.4 package.scala 96:25:@51683.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@51685.4]
  assign _T_479 = x664_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@51694.4]
  assign _T_480 = ~ x664_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@51695.4]
  assign _T_547 = x668_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@51860.4]
  assign x668_inr_UnitPipe_sigsIn_forwardpressure = io_in_x650_valid | x668_inr_UnitPipe_sm_io_doneLatch; // @[sm_x669_outr_UnitPipe.scala 101:55:@51867.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@51894.4 package.scala 96:25:@51895.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@51902.4 package.scala 96:25:@51903.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@51905.4]
  assign x668_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@51906.4]
  assign io_in_x650_ready = x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1_io_in_x650_ready; // @[sm_x668_inr_UnitPipe.scala 46:23:@51963.4]
  assign io_in_x649_valid = x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_valid; // @[sm_x664_inr_Foreach.scala 49:23:@51762.4]
  assign io_in_x649_bits_wdata_0 = x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_bits_wdata_0; // @[sm_x664_inr_Foreach.scala 49:23:@51761.4]
  assign io_in_x649_bits_wstrb = x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x649_bits_wstrb; // @[sm_x664_inr_Foreach.scala 49:23:@51760.4]
  assign io_in_x648_valid = x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_valid; // @[sm_x655_inr_UnitPipe.scala 49:23:@51518.4]
  assign io_in_x648_bits_addr = x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_bits_addr; // @[sm_x655_inr_UnitPipe.scala 49:23:@51517.4]
  assign io_in_x648_bits_size = x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x648_bits_size; // @[sm_x655_inr_UnitPipe.scala 49:23:@51516.4]
  assign io_in_x355_outbuf_0_rPort_0_ofs_0 = x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@51767.4]
  assign io_in_x355_outbuf_0_rPort_0_en_0 = x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@51766.4]
  assign io_in_x355_outbuf_0_rPort_0_backpressure = x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@51765.4]
  assign io_sigsOut_smDoneIn_0 = x655_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@51465.4]
  assign io_sigsOut_smDoneIn_1 = x664_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@51692.4]
  assign io_sigsOut_smDoneIn_2 = x668_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@51912.4]
  assign io_sigsOut_smCtrCopyDone_0 = x655_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@51479.4]
  assign io_sigsOut_smCtrCopyDone_1 = x664_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@51711.4]
  assign io_sigsOut_smCtrCopyDone_2 = x668_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@51926.4]
  assign x655_inr_UnitPipe_sm_clock = clock; // @[:@51386.4]
  assign x655_inr_UnitPipe_sm_reset = reset; // @[:@51387.4]
  assign x655_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@51462.4]
  assign x655_inr_UnitPipe_sm_io_ctrDone = x655_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x669_outr_UnitPipe.scala 77:39:@51417.4]
  assign x655_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@51464.4]
  assign x655_inr_UnitPipe_sm_io_backpressure = io_in_x648_ready | x655_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@51436.4]
  assign RetimeWrapper_clock = clock; // @[:@51443.4]
  assign RetimeWrapper_reset = reset; // @[:@51444.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@51446.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@51445.4]
  assign RetimeWrapper_1_clock = clock; // @[:@51451.4]
  assign RetimeWrapper_1_reset = reset; // @[:@51452.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@51454.4]
  assign RetimeWrapper_1_io_in = x655_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@51453.4]
  assign x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_in_x351_outdram_number = io_in_x351_outdram_number; // @[sm_x655_inr_UnitPipe.scala 50:31:@51520.4]
  assign x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x648_ready | x655_inr_UnitPipe_sm_io_doneLatch; // @[sm_x655_inr_UnitPipe.scala 74:22:@51535.4]
  assign x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x655_inr_UnitPipe_sm_io_datapathEn; // @[sm_x655_inr_UnitPipe.scala 74:22:@51533.4]
  assign x655_inr_UnitPipe_kernelx655_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x655_inr_UnitPipe.scala 73:18:@51521.4]
  assign x657_ctrchain_clock = clock; // @[:@51549.4]
  assign x657_ctrchain_reset = reset; // @[:@51550.4]
  assign x657_ctrchain_io_input_reset = x664_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@51710.4]
  assign x657_ctrchain_io_input_enable = x664_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@51662.4 SpatialBlocks.scala 159:42:@51709.4]
  assign x664_inr_Foreach_sm_clock = clock; // @[:@51602.4]
  assign x664_inr_Foreach_sm_reset = reset; // @[:@51603.4]
  assign x664_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@51689.4]
  assign x664_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x669_outr_UnitPipe.scala 90:38:@51637.4]
  assign x664_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@51691.4]
  assign x664_inr_Foreach_sm_io_backpressure = io_in_x649_ready | x664_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@51663.4]
  assign x664_inr_Foreach_sm_io_break = 1'h0; // @[sm_x669_outr_UnitPipe.scala 94:36:@51643.4]
  assign RetimeWrapper_2_clock = clock; // @[:@51630.4]
  assign RetimeWrapper_2_reset = reset; // @[:@51631.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@51633.4]
  assign RetimeWrapper_2_io_in = x657_ctrchain_io_output_done; // @[package.scala 94:16:@51632.4]
  assign RetimeWrapper_3_clock = clock; // @[:@51670.4]
  assign RetimeWrapper_3_reset = reset; // @[:@51671.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@51673.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@51672.4]
  assign RetimeWrapper_4_clock = clock; // @[:@51678.4]
  assign RetimeWrapper_4_reset = reset; // @[:@51679.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@51681.4]
  assign RetimeWrapper_4_io_in = x664_inr_Foreach_sm_io_done; // @[package.scala 94:16:@51680.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_clock = clock; // @[:@51713.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_reset = reset; // @[:@51714.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_in_x355_outbuf_0_rPort_0_output_0 = io_in_x355_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@51764.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x649_ready | x664_inr_Foreach_sm_io_doneLatch; // @[sm_x664_inr_Foreach.scala 83:22:@51783.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x664_inr_Foreach.scala 83:22:@51781.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_break = x664_inr_Foreach_sm_io_break; // @[sm_x664_inr_Foreach.scala 83:22:@51779.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x657_ctrchain_io_output_counts_0[22]}},x657_ctrchain_io_output_counts_0}; // @[sm_x664_inr_Foreach.scala 83:22:@51774.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x657_ctrchain_io_output_oobs_0; // @[sm_x664_inr_Foreach.scala 83:22:@51773.4]
  assign x664_inr_Foreach_kernelx664_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x664_inr_Foreach.scala 82:18:@51769.4]
  assign x668_inr_UnitPipe_sm_clock = clock; // @[:@51833.4]
  assign x668_inr_UnitPipe_sm_reset = reset; // @[:@51834.4]
  assign x668_inr_UnitPipe_sm_io_enable = x668_inr_UnitPipe_sigsIn_baseEn & x668_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@51909.4]
  assign x668_inr_UnitPipe_sm_io_ctrDone = x668_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x669_outr_UnitPipe.scala 99:39:@51864.4]
  assign x668_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@51911.4]
  assign RetimeWrapper_5_clock = clock; // @[:@51890.4]
  assign RetimeWrapper_5_reset = reset; // @[:@51891.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@51893.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@51892.4]
  assign RetimeWrapper_6_clock = clock; // @[:@51898.4]
  assign RetimeWrapper_6_reset = reset; // @[:@51899.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@51901.4]
  assign RetimeWrapper_6_io_in = x668_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@51900.4]
  assign x668_inr_UnitPipe_kernelx668_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x668_inr_UnitPipe_sm_io_datapathEn; // @[sm_x668_inr_UnitPipe.scala 65:22:@51976.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x724_kernelx724_concrete1( // @[:@51992.2]
  input          clock, // @[:@51993.4]
  input          reset, // @[:@51994.4]
  input          io_in_x353_TVALID, // @[:@51995.4]
  output         io_in_x353_TREADY, // @[:@51995.4]
  input  [255:0] io_in_x353_TDATA, // @[:@51995.4]
  input  [7:0]   io_in_x353_TID, // @[:@51995.4]
  input  [7:0]   io_in_x353_TDEST, // @[:@51995.4]
  output         io_in_x650_ready, // @[:@51995.4]
  input          io_in_x650_valid, // @[:@51995.4]
  input          io_in_x649_ready, // @[:@51995.4]
  output         io_in_x649_valid, // @[:@51995.4]
  output [31:0]  io_in_x649_bits_wdata_0, // @[:@51995.4]
  output         io_in_x649_bits_wstrb, // @[:@51995.4]
  input          io_in_x648_ready, // @[:@51995.4]
  output         io_in_x648_valid, // @[:@51995.4]
  output [63:0]  io_in_x648_bits_addr, // @[:@51995.4]
  output [31:0]  io_in_x648_bits_size, // @[:@51995.4]
  output [20:0]  io_in_x355_outbuf_0_rPort_0_ofs_0, // @[:@51995.4]
  output         io_in_x355_outbuf_0_rPort_0_en_0, // @[:@51995.4]
  output         io_in_x355_outbuf_0_rPort_0_backpressure, // @[:@51995.4]
  input  [31:0]  io_in_x355_outbuf_0_rPort_0_output_0, // @[:@51995.4]
  input  [63:0]  io_in_x351_outdram_number, // @[:@51995.4]
  output         io_in_x354_TVALID, // @[:@51995.4]
  input          io_in_x354_TREADY, // @[:@51995.4]
  output [255:0] io_in_x354_TDATA, // @[:@51995.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@51995.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@51995.4]
  input          io_sigsIn_smChildAcks_0, // @[:@51995.4]
  input          io_sigsIn_smChildAcks_1, // @[:@51995.4]
  output         io_sigsOut_smDoneIn_0, // @[:@51995.4]
  output         io_sigsOut_smDoneIn_1, // @[:@51995.4]
  input          io_rr // @[:@51995.4]
);
  wire  x647_outr_UnitPipe_sm_clock; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_reset; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_enable; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_done; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_parentAck; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_childAck_0; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_childAck_1; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  x647_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@52130.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@52130.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@52130.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@52130.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@52130.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@52138.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@52138.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@52138.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@52138.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@52138.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_clock; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_reset; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TVALID; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TREADY; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire [255:0] x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TDATA; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire [7:0] x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TID; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire [7:0] x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TDEST; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TVALID; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TREADY; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire [255:0] x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TDATA; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_rr; // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
  wire  x669_outr_UnitPipe_sm_clock; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_reset; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_enable; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_done; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_parentAck; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_childAck_0; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_childAck_1; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_childAck_2; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  x669_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@52419.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@52419.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@52419.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@52419.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@52419.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@52427.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@52427.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@52427.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@52427.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@52427.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_clock; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_reset; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x650_ready; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x650_valid; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_ready; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_valid; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire [31:0] x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_bits_wdata_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_bits_wstrb; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_ready; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_valid; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire [63:0] x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_bits_addr; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire [31:0] x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_bits_size; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire [20:0] x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_en_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire [31:0] x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_output_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire [63:0] x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x351_outdram_number; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_rr; // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
  wire  _T_408; // @[package.scala 96:25:@52135.4 package.scala 96:25:@52136.4]
  wire  _T_414; // @[package.scala 96:25:@52143.4 package.scala 96:25:@52144.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@52146.4]
  wire  _T_508; // @[package.scala 96:25:@52424.4 package.scala 96:25:@52425.4]
  wire  _T_514; // @[package.scala 96:25:@52432.4 package.scala 96:25:@52433.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@52435.4]
  x647_outr_UnitPipe_sm x647_outr_UnitPipe_sm ( // @[sm_x647_outr_UnitPipe.scala 32:18:@52068.4]
    .clock(x647_outr_UnitPipe_sm_clock),
    .reset(x647_outr_UnitPipe_sm_reset),
    .io_enable(x647_outr_UnitPipe_sm_io_enable),
    .io_done(x647_outr_UnitPipe_sm_io_done),
    .io_parentAck(x647_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x647_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x647_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x647_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x647_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x647_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x647_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x647_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x647_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@52130.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@52138.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1 x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1 ( // @[sm_x647_outr_UnitPipe.scala 87:24:@52169.4]
    .clock(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_clock),
    .reset(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_reset),
    .io_in_x353_TVALID(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TVALID),
    .io_in_x353_TREADY(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TREADY),
    .io_in_x353_TDATA(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TDATA),
    .io_in_x353_TID(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TID),
    .io_in_x353_TDEST(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TDEST),
    .io_in_x354_TVALID(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TVALID),
    .io_in_x354_TREADY(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TREADY),
    .io_in_x354_TDATA(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TDATA),
    .io_sigsIn_smEnableOuts_0(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_rr)
  );
  x669_outr_UnitPipe_sm x669_outr_UnitPipe_sm ( // @[sm_x669_outr_UnitPipe.scala 36:18:@52347.4]
    .clock(x669_outr_UnitPipe_sm_clock),
    .reset(x669_outr_UnitPipe_sm_reset),
    .io_enable(x669_outr_UnitPipe_sm_io_enable),
    .io_done(x669_outr_UnitPipe_sm_io_done),
    .io_parentAck(x669_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x669_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x669_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x669_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x669_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x669_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x669_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x669_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x669_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x669_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x669_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x669_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x669_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@52419.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@52427.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1 x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1 ( // @[sm_x669_outr_UnitPipe.scala 108:24:@52459.4]
    .clock(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_clock),
    .reset(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_reset),
    .io_in_x650_ready(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x650_ready),
    .io_in_x650_valid(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x650_valid),
    .io_in_x649_ready(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_ready),
    .io_in_x649_valid(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_valid),
    .io_in_x649_bits_wdata_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_bits_wdata_0),
    .io_in_x649_bits_wstrb(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_bits_wstrb),
    .io_in_x648_ready(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_ready),
    .io_in_x648_valid(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_valid),
    .io_in_x648_bits_addr(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_bits_addr),
    .io_in_x648_bits_size(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_bits_size),
    .io_in_x355_outbuf_0_rPort_0_ofs_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0),
    .io_in_x355_outbuf_0_rPort_0_en_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_en_0),
    .io_in_x355_outbuf_0_rPort_0_backpressure(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure),
    .io_in_x355_outbuf_0_rPort_0_output_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_output_0),
    .io_in_x351_outdram_number(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x351_outdram_number),
    .io_sigsIn_smEnableOuts_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@52135.4 package.scala 96:25:@52136.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@52143.4 package.scala 96:25:@52144.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@52146.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@52424.4 package.scala 96:25:@52425.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@52432.4 package.scala 96:25:@52433.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@52435.4]
  assign io_in_x353_TREADY = x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TREADY; // @[sm_x647_outr_UnitPipe.scala 48:23:@52237.4]
  assign io_in_x650_ready = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x650_ready; // @[sm_x669_outr_UnitPipe.scala 58:23:@52541.4]
  assign io_in_x649_valid = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_valid; // @[sm_x669_outr_UnitPipe.scala 59:23:@52544.4]
  assign io_in_x649_bits_wdata_0 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_bits_wdata_0; // @[sm_x669_outr_UnitPipe.scala 59:23:@52543.4]
  assign io_in_x649_bits_wstrb = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_bits_wstrb; // @[sm_x669_outr_UnitPipe.scala 59:23:@52542.4]
  assign io_in_x648_valid = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_valid; // @[sm_x669_outr_UnitPipe.scala 60:23:@52548.4]
  assign io_in_x648_bits_addr = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_bits_addr; // @[sm_x669_outr_UnitPipe.scala 60:23:@52547.4]
  assign io_in_x648_bits_size = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_bits_size; // @[sm_x669_outr_UnitPipe.scala 60:23:@52546.4]
  assign io_in_x355_outbuf_0_rPort_0_ofs_0 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@52553.4]
  assign io_in_x355_outbuf_0_rPort_0_en_0 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@52552.4]
  assign io_in_x355_outbuf_0_rPort_0_backpressure = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@52551.4]
  assign io_in_x354_TVALID = x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TVALID; // @[sm_x647_outr_UnitPipe.scala 49:23:@52247.4]
  assign io_in_x354_TDATA = x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TDATA; // @[sm_x647_outr_UnitPipe.scala 49:23:@52245.4]
  assign io_sigsOut_smDoneIn_0 = x647_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@52153.4]
  assign io_sigsOut_smDoneIn_1 = x669_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@52442.4]
  assign x647_outr_UnitPipe_sm_clock = clock; // @[:@52069.4]
  assign x647_outr_UnitPipe_sm_reset = reset; // @[:@52070.4]
  assign x647_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@52150.4]
  assign x647_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@52152.4]
  assign x647_outr_UnitPipe_sm_io_doneIn_0 = x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@52120.4]
  assign x647_outr_UnitPipe_sm_io_doneIn_1 = x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@52121.4]
  assign x647_outr_UnitPipe_sm_io_ctrCopyDone_0 = x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@52167.4]
  assign x647_outr_UnitPipe_sm_io_ctrCopyDone_1 = x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@52168.4]
  assign RetimeWrapper_clock = clock; // @[:@52131.4]
  assign RetimeWrapper_reset = reset; // @[:@52132.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@52134.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@52133.4]
  assign RetimeWrapper_1_clock = clock; // @[:@52139.4]
  assign RetimeWrapper_1_reset = reset; // @[:@52140.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@52142.4]
  assign RetimeWrapper_1_io_in = x647_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@52141.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_clock = clock; // @[:@52170.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_reset = reset; // @[:@52171.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TVALID = io_in_x353_TVALID; // @[sm_x647_outr_UnitPipe.scala 48:23:@52238.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TDATA = io_in_x353_TDATA; // @[sm_x647_outr_UnitPipe.scala 48:23:@52236.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TID = io_in_x353_TID; // @[sm_x647_outr_UnitPipe.scala 48:23:@52232.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x353_TDEST = io_in_x353_TDEST; // @[sm_x647_outr_UnitPipe.scala 48:23:@52231.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_in_x354_TREADY = io_in_x354_TREADY; // @[sm_x647_outr_UnitPipe.scala 49:23:@52246.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x647_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x647_outr_UnitPipe.scala 92:22:@52263.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x647_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x647_outr_UnitPipe.scala 92:22:@52264.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x647_outr_UnitPipe_sm_io_childAck_0; // @[sm_x647_outr_UnitPipe.scala 92:22:@52259.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x647_outr_UnitPipe_sm_io_childAck_1; // @[sm_x647_outr_UnitPipe.scala 92:22:@52260.4]
  assign x647_outr_UnitPipe_kernelx647_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x647_outr_UnitPipe.scala 91:18:@52248.4]
  assign x669_outr_UnitPipe_sm_clock = clock; // @[:@52348.4]
  assign x669_outr_UnitPipe_sm_reset = reset; // @[:@52349.4]
  assign x669_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@52439.4]
  assign x669_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@52441.4]
  assign x669_outr_UnitPipe_sm_io_doneIn_0 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@52407.4]
  assign x669_outr_UnitPipe_sm_io_doneIn_1 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@52408.4]
  assign x669_outr_UnitPipe_sm_io_doneIn_2 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@52409.4]
  assign x669_outr_UnitPipe_sm_io_ctrCopyDone_0 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@52456.4]
  assign x669_outr_UnitPipe_sm_io_ctrCopyDone_1 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@52457.4]
  assign x669_outr_UnitPipe_sm_io_ctrCopyDone_2 = x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@52458.4]
  assign RetimeWrapper_2_clock = clock; // @[:@52420.4]
  assign RetimeWrapper_2_reset = reset; // @[:@52421.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@52423.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@52422.4]
  assign RetimeWrapper_3_clock = clock; // @[:@52428.4]
  assign RetimeWrapper_3_reset = reset; // @[:@52429.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@52431.4]
  assign RetimeWrapper_3_io_in = x669_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@52430.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_clock = clock; // @[:@52460.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_reset = reset; // @[:@52461.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x650_valid = io_in_x650_valid; // @[sm_x669_outr_UnitPipe.scala 58:23:@52540.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x649_ready = io_in_x649_ready; // @[sm_x669_outr_UnitPipe.scala 59:23:@52545.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x648_ready = io_in_x648_ready; // @[sm_x669_outr_UnitPipe.scala 60:23:@52549.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x355_outbuf_0_rPort_0_output_0 = io_in_x355_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@52550.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_in_x351_outdram_number = io_in_x351_outdram_number; // @[sm_x669_outr_UnitPipe.scala 62:31:@52555.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x669_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x669_outr_UnitPipe.scala 113:22:@52578.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x669_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x669_outr_UnitPipe.scala 113:22:@52579.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x669_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x669_outr_UnitPipe.scala 113:22:@52580.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x669_outr_UnitPipe_sm_io_childAck_0; // @[sm_x669_outr_UnitPipe.scala 113:22:@52572.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x669_outr_UnitPipe_sm_io_childAck_1; // @[sm_x669_outr_UnitPipe.scala 113:22:@52573.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x669_outr_UnitPipe_sm_io_childAck_2; // @[sm_x669_outr_UnitPipe.scala 113:22:@52574.4]
  assign x669_outr_UnitPipe_kernelx669_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x669_outr_UnitPipe.scala 112:18:@52556.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@52608.2]
  input          clock, // @[:@52609.4]
  input          reset, // @[:@52610.4]
  input          io_in_x353_TVALID, // @[:@52611.4]
  output         io_in_x353_TREADY, // @[:@52611.4]
  input  [255:0] io_in_x353_TDATA, // @[:@52611.4]
  input  [7:0]   io_in_x353_TID, // @[:@52611.4]
  input  [7:0]   io_in_x353_TDEST, // @[:@52611.4]
  output         io_in_x650_ready, // @[:@52611.4]
  input          io_in_x650_valid, // @[:@52611.4]
  input          io_in_x649_ready, // @[:@52611.4]
  output         io_in_x649_valid, // @[:@52611.4]
  output [31:0]  io_in_x649_bits_wdata_0, // @[:@52611.4]
  output         io_in_x649_bits_wstrb, // @[:@52611.4]
  input          io_in_x648_ready, // @[:@52611.4]
  output         io_in_x648_valid, // @[:@52611.4]
  output [63:0]  io_in_x648_bits_addr, // @[:@52611.4]
  output [31:0]  io_in_x648_bits_size, // @[:@52611.4]
  input  [63:0]  io_in_x351_outdram_number, // @[:@52611.4]
  output         io_in_x354_TVALID, // @[:@52611.4]
  input          io_in_x354_TREADY, // @[:@52611.4]
  output [255:0] io_in_x354_TDATA, // @[:@52611.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@52611.4]
  input          io_sigsIn_smChildAcks_0, // @[:@52611.4]
  output         io_sigsOut_smDoneIn_0, // @[:@52611.4]
  input          io_rr // @[:@52611.4]
);
  wire  x355_outbuf_0_clock; // @[m_x355_outbuf_0.scala 27:17:@52621.4]
  wire  x355_outbuf_0_reset; // @[m_x355_outbuf_0.scala 27:17:@52621.4]
  wire [20:0] x355_outbuf_0_io_rPort_0_ofs_0; // @[m_x355_outbuf_0.scala 27:17:@52621.4]
  wire  x355_outbuf_0_io_rPort_0_en_0; // @[m_x355_outbuf_0.scala 27:17:@52621.4]
  wire  x355_outbuf_0_io_rPort_0_backpressure; // @[m_x355_outbuf_0.scala 27:17:@52621.4]
  wire [31:0] x355_outbuf_0_io_rPort_0_output_0; // @[m_x355_outbuf_0.scala 27:17:@52621.4]
  wire  x724_sm_clock; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_reset; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_enable; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_done; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_ctrDone; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_ctrInc; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_parentAck; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_doneIn_0; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_doneIn_1; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_enableOut_0; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_enableOut_1; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_childAck_0; // @[sm_x724.scala 37:18:@52679.4]
  wire  x724_sm_io_childAck_1; // @[sm_x724.scala 37:18:@52679.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@52746.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@52746.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@52746.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@52746.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@52746.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@52754.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@52754.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@52754.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@52754.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@52754.4]
  wire  x724_kernelx724_concrete1_clock; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_reset; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x353_TVALID; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x353_TREADY; // @[sm_x724.scala 102:24:@52783.4]
  wire [255:0] x724_kernelx724_concrete1_io_in_x353_TDATA; // @[sm_x724.scala 102:24:@52783.4]
  wire [7:0] x724_kernelx724_concrete1_io_in_x353_TID; // @[sm_x724.scala 102:24:@52783.4]
  wire [7:0] x724_kernelx724_concrete1_io_in_x353_TDEST; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x650_ready; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x650_valid; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x649_ready; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x649_valid; // @[sm_x724.scala 102:24:@52783.4]
  wire [31:0] x724_kernelx724_concrete1_io_in_x649_bits_wdata_0; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x649_bits_wstrb; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x648_ready; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x648_valid; // @[sm_x724.scala 102:24:@52783.4]
  wire [63:0] x724_kernelx724_concrete1_io_in_x648_bits_addr; // @[sm_x724.scala 102:24:@52783.4]
  wire [31:0] x724_kernelx724_concrete1_io_in_x648_bits_size; // @[sm_x724.scala 102:24:@52783.4]
  wire [20:0] x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_en_0; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure; // @[sm_x724.scala 102:24:@52783.4]
  wire [31:0] x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_output_0; // @[sm_x724.scala 102:24:@52783.4]
  wire [63:0] x724_kernelx724_concrete1_io_in_x351_outdram_number; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x354_TVALID; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_in_x354_TREADY; // @[sm_x724.scala 102:24:@52783.4]
  wire [255:0] x724_kernelx724_concrete1_io_in_x354_TDATA; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x724.scala 102:24:@52783.4]
  wire  x724_kernelx724_concrete1_io_rr; // @[sm_x724.scala 102:24:@52783.4]
  wire  _T_266; // @[package.scala 100:49:@52712.4]
  reg  _T_269; // @[package.scala 48:56:@52713.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@52751.4 package.scala 96:25:@52752.4]
  wire  _T_289; // @[package.scala 96:25:@52759.4 package.scala 96:25:@52760.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@52762.4]
  x355_outbuf_0 x355_outbuf_0 ( // @[m_x355_outbuf_0.scala 27:17:@52621.4]
    .clock(x355_outbuf_0_clock),
    .reset(x355_outbuf_0_reset),
    .io_rPort_0_ofs_0(x355_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x355_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x355_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x355_outbuf_0_io_rPort_0_output_0)
  );
  x724_sm x724_sm ( // @[sm_x724.scala 37:18:@52679.4]
    .clock(x724_sm_clock),
    .reset(x724_sm_reset),
    .io_enable(x724_sm_io_enable),
    .io_done(x724_sm_io_done),
    .io_ctrDone(x724_sm_io_ctrDone),
    .io_ctrInc(x724_sm_io_ctrInc),
    .io_parentAck(x724_sm_io_parentAck),
    .io_doneIn_0(x724_sm_io_doneIn_0),
    .io_doneIn_1(x724_sm_io_doneIn_1),
    .io_enableOut_0(x724_sm_io_enableOut_0),
    .io_enableOut_1(x724_sm_io_enableOut_1),
    .io_childAck_0(x724_sm_io_childAck_0),
    .io_childAck_1(x724_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@52746.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@52754.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x724_kernelx724_concrete1 x724_kernelx724_concrete1 ( // @[sm_x724.scala 102:24:@52783.4]
    .clock(x724_kernelx724_concrete1_clock),
    .reset(x724_kernelx724_concrete1_reset),
    .io_in_x353_TVALID(x724_kernelx724_concrete1_io_in_x353_TVALID),
    .io_in_x353_TREADY(x724_kernelx724_concrete1_io_in_x353_TREADY),
    .io_in_x353_TDATA(x724_kernelx724_concrete1_io_in_x353_TDATA),
    .io_in_x353_TID(x724_kernelx724_concrete1_io_in_x353_TID),
    .io_in_x353_TDEST(x724_kernelx724_concrete1_io_in_x353_TDEST),
    .io_in_x650_ready(x724_kernelx724_concrete1_io_in_x650_ready),
    .io_in_x650_valid(x724_kernelx724_concrete1_io_in_x650_valid),
    .io_in_x649_ready(x724_kernelx724_concrete1_io_in_x649_ready),
    .io_in_x649_valid(x724_kernelx724_concrete1_io_in_x649_valid),
    .io_in_x649_bits_wdata_0(x724_kernelx724_concrete1_io_in_x649_bits_wdata_0),
    .io_in_x649_bits_wstrb(x724_kernelx724_concrete1_io_in_x649_bits_wstrb),
    .io_in_x648_ready(x724_kernelx724_concrete1_io_in_x648_ready),
    .io_in_x648_valid(x724_kernelx724_concrete1_io_in_x648_valid),
    .io_in_x648_bits_addr(x724_kernelx724_concrete1_io_in_x648_bits_addr),
    .io_in_x648_bits_size(x724_kernelx724_concrete1_io_in_x648_bits_size),
    .io_in_x355_outbuf_0_rPort_0_ofs_0(x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0),
    .io_in_x355_outbuf_0_rPort_0_en_0(x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_en_0),
    .io_in_x355_outbuf_0_rPort_0_backpressure(x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure),
    .io_in_x355_outbuf_0_rPort_0_output_0(x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_output_0),
    .io_in_x351_outdram_number(x724_kernelx724_concrete1_io_in_x351_outdram_number),
    .io_in_x354_TVALID(x724_kernelx724_concrete1_io_in_x354_TVALID),
    .io_in_x354_TREADY(x724_kernelx724_concrete1_io_in_x354_TREADY),
    .io_in_x354_TDATA(x724_kernelx724_concrete1_io_in_x354_TDATA),
    .io_sigsIn_smEnableOuts_0(x724_kernelx724_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x724_kernelx724_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x724_kernelx724_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x724_kernelx724_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x724_kernelx724_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x724_kernelx724_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x724_kernelx724_concrete1_io_rr)
  );
  assign _T_266 = x724_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@52712.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@52751.4 package.scala 96:25:@52752.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@52759.4 package.scala 96:25:@52760.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@52762.4]
  assign io_in_x353_TREADY = x724_kernelx724_concrete1_io_in_x353_TREADY; // @[sm_x724.scala 63:23:@52869.4]
  assign io_in_x650_ready = x724_kernelx724_concrete1_io_in_x650_ready; // @[sm_x724.scala 64:23:@52873.4]
  assign io_in_x649_valid = x724_kernelx724_concrete1_io_in_x649_valid; // @[sm_x724.scala 65:23:@52876.4]
  assign io_in_x649_bits_wdata_0 = x724_kernelx724_concrete1_io_in_x649_bits_wdata_0; // @[sm_x724.scala 65:23:@52875.4]
  assign io_in_x649_bits_wstrb = x724_kernelx724_concrete1_io_in_x649_bits_wstrb; // @[sm_x724.scala 65:23:@52874.4]
  assign io_in_x648_valid = x724_kernelx724_concrete1_io_in_x648_valid; // @[sm_x724.scala 66:23:@52880.4]
  assign io_in_x648_bits_addr = x724_kernelx724_concrete1_io_in_x648_bits_addr; // @[sm_x724.scala 66:23:@52879.4]
  assign io_in_x648_bits_size = x724_kernelx724_concrete1_io_in_x648_bits_size; // @[sm_x724.scala 66:23:@52878.4]
  assign io_in_x354_TVALID = x724_kernelx724_concrete1_io_in_x354_TVALID; // @[sm_x724.scala 69:23:@52896.4]
  assign io_in_x354_TDATA = x724_kernelx724_concrete1_io_in_x354_TDATA; // @[sm_x724.scala 69:23:@52894.4]
  assign io_sigsOut_smDoneIn_0 = x724_sm_io_done; // @[SpatialBlocks.scala 156:53:@52769.4]
  assign x355_outbuf_0_clock = clock; // @[:@52622.4]
  assign x355_outbuf_0_reset = reset; // @[:@52623.4]
  assign x355_outbuf_0_io_rPort_0_ofs_0 = x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@52885.4]
  assign x355_outbuf_0_io_rPort_0_en_0 = x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@52884.4]
  assign x355_outbuf_0_io_rPort_0_backpressure = x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@52883.4]
  assign x724_sm_clock = clock; // @[:@52680.4]
  assign x724_sm_reset = reset; // @[:@52681.4]
  assign x724_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@52766.4]
  assign x724_sm_io_ctrDone = x724_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@52716.4]
  assign x724_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@52768.4]
  assign x724_sm_io_doneIn_0 = x724_kernelx724_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@52736.4]
  assign x724_sm_io_doneIn_1 = x724_kernelx724_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@52737.4]
  assign RetimeWrapper_clock = clock; // @[:@52747.4]
  assign RetimeWrapper_reset = reset; // @[:@52748.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@52750.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@52749.4]
  assign RetimeWrapper_1_clock = clock; // @[:@52755.4]
  assign RetimeWrapper_1_reset = reset; // @[:@52756.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@52758.4]
  assign RetimeWrapper_1_io_in = x724_sm_io_done; // @[package.scala 94:16:@52757.4]
  assign x724_kernelx724_concrete1_clock = clock; // @[:@52784.4]
  assign x724_kernelx724_concrete1_reset = reset; // @[:@52785.4]
  assign x724_kernelx724_concrete1_io_in_x353_TVALID = io_in_x353_TVALID; // @[sm_x724.scala 63:23:@52870.4]
  assign x724_kernelx724_concrete1_io_in_x353_TDATA = io_in_x353_TDATA; // @[sm_x724.scala 63:23:@52868.4]
  assign x724_kernelx724_concrete1_io_in_x353_TID = io_in_x353_TID; // @[sm_x724.scala 63:23:@52864.4]
  assign x724_kernelx724_concrete1_io_in_x353_TDEST = io_in_x353_TDEST; // @[sm_x724.scala 63:23:@52863.4]
  assign x724_kernelx724_concrete1_io_in_x650_valid = io_in_x650_valid; // @[sm_x724.scala 64:23:@52872.4]
  assign x724_kernelx724_concrete1_io_in_x649_ready = io_in_x649_ready; // @[sm_x724.scala 65:23:@52877.4]
  assign x724_kernelx724_concrete1_io_in_x648_ready = io_in_x648_ready; // @[sm_x724.scala 66:23:@52881.4]
  assign x724_kernelx724_concrete1_io_in_x355_outbuf_0_rPort_0_output_0 = x355_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@52882.4]
  assign x724_kernelx724_concrete1_io_in_x351_outdram_number = io_in_x351_outdram_number; // @[sm_x724.scala 68:31:@52887.4]
  assign x724_kernelx724_concrete1_io_in_x354_TREADY = io_in_x354_TREADY; // @[sm_x724.scala 69:23:@52895.4]
  assign x724_kernelx724_concrete1_io_sigsIn_smEnableOuts_0 = x724_sm_io_enableOut_0; // @[sm_x724.scala 107:22:@52907.4]
  assign x724_kernelx724_concrete1_io_sigsIn_smEnableOuts_1 = x724_sm_io_enableOut_1; // @[sm_x724.scala 107:22:@52908.4]
  assign x724_kernelx724_concrete1_io_sigsIn_smChildAcks_0 = x724_sm_io_childAck_0; // @[sm_x724.scala 107:22:@52903.4]
  assign x724_kernelx724_concrete1_io_sigsIn_smChildAcks_1 = x724_sm_io_childAck_1; // @[sm_x724.scala 107:22:@52904.4]
  assign x724_kernelx724_concrete1_io_rr = io_rr; // @[sm_x724.scala 106:18:@52897.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@52930.2]
  input          clock, // @[:@52931.4]
  input          reset, // @[:@52932.4]
  input          io_enable, // @[:@52933.4]
  output         io_done, // @[:@52933.4]
  input          io_reset, // @[:@52933.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@52933.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@52933.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@52933.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@52933.4]
  output         io_memStreams_loads_0_data_ready, // @[:@52933.4]
  input          io_memStreams_loads_0_data_valid, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@52933.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@52933.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@52933.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@52933.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@52933.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@52933.4]
  input          io_memStreams_stores_0_data_ready, // @[:@52933.4]
  output         io_memStreams_stores_0_data_valid, // @[:@52933.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@52933.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@52933.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@52933.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@52933.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@52933.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@52933.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@52933.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@52933.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@52933.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@52933.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@52933.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@52933.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@52933.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@52933.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@52933.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@52933.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@52933.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@52933.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@52933.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@52933.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@52933.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@52933.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@52933.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@52933.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@52933.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@52933.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@52933.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@52933.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@52933.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@52933.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@52933.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@52933.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@52933.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@52933.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@52933.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@52933.4]
  output         io_heap_0_req_valid, // @[:@52933.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@52933.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@52933.4]
  input          io_heap_0_resp_valid, // @[:@52933.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@52933.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@52933.4]
  input  [63:0]  io_argIns_0, // @[:@52933.4]
  input  [63:0]  io_argIns_1, // @[:@52933.4]
  input          io_argOuts_0_port_ready, // @[:@52933.4]
  output         io_argOuts_0_port_valid, // @[:@52933.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@52933.4]
  input  [63:0]  io_argOuts_0_echo // @[:@52933.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@53081.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@53081.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@53081.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@53081.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@53099.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@53099.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@53099.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@53099.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@53099.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@53108.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@53108.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@53108.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@53108.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@53108.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@53108.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@53147.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@53179.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@53179.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@53179.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@53179.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@53179.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x353_TVALID; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x353_TREADY; // @[sm_RootController.scala 91:24:@53241.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x353_TDATA; // @[sm_RootController.scala 91:24:@53241.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x353_TID; // @[sm_RootController.scala 91:24:@53241.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x353_TDEST; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x650_ready; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x650_valid; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x649_ready; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x649_valid; // @[sm_RootController.scala 91:24:@53241.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x649_bits_wdata_0; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x649_bits_wstrb; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x648_ready; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x648_valid; // @[sm_RootController.scala 91:24:@53241.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x648_bits_addr; // @[sm_RootController.scala 91:24:@53241.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x648_bits_size; // @[sm_RootController.scala 91:24:@53241.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x351_outdram_number; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x354_TVALID; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_in_x354_TREADY; // @[sm_RootController.scala 91:24:@53241.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x354_TDATA; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@53241.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@53241.4]
  wire  _T_599; // @[package.scala 96:25:@53104.4 package.scala 96:25:@53105.4]
  wire  _T_664; // @[Main.scala 46:50:@53175.4]
  wire  _T_665; // @[Main.scala 46:59:@53176.4]
  wire  _T_677; // @[package.scala 100:49:@53196.4]
  reg  _T_680; // @[package.scala 48:56:@53197.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@53081.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@53099.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@53108.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@53147.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@53179.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@53241.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x353_TVALID(RootController_kernelRootController_concrete1_io_in_x353_TVALID),
    .io_in_x353_TREADY(RootController_kernelRootController_concrete1_io_in_x353_TREADY),
    .io_in_x353_TDATA(RootController_kernelRootController_concrete1_io_in_x353_TDATA),
    .io_in_x353_TID(RootController_kernelRootController_concrete1_io_in_x353_TID),
    .io_in_x353_TDEST(RootController_kernelRootController_concrete1_io_in_x353_TDEST),
    .io_in_x650_ready(RootController_kernelRootController_concrete1_io_in_x650_ready),
    .io_in_x650_valid(RootController_kernelRootController_concrete1_io_in_x650_valid),
    .io_in_x649_ready(RootController_kernelRootController_concrete1_io_in_x649_ready),
    .io_in_x649_valid(RootController_kernelRootController_concrete1_io_in_x649_valid),
    .io_in_x649_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x649_bits_wdata_0),
    .io_in_x649_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x649_bits_wstrb),
    .io_in_x648_ready(RootController_kernelRootController_concrete1_io_in_x648_ready),
    .io_in_x648_valid(RootController_kernelRootController_concrete1_io_in_x648_valid),
    .io_in_x648_bits_addr(RootController_kernelRootController_concrete1_io_in_x648_bits_addr),
    .io_in_x648_bits_size(RootController_kernelRootController_concrete1_io_in_x648_bits_size),
    .io_in_x351_outdram_number(RootController_kernelRootController_concrete1_io_in_x351_outdram_number),
    .io_in_x354_TVALID(RootController_kernelRootController_concrete1_io_in_x354_TVALID),
    .io_in_x354_TREADY(RootController_kernelRootController_concrete1_io_in_x354_TREADY),
    .io_in_x354_TDATA(RootController_kernelRootController_concrete1_io_in_x354_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@53104.4 package.scala 96:25:@53105.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@53175.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@53176.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@53196.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@53195.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x648_valid; // @[sm_RootController.scala 63:23:@53320.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x648_bits_addr; // @[sm_RootController.scala 63:23:@53319.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x648_bits_size; // @[sm_RootController.scala 63:23:@53318.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x649_valid; // @[sm_RootController.scala 62:23:@53316.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x649_bits_wdata_0; // @[sm_RootController.scala 62:23:@53315.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x649_bits_wstrb; // @[sm_RootController.scala 62:23:@53314.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x650_ready; // @[sm_RootController.scala 61:23:@53313.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x353_TREADY; // @[sm_RootController.scala 60:23:@53309.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x354_TVALID; // @[sm_RootController.scala 65:23:@53331.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x354_TDATA; // @[sm_RootController.scala 65:23:@53329.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 65:23:@53328.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 65:23:@53327.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 65:23:@53326.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 65:23:@53325.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 65:23:@53324.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 65:23:@53323.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@53082.4]
  assign SingleCounter_reset = reset; // @[:@53083.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@53097.4]
  assign RetimeWrapper_clock = clock; // @[:@53100.4]
  assign RetimeWrapper_reset = reset; // @[:@53101.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@53103.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@53102.4]
  assign SRFF_clock = clock; // @[:@53109.4]
  assign SRFF_reset = reset; // @[:@53110.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@53359.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@53193.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@53194.4]
  assign RootController_sm_clock = clock; // @[:@53148.4]
  assign RootController_sm_reset = reset; // @[:@53149.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@53192.4 SpatialBlocks.scala 140:18:@53226.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@53220.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@53200.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@53188.4 SpatialBlocks.scala 142:21:@53228.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@53217.4]
  assign RetimeWrapper_1_clock = clock; // @[:@53180.4]
  assign RetimeWrapper_1_reset = reset; // @[:@53181.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@53183.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@53182.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@53242.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@53243.4]
  assign RootController_kernelRootController_concrete1_io_in_x353_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 60:23:@53310.4]
  assign RootController_kernelRootController_concrete1_io_in_x353_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 60:23:@53308.4]
  assign RootController_kernelRootController_concrete1_io_in_x353_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 60:23:@53304.4]
  assign RootController_kernelRootController_concrete1_io_in_x353_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 60:23:@53303.4]
  assign RootController_kernelRootController_concrete1_io_in_x650_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 61:23:@53312.4]
  assign RootController_kernelRootController_concrete1_io_in_x649_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 62:23:@53317.4]
  assign RootController_kernelRootController_concrete1_io_in_x648_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 63:23:@53321.4]
  assign RootController_kernelRootController_concrete1_io_in_x351_outdram_number = io_argIns_1; // @[sm_RootController.scala 64:31:@53322.4]
  assign RootController_kernelRootController_concrete1_io_in_x354_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 65:23:@53330.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@53340.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@53338.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@53332.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@53361.2]
  input        clock, // @[:@53362.4]
  input        reset, // @[:@53363.4]
  input        io_enable, // @[:@53364.4]
  output [5:0] io_out, // @[:@53364.4]
  output [5:0] io_next // @[:@53364.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@53366.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@53367.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@53368.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@53373.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@53367.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@53368.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@53373.6]
  assign io_out = count; // @[Counter.scala 25:10:@53376.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@53377.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_25( // @[:@53413.2]
  input         clock, // @[:@53414.4]
  input         reset, // @[:@53415.4]
  input  [5:0]  io_raddr, // @[:@53416.4]
  input         io_wen, // @[:@53416.4]
  input  [5:0]  io_waddr, // @[:@53416.4]
  input  [63:0] io_wdata_addr, // @[:@53416.4]
  input  [31:0] io_wdata_size, // @[:@53416.4]
  output [63:0] io_rdata_addr, // @[:@53416.4]
  output [31:0] io_rdata_size // @[:@53416.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@53418.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@53418.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@53418.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@53418.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@53418.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@53418.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@53418.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@53418.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@53418.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@53432.4]
  wire  _T_20; // @[SRAM.scala 182:49:@53437.4]
  wire  _T_21; // @[SRAM.scala 182:37:@53438.4]
  reg  _T_24; // @[SRAM.scala 182:29:@53439.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@53442.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@53444.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@53418.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@53432.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@53437.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@53438.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@53444.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@53453.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@53452.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@53433.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@53434.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@53430.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@53436.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@53435.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@53431.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@53429.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@53428.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@53455.2]
  input         clock, // @[:@53456.4]
  input         reset, // @[:@53457.4]
  output        io_in_ready, // @[:@53458.4]
  input         io_in_valid, // @[:@53458.4]
  input  [63:0] io_in_bits_addr, // @[:@53458.4]
  input  [31:0] io_in_bits_size, // @[:@53458.4]
  input         io_out_ready, // @[:@53458.4]
  output        io_out_valid, // @[:@53458.4]
  output [63:0] io_out_bits_addr, // @[:@53458.4]
  output [31:0] io_out_bits_size // @[:@53458.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@53854.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@53854.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@53854.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@53854.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@53854.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@53864.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@53864.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@53864.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@53864.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@53864.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@53879.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@53879.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@53879.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@53879.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@53879.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@53879.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@53879.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@53879.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@53879.4]
  wire  writeEn; // @[FIFO.scala 30:29:@53852.4]
  wire  readEn; // @[FIFO.scala 31:29:@53853.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@53874.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@53875.4]
  wire  _T_824; // @[FIFO.scala 45:27:@53876.4]
  wire  empty; // @[FIFO.scala 45:24:@53877.4]
  wire  full; // @[FIFO.scala 46:23:@53878.4]
  wire  _T_827; // @[FIFO.scala 83:17:@53891.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@53892.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@53854.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@53864.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_25 SRAM ( // @[FIFO.scala 73:19:@53879.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@53852.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@53853.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@53875.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@53876.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@53877.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@53878.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@53891.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@53892.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@53898.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@53896.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@53889.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@53888.4]
  assign enqCounter_clock = clock; // @[:@53855.4]
  assign enqCounter_reset = reset; // @[:@53856.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@53862.4]
  assign deqCounter_clock = clock; // @[:@53865.4]
  assign deqCounter_reset = reset; // @[:@53866.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@53872.4]
  assign SRAM_clock = clock; // @[:@53880.4]
  assign SRAM_reset = reset; // @[:@53881.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@53883.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@53884.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@53885.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@53887.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@53886.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@53900.2]
  input        clock, // @[:@53901.4]
  input        reset, // @[:@53902.4]
  input        io_enable, // @[:@53903.4]
  output [3:0] io_out // @[:@53903.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@53905.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@53906.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@53907.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@53912.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@53906.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@53907.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@53912.6]
  assign io_out = count; // @[Counter.scala 25:10:@53915.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@53936.2]
  input        clock, // @[:@53937.4]
  input        reset, // @[:@53938.4]
  input        io_reset, // @[:@53939.4]
  input        io_enable, // @[:@53939.4]
  input  [1:0] io_stride, // @[:@53939.4]
  output [1:0] io_out, // @[:@53939.4]
  output [1:0] io_next // @[:@53939.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@53941.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@53942.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@53943.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@53948.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@53944.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@53942.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@53943.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@53948.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@53944.4]
  assign io_out = count; // @[Counter.scala 25:10:@53951.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@53952.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_26( // @[:@53988.2]
  input         clock, // @[:@53989.4]
  input         reset, // @[:@53990.4]
  input  [1:0]  io_raddr, // @[:@53991.4]
  input         io_wen, // @[:@53991.4]
  input  [1:0]  io_waddr, // @[:@53991.4]
  input  [31:0] io_wdata, // @[:@53991.4]
  output [31:0] io_rdata, // @[:@53991.4]
  input         io_backpressure // @[:@53991.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@53993.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@53993.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@53993.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@53993.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@53993.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@53993.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@53993.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@53993.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@53993.4]
  wire  _T_19; // @[SRAM.scala 182:49:@54011.4]
  wire  _T_20; // @[SRAM.scala 182:37:@54012.4]
  reg  _T_23; // @[SRAM.scala 182:29:@54013.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@54015.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@53993.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@54011.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@54012.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@54020.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@54007.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@54008.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@54005.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@54010.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@54009.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@54006.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@54004.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@54003.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@54022.2]
  input         clock, // @[:@54023.4]
  input         reset, // @[:@54024.4]
  output        io_in_ready, // @[:@54025.4]
  input         io_in_valid, // @[:@54025.4]
  input  [31:0] io_in_bits, // @[:@54025.4]
  input         io_out_ready, // @[:@54025.4]
  output        io_out_valid, // @[:@54025.4]
  output [31:0] io_out_bits // @[:@54025.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@54051.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@54051.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@54051.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@54051.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@54051.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@54051.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@54051.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@54061.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@54061.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@54061.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@54061.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@54061.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@54061.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@54061.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@54076.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@54076.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@54076.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@54076.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@54076.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@54076.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@54076.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@54076.4]
  wire  writeEn; // @[FIFO.scala 30:29:@54049.4]
  wire  readEn; // @[FIFO.scala 31:29:@54050.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@54071.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@54072.4]
  wire  _T_104; // @[FIFO.scala 45:27:@54073.4]
  wire  empty; // @[FIFO.scala 45:24:@54074.4]
  wire  full; // @[FIFO.scala 46:23:@54075.4]
  wire  _T_107; // @[FIFO.scala 83:17:@54086.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@54087.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@54051.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@54061.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_26 SRAM ( // @[FIFO.scala 73:19:@54076.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@54049.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@54050.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@54072.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@54073.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@54074.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@54075.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@54086.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@54087.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@54093.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@54091.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@54084.4]
  assign enqCounter_clock = clock; // @[:@54052.4]
  assign enqCounter_reset = reset; // @[:@54053.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@54059.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@54060.4]
  assign deqCounter_clock = clock; // @[:@54062.4]
  assign deqCounter_reset = reset; // @[:@54063.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@54069.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@54070.4]
  assign SRAM_clock = clock; // @[:@54077.4]
  assign SRAM_reset = reset; // @[:@54078.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@54080.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@54081.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@54082.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@54083.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@54085.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@56480.2]
  input         clock, // @[:@56481.4]
  input         reset, // @[:@56482.4]
  output        io_in_ready, // @[:@56483.4]
  input         io_in_valid, // @[:@56483.4]
  input  [31:0] io_in_bits_0, // @[:@56483.4]
  input         io_out_ready, // @[:@56483.4]
  output        io_out_valid, // @[:@56483.4]
  output [31:0] io_out_bits_0, // @[:@56483.4]
  output [31:0] io_out_bits_1, // @[:@56483.4]
  output [31:0] io_out_bits_2, // @[:@56483.4]
  output [31:0] io_out_bits_3, // @[:@56483.4]
  output [31:0] io_out_bits_4, // @[:@56483.4]
  output [31:0] io_out_bits_5, // @[:@56483.4]
  output [31:0] io_out_bits_6, // @[:@56483.4]
  output [31:0] io_out_bits_7, // @[:@56483.4]
  output [31:0] io_out_bits_8, // @[:@56483.4]
  output [31:0] io_out_bits_9, // @[:@56483.4]
  output [31:0] io_out_bits_10, // @[:@56483.4]
  output [31:0] io_out_bits_11, // @[:@56483.4]
  output [31:0] io_out_bits_12, // @[:@56483.4]
  output [31:0] io_out_bits_13, // @[:@56483.4]
  output [31:0] io_out_bits_14, // @[:@56483.4]
  output [31:0] io_out_bits_15 // @[:@56483.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@56487.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@56487.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@56487.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@56487.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@56498.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@56498.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@56498.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@56498.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@56511.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@56511.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@56511.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@56511.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@56511.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@56511.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@56511.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@56511.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@56546.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@56546.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@56546.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@56546.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@56546.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@56546.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@56546.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@56546.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@56581.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@56581.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@56581.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@56581.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@56581.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@56581.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@56581.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@56581.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@56616.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@56616.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@56616.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@56616.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@56616.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@56616.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@56616.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@56616.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@56651.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@56651.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@56651.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@56651.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@56651.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@56651.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@56651.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@56651.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@56686.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@56686.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@56686.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@56686.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@56686.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@56686.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@56686.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@56686.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@56721.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@56721.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@56721.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@56721.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@56721.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@56721.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@56721.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@56721.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@56756.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@56756.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@56756.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@56756.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@56756.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@56756.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@56756.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@56756.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@56791.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@56791.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@56791.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@56791.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@56791.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@56791.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@56791.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@56791.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@56826.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@56826.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@56826.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@56826.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@56826.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@56826.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@56826.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@56826.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@56861.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@56861.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@56861.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@56861.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@56861.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@56861.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@56861.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@56861.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@56896.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@56896.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@56896.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@56896.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@56896.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@56896.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@56896.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@56896.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@56931.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@56931.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@56931.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@56931.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@56931.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@56931.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@56931.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@56931.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@56966.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@56966.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@56966.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@56966.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@56966.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@56966.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@56966.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@56966.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@57001.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@57001.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@57001.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@57001.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@57001.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@57001.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@57001.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@57001.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@57036.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@57036.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@57036.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@57036.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@57036.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@57036.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@57036.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@57036.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@56486.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@56509.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@56536.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@56571.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@56606.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@56641.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@56676.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@56711.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@56746.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@56781.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@56816.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@56851.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@56886.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@56921.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@56956.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@56991.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@57026.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@57061.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57072.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57073.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57074.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57075.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57076.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57077.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57078.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57079.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57080.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57081.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57082.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57083.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57084.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57085.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57086.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@57103.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57087.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@57122.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@57123.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@57124.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@57125.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@57126.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@57127.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@57128.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@57129.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@57130.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@57131.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@57132.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@57133.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@57134.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@57135.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@56487.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@56498.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@56511.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@56546.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@56581.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@56616.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@56651.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@56686.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@56721.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@56756.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@56791.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@56826.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@56861.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@56896.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@56931.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@56966.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@57001.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@57036.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@56486.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@56509.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@56536.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@56571.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@56606.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@56641.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@56676.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@56711.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@56746.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@56781.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@56816.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@56851.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@56886.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@56921.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@56956.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@56991.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@57026.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@57061.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57072.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57073.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57074.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57075.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57076.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57077.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57078.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57079.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57080.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57081.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57082.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57083.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57084.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57085.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57086.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@57103.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@57071.4 FIFOVec.scala 49:42:@57087.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@57122.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@57123.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@57124.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@57125.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@57126.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@57127.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@57128.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@57129.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@57130.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@57131.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@57132.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@57133.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@57134.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@57135.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@57104.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@57138.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@57446.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@57447.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@57448.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@57449.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@57450.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@57451.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@57452.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@57453.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@57454.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@57455.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@57456.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@57457.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@57458.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@57459.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@57460.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@57461.4]
  assign enqCounter_clock = clock; // @[:@56488.4]
  assign enqCounter_reset = reset; // @[:@56489.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@56496.4]
  assign deqCounter_clock = clock; // @[:@56499.4]
  assign deqCounter_reset = reset; // @[:@56500.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@56507.4]
  assign fifos_0_clock = clock; // @[:@56512.4]
  assign fifos_0_reset = reset; // @[:@56513.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@56539.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56541.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56545.4]
  assign fifos_1_clock = clock; // @[:@56547.4]
  assign fifos_1_reset = reset; // @[:@56548.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@56574.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56576.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56580.4]
  assign fifos_2_clock = clock; // @[:@56582.4]
  assign fifos_2_reset = reset; // @[:@56583.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@56609.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56611.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56615.4]
  assign fifos_3_clock = clock; // @[:@56617.4]
  assign fifos_3_reset = reset; // @[:@56618.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@56644.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56646.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56650.4]
  assign fifos_4_clock = clock; // @[:@56652.4]
  assign fifos_4_reset = reset; // @[:@56653.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@56679.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56681.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56685.4]
  assign fifos_5_clock = clock; // @[:@56687.4]
  assign fifos_5_reset = reset; // @[:@56688.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@56714.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56716.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56720.4]
  assign fifos_6_clock = clock; // @[:@56722.4]
  assign fifos_6_reset = reset; // @[:@56723.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@56749.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56751.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56755.4]
  assign fifos_7_clock = clock; // @[:@56757.4]
  assign fifos_7_reset = reset; // @[:@56758.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@56784.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56786.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56790.4]
  assign fifos_8_clock = clock; // @[:@56792.4]
  assign fifos_8_reset = reset; // @[:@56793.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@56819.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56821.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56825.4]
  assign fifos_9_clock = clock; // @[:@56827.4]
  assign fifos_9_reset = reset; // @[:@56828.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@56854.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56856.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56860.4]
  assign fifos_10_clock = clock; // @[:@56862.4]
  assign fifos_10_reset = reset; // @[:@56863.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@56889.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56891.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56895.4]
  assign fifos_11_clock = clock; // @[:@56897.4]
  assign fifos_11_reset = reset; // @[:@56898.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@56924.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56926.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56930.4]
  assign fifos_12_clock = clock; // @[:@56932.4]
  assign fifos_12_reset = reset; // @[:@56933.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@56959.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56961.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@56965.4]
  assign fifos_13_clock = clock; // @[:@56967.4]
  assign fifos_13_reset = reset; // @[:@56968.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@56994.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@56996.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@57000.4]
  assign fifos_14_clock = clock; // @[:@57002.4]
  assign fifos_14_reset = reset; // @[:@57003.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@57029.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@57031.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@57035.4]
  assign fifos_15_clock = clock; // @[:@57037.4]
  assign fifos_15_reset = reset; // @[:@57038.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@57064.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@57066.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@57070.4]
endmodule
module FFRAM( // @[:@57535.2]
  input        clock, // @[:@57536.4]
  input        reset, // @[:@57537.4]
  input  [1:0] io_raddr, // @[:@57538.4]
  input        io_wen, // @[:@57538.4]
  input  [1:0] io_waddr, // @[:@57538.4]
  input        io_wdata, // @[:@57538.4]
  output       io_rdata, // @[:@57538.4]
  input        io_banks_0_wdata_valid, // @[:@57538.4]
  input        io_banks_0_wdata_bits, // @[:@57538.4]
  input        io_banks_1_wdata_valid, // @[:@57538.4]
  input        io_banks_1_wdata_bits, // @[:@57538.4]
  input        io_banks_2_wdata_valid, // @[:@57538.4]
  input        io_banks_2_wdata_bits, // @[:@57538.4]
  input        io_banks_3_wdata_valid, // @[:@57538.4]
  input        io_banks_3_wdata_bits // @[:@57538.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@57542.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@57543.4]
  wire  _T_89; // @[SRAM.scala 148:25:@57544.4]
  wire  _T_90; // @[SRAM.scala 148:15:@57545.4]
  wire  _T_91; // @[SRAM.scala 149:15:@57547.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@57546.4]
  reg  regs_1; // @[SRAM.scala 145:20:@57553.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@57554.4]
  wire  _T_98; // @[SRAM.scala 148:25:@57555.4]
  wire  _T_99; // @[SRAM.scala 148:15:@57556.4]
  wire  _T_100; // @[SRAM.scala 149:15:@57558.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@57557.4]
  reg  regs_2; // @[SRAM.scala 145:20:@57564.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@57565.4]
  wire  _T_107; // @[SRAM.scala 148:25:@57566.4]
  wire  _T_108; // @[SRAM.scala 148:15:@57567.4]
  wire  _T_109; // @[SRAM.scala 149:15:@57569.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@57568.4]
  reg  regs_3; // @[SRAM.scala 145:20:@57575.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@57576.4]
  wire  _T_116; // @[SRAM.scala 148:25:@57577.4]
  wire  _T_117; // @[SRAM.scala 148:15:@57578.4]
  wire  _T_118; // @[SRAM.scala 149:15:@57580.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@57579.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@57589.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@57589.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@57543.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@57544.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@57545.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@57547.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@57546.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@57554.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@57555.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@57556.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@57558.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@57557.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@57565.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@57566.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@57567.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@57569.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@57568.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@57576.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@57577.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@57578.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@57580.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@57579.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@57589.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@57589.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@57589.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@57591.2]
  input   clock, // @[:@57592.4]
  input   reset, // @[:@57593.4]
  output  io_in_ready, // @[:@57594.4]
  input   io_in_valid, // @[:@57594.4]
  input   io_in_bits, // @[:@57594.4]
  input   io_out_ready, // @[:@57594.4]
  output  io_out_valid, // @[:@57594.4]
  output  io_out_bits // @[:@57594.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@57620.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@57620.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@57620.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@57620.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@57620.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@57620.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@57620.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@57630.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@57630.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@57630.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@57630.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@57630.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@57630.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@57630.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@57645.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@57645.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@57645.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@57645.4]
  wire  writeEn; // @[FIFO.scala 30:29:@57618.4]
  wire  readEn; // @[FIFO.scala 31:29:@57619.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@57640.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@57641.4]
  wire  _T_104; // @[FIFO.scala 45:27:@57642.4]
  wire  empty; // @[FIFO.scala 45:24:@57643.4]
  wire  full; // @[FIFO.scala 46:23:@57644.4]
  wire  _T_157; // @[FIFO.scala 83:17:@57731.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@57732.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@57620.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@57630.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@57645.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@57618.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@57619.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@57641.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@57642.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@57643.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@57644.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@57731.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@57732.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@57738.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@57736.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@57670.4]
  assign enqCounter_clock = clock; // @[:@57621.4]
  assign enqCounter_reset = reset; // @[:@57622.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@57628.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@57629.4]
  assign deqCounter_clock = clock; // @[:@57631.4]
  assign deqCounter_reset = reset; // @[:@57632.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@57638.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@57639.4]
  assign FFRAM_clock = clock; // @[:@57646.4]
  assign FFRAM_reset = reset; // @[:@57647.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@57666.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@57667.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@57668.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@57669.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@57672.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@57671.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@57675.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@57674.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@57678.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@57677.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@57681.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@57680.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@61355.2]
  input   clock, // @[:@61356.4]
  input   reset, // @[:@61357.4]
  output  io_in_ready, // @[:@61358.4]
  input   io_in_valid, // @[:@61358.4]
  input   io_in_bits_0, // @[:@61358.4]
  input   io_out_ready, // @[:@61358.4]
  output  io_out_valid, // @[:@61358.4]
  output  io_out_bits_0, // @[:@61358.4]
  output  io_out_bits_1, // @[:@61358.4]
  output  io_out_bits_2, // @[:@61358.4]
  output  io_out_bits_3, // @[:@61358.4]
  output  io_out_bits_4, // @[:@61358.4]
  output  io_out_bits_5, // @[:@61358.4]
  output  io_out_bits_6, // @[:@61358.4]
  output  io_out_bits_7, // @[:@61358.4]
  output  io_out_bits_8, // @[:@61358.4]
  output  io_out_bits_9, // @[:@61358.4]
  output  io_out_bits_10, // @[:@61358.4]
  output  io_out_bits_11, // @[:@61358.4]
  output  io_out_bits_12, // @[:@61358.4]
  output  io_out_bits_13, // @[:@61358.4]
  output  io_out_bits_14, // @[:@61358.4]
  output  io_out_bits_15 // @[:@61358.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@61362.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@61362.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@61362.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@61362.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@61373.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@61373.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@61373.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@61373.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@61386.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@61421.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@61456.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@61491.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@61526.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@61561.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@61596.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@61631.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@61666.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@61701.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@61736.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@61771.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@61806.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@61841.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@61876.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@61911.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@61911.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@61911.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@61911.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@61911.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@61911.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@61911.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@61911.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@61361.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@61384.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@61411.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@61446.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@61481.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@61516.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@61551.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@61586.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@61621.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@61656.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@61691.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@61726.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@61761.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@61796.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@61831.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@61866.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@61901.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@61936.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61947.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61948.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61949.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61950.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61951.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61952.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61953.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61954.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61955.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61956.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61957.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61958.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61959.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61960.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61961.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@61978.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61962.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@61997.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@61998.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@61999.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@62000.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@62001.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@62002.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@62003.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@62004.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@62005.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@62006.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@62007.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@62008.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@62009.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@62010.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@61362.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@61373.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@61386.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@61421.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@61456.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@61491.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@61526.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@61561.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@61596.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@61631.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@61666.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@61701.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@61736.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@61771.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@61806.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@61841.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@61876.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@61911.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@61361.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@61384.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@61411.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@61446.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@61481.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@61516.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@61551.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@61586.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@61621.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@61656.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@61691.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@61726.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@61761.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@61796.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@61831.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@61866.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@61901.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@61936.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61947.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61948.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61949.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61950.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61951.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61952.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61953.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61954.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61955.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61956.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61957.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61958.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61959.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61960.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61961.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@61978.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@61946.4 FIFOVec.scala 49:42:@61962.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@61997.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@61998.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@61999.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@62000.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@62001.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@62002.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@62003.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@62004.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@62005.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@62006.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@62007.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@62008.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@62009.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@62010.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@61979.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@62013.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@62321.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@62322.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@62323.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@62324.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@62325.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@62326.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@62327.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@62328.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@62329.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@62330.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@62331.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@62332.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@62333.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@62334.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@62335.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@62336.4]
  assign enqCounter_clock = clock; // @[:@61363.4]
  assign enqCounter_reset = reset; // @[:@61364.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@61371.4]
  assign deqCounter_clock = clock; // @[:@61374.4]
  assign deqCounter_reset = reset; // @[:@61375.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@61382.4]
  assign fifos_0_clock = clock; // @[:@61387.4]
  assign fifos_0_reset = reset; // @[:@61388.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@61414.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61416.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61420.4]
  assign fifos_1_clock = clock; // @[:@61422.4]
  assign fifos_1_reset = reset; // @[:@61423.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@61449.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61451.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61455.4]
  assign fifos_2_clock = clock; // @[:@61457.4]
  assign fifos_2_reset = reset; // @[:@61458.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@61484.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61486.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61490.4]
  assign fifos_3_clock = clock; // @[:@61492.4]
  assign fifos_3_reset = reset; // @[:@61493.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@61519.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61521.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61525.4]
  assign fifos_4_clock = clock; // @[:@61527.4]
  assign fifos_4_reset = reset; // @[:@61528.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@61554.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61556.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61560.4]
  assign fifos_5_clock = clock; // @[:@61562.4]
  assign fifos_5_reset = reset; // @[:@61563.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@61589.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61591.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61595.4]
  assign fifos_6_clock = clock; // @[:@61597.4]
  assign fifos_6_reset = reset; // @[:@61598.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@61624.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61626.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61630.4]
  assign fifos_7_clock = clock; // @[:@61632.4]
  assign fifos_7_reset = reset; // @[:@61633.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@61659.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61661.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61665.4]
  assign fifos_8_clock = clock; // @[:@61667.4]
  assign fifos_8_reset = reset; // @[:@61668.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@61694.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61696.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61700.4]
  assign fifos_9_clock = clock; // @[:@61702.4]
  assign fifos_9_reset = reset; // @[:@61703.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@61729.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61731.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61735.4]
  assign fifos_10_clock = clock; // @[:@61737.4]
  assign fifos_10_reset = reset; // @[:@61738.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@61764.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61766.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61770.4]
  assign fifos_11_clock = clock; // @[:@61772.4]
  assign fifos_11_reset = reset; // @[:@61773.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@61799.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61801.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61805.4]
  assign fifos_12_clock = clock; // @[:@61807.4]
  assign fifos_12_reset = reset; // @[:@61808.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@61834.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61836.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61840.4]
  assign fifos_13_clock = clock; // @[:@61842.4]
  assign fifos_13_reset = reset; // @[:@61843.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@61869.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61871.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61875.4]
  assign fifos_14_clock = clock; // @[:@61877.4]
  assign fifos_14_reset = reset; // @[:@61878.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@61904.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61906.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61910.4]
  assign fifos_15_clock = clock; // @[:@61912.4]
  assign fifos_15_reset = reset; // @[:@61913.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@61939.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@61941.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@61945.4]
endmodule
module FIFOWidthConvert( // @[:@62338.2]
  input         clock, // @[:@62339.4]
  input         reset, // @[:@62340.4]
  output        io_in_ready, // @[:@62341.4]
  input         io_in_valid, // @[:@62341.4]
  input  [31:0] io_in_bits_data_0, // @[:@62341.4]
  input         io_in_bits_strobe, // @[:@62341.4]
  input         io_out_ready, // @[:@62341.4]
  output        io_out_valid, // @[:@62341.4]
  output [31:0] io_out_bits_data_0, // @[:@62341.4]
  output [31:0] io_out_bits_data_1, // @[:@62341.4]
  output [31:0] io_out_bits_data_2, // @[:@62341.4]
  output [31:0] io_out_bits_data_3, // @[:@62341.4]
  output [31:0] io_out_bits_data_4, // @[:@62341.4]
  output [31:0] io_out_bits_data_5, // @[:@62341.4]
  output [31:0] io_out_bits_data_6, // @[:@62341.4]
  output [31:0] io_out_bits_data_7, // @[:@62341.4]
  output [31:0] io_out_bits_data_8, // @[:@62341.4]
  output [31:0] io_out_bits_data_9, // @[:@62341.4]
  output [31:0] io_out_bits_data_10, // @[:@62341.4]
  output [31:0] io_out_bits_data_11, // @[:@62341.4]
  output [31:0] io_out_bits_data_12, // @[:@62341.4]
  output [31:0] io_out_bits_data_13, // @[:@62341.4]
  output [31:0] io_out_bits_data_14, // @[:@62341.4]
  output [31:0] io_out_bits_data_15, // @[:@62341.4]
  output [63:0] io_out_bits_strobe // @[:@62341.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@62343.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@62384.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@62443.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@62449.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@62507.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@62513.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@62514.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@62518.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@62522.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@62526.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@62530.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@62534.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@62538.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@62542.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@62546.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@62550.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@62554.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@62558.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@62562.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@62566.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@62570.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@62574.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@62651.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@62660.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@62669.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@62678.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@62687.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@62696.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@62704.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@62343.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@62384.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@62443.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@62449.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@62507.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@62513.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@62514.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@62518.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@62522.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@62526.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@62530.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@62534.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@62538.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@62542.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@62546.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@62550.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@62554.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@62558.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@62562.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@62566.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@62570.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@62574.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@62651.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@62660.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@62669.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@62678.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@62687.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@62696.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@62704.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@62433.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@62434.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@62483.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@62484.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@62485.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@62486.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@62487.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@62488.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@62489.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@62490.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@62491.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@62492.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@62493.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@62494.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@62495.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@62496.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@62497.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@62498.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@62706.4]
  assign FIFOVec_clock = clock; // @[:@62344.4]
  assign FIFOVec_reset = reset; // @[:@62345.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@62430.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@62429.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@62707.4]
  assign FIFOVec_1_clock = clock; // @[:@62385.4]
  assign FIFOVec_1_reset = reset; // @[:@62386.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@62432.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@62431.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@62708.4]
endmodule
module FFRAM_16( // @[:@62746.2]
  input        clock, // @[:@62747.4]
  input        reset, // @[:@62748.4]
  input  [5:0] io_raddr, // @[:@62749.4]
  input        io_wen, // @[:@62749.4]
  input  [5:0] io_waddr, // @[:@62749.4]
  input        io_wdata, // @[:@62749.4]
  output       io_rdata, // @[:@62749.4]
  input        io_banks_0_wdata_valid, // @[:@62749.4]
  input        io_banks_0_wdata_bits, // @[:@62749.4]
  input        io_banks_1_wdata_valid, // @[:@62749.4]
  input        io_banks_1_wdata_bits, // @[:@62749.4]
  input        io_banks_2_wdata_valid, // @[:@62749.4]
  input        io_banks_2_wdata_bits, // @[:@62749.4]
  input        io_banks_3_wdata_valid, // @[:@62749.4]
  input        io_banks_3_wdata_bits, // @[:@62749.4]
  input        io_banks_4_wdata_valid, // @[:@62749.4]
  input        io_banks_4_wdata_bits, // @[:@62749.4]
  input        io_banks_5_wdata_valid, // @[:@62749.4]
  input        io_banks_5_wdata_bits, // @[:@62749.4]
  input        io_banks_6_wdata_valid, // @[:@62749.4]
  input        io_banks_6_wdata_bits, // @[:@62749.4]
  input        io_banks_7_wdata_valid, // @[:@62749.4]
  input        io_banks_7_wdata_bits, // @[:@62749.4]
  input        io_banks_8_wdata_valid, // @[:@62749.4]
  input        io_banks_8_wdata_bits, // @[:@62749.4]
  input        io_banks_9_wdata_valid, // @[:@62749.4]
  input        io_banks_9_wdata_bits, // @[:@62749.4]
  input        io_banks_10_wdata_valid, // @[:@62749.4]
  input        io_banks_10_wdata_bits, // @[:@62749.4]
  input        io_banks_11_wdata_valid, // @[:@62749.4]
  input        io_banks_11_wdata_bits, // @[:@62749.4]
  input        io_banks_12_wdata_valid, // @[:@62749.4]
  input        io_banks_12_wdata_bits, // @[:@62749.4]
  input        io_banks_13_wdata_valid, // @[:@62749.4]
  input        io_banks_13_wdata_bits, // @[:@62749.4]
  input        io_banks_14_wdata_valid, // @[:@62749.4]
  input        io_banks_14_wdata_bits, // @[:@62749.4]
  input        io_banks_15_wdata_valid, // @[:@62749.4]
  input        io_banks_15_wdata_bits, // @[:@62749.4]
  input        io_banks_16_wdata_valid, // @[:@62749.4]
  input        io_banks_16_wdata_bits, // @[:@62749.4]
  input        io_banks_17_wdata_valid, // @[:@62749.4]
  input        io_banks_17_wdata_bits, // @[:@62749.4]
  input        io_banks_18_wdata_valid, // @[:@62749.4]
  input        io_banks_18_wdata_bits, // @[:@62749.4]
  input        io_banks_19_wdata_valid, // @[:@62749.4]
  input        io_banks_19_wdata_bits, // @[:@62749.4]
  input        io_banks_20_wdata_valid, // @[:@62749.4]
  input        io_banks_20_wdata_bits, // @[:@62749.4]
  input        io_banks_21_wdata_valid, // @[:@62749.4]
  input        io_banks_21_wdata_bits, // @[:@62749.4]
  input        io_banks_22_wdata_valid, // @[:@62749.4]
  input        io_banks_22_wdata_bits, // @[:@62749.4]
  input        io_banks_23_wdata_valid, // @[:@62749.4]
  input        io_banks_23_wdata_bits, // @[:@62749.4]
  input        io_banks_24_wdata_valid, // @[:@62749.4]
  input        io_banks_24_wdata_bits, // @[:@62749.4]
  input        io_banks_25_wdata_valid, // @[:@62749.4]
  input        io_banks_25_wdata_bits, // @[:@62749.4]
  input        io_banks_26_wdata_valid, // @[:@62749.4]
  input        io_banks_26_wdata_bits, // @[:@62749.4]
  input        io_banks_27_wdata_valid, // @[:@62749.4]
  input        io_banks_27_wdata_bits, // @[:@62749.4]
  input        io_banks_28_wdata_valid, // @[:@62749.4]
  input        io_banks_28_wdata_bits, // @[:@62749.4]
  input        io_banks_29_wdata_valid, // @[:@62749.4]
  input        io_banks_29_wdata_bits, // @[:@62749.4]
  input        io_banks_30_wdata_valid, // @[:@62749.4]
  input        io_banks_30_wdata_bits, // @[:@62749.4]
  input        io_banks_31_wdata_valid, // @[:@62749.4]
  input        io_banks_31_wdata_bits, // @[:@62749.4]
  input        io_banks_32_wdata_valid, // @[:@62749.4]
  input        io_banks_32_wdata_bits, // @[:@62749.4]
  input        io_banks_33_wdata_valid, // @[:@62749.4]
  input        io_banks_33_wdata_bits, // @[:@62749.4]
  input        io_banks_34_wdata_valid, // @[:@62749.4]
  input        io_banks_34_wdata_bits, // @[:@62749.4]
  input        io_banks_35_wdata_valid, // @[:@62749.4]
  input        io_banks_35_wdata_bits, // @[:@62749.4]
  input        io_banks_36_wdata_valid, // @[:@62749.4]
  input        io_banks_36_wdata_bits, // @[:@62749.4]
  input        io_banks_37_wdata_valid, // @[:@62749.4]
  input        io_banks_37_wdata_bits, // @[:@62749.4]
  input        io_banks_38_wdata_valid, // @[:@62749.4]
  input        io_banks_38_wdata_bits, // @[:@62749.4]
  input        io_banks_39_wdata_valid, // @[:@62749.4]
  input        io_banks_39_wdata_bits, // @[:@62749.4]
  input        io_banks_40_wdata_valid, // @[:@62749.4]
  input        io_banks_40_wdata_bits, // @[:@62749.4]
  input        io_banks_41_wdata_valid, // @[:@62749.4]
  input        io_banks_41_wdata_bits, // @[:@62749.4]
  input        io_banks_42_wdata_valid, // @[:@62749.4]
  input        io_banks_42_wdata_bits, // @[:@62749.4]
  input        io_banks_43_wdata_valid, // @[:@62749.4]
  input        io_banks_43_wdata_bits, // @[:@62749.4]
  input        io_banks_44_wdata_valid, // @[:@62749.4]
  input        io_banks_44_wdata_bits, // @[:@62749.4]
  input        io_banks_45_wdata_valid, // @[:@62749.4]
  input        io_banks_45_wdata_bits, // @[:@62749.4]
  input        io_banks_46_wdata_valid, // @[:@62749.4]
  input        io_banks_46_wdata_bits, // @[:@62749.4]
  input        io_banks_47_wdata_valid, // @[:@62749.4]
  input        io_banks_47_wdata_bits, // @[:@62749.4]
  input        io_banks_48_wdata_valid, // @[:@62749.4]
  input        io_banks_48_wdata_bits, // @[:@62749.4]
  input        io_banks_49_wdata_valid, // @[:@62749.4]
  input        io_banks_49_wdata_bits, // @[:@62749.4]
  input        io_banks_50_wdata_valid, // @[:@62749.4]
  input        io_banks_50_wdata_bits, // @[:@62749.4]
  input        io_banks_51_wdata_valid, // @[:@62749.4]
  input        io_banks_51_wdata_bits, // @[:@62749.4]
  input        io_banks_52_wdata_valid, // @[:@62749.4]
  input        io_banks_52_wdata_bits, // @[:@62749.4]
  input        io_banks_53_wdata_valid, // @[:@62749.4]
  input        io_banks_53_wdata_bits, // @[:@62749.4]
  input        io_banks_54_wdata_valid, // @[:@62749.4]
  input        io_banks_54_wdata_bits, // @[:@62749.4]
  input        io_banks_55_wdata_valid, // @[:@62749.4]
  input        io_banks_55_wdata_bits, // @[:@62749.4]
  input        io_banks_56_wdata_valid, // @[:@62749.4]
  input        io_banks_56_wdata_bits, // @[:@62749.4]
  input        io_banks_57_wdata_valid, // @[:@62749.4]
  input        io_banks_57_wdata_bits, // @[:@62749.4]
  input        io_banks_58_wdata_valid, // @[:@62749.4]
  input        io_banks_58_wdata_bits, // @[:@62749.4]
  input        io_banks_59_wdata_valid, // @[:@62749.4]
  input        io_banks_59_wdata_bits, // @[:@62749.4]
  input        io_banks_60_wdata_valid, // @[:@62749.4]
  input        io_banks_60_wdata_bits, // @[:@62749.4]
  input        io_banks_61_wdata_valid, // @[:@62749.4]
  input        io_banks_61_wdata_bits, // @[:@62749.4]
  input        io_banks_62_wdata_valid, // @[:@62749.4]
  input        io_banks_62_wdata_bits, // @[:@62749.4]
  input        io_banks_63_wdata_valid, // @[:@62749.4]
  input        io_banks_63_wdata_bits // @[:@62749.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@62753.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@62754.4]
  wire  _T_689; // @[SRAM.scala 148:25:@62755.4]
  wire  _T_690; // @[SRAM.scala 148:15:@62756.4]
  wire  _T_691; // @[SRAM.scala 149:15:@62758.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@62757.4]
  reg  regs_1; // @[SRAM.scala 145:20:@62764.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@62765.4]
  wire  _T_698; // @[SRAM.scala 148:25:@62766.4]
  wire  _T_699; // @[SRAM.scala 148:15:@62767.4]
  wire  _T_700; // @[SRAM.scala 149:15:@62769.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@62768.4]
  reg  regs_2; // @[SRAM.scala 145:20:@62775.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@62776.4]
  wire  _T_707; // @[SRAM.scala 148:25:@62777.4]
  wire  _T_708; // @[SRAM.scala 148:15:@62778.4]
  wire  _T_709; // @[SRAM.scala 149:15:@62780.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@62779.4]
  reg  regs_3; // @[SRAM.scala 145:20:@62786.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@62787.4]
  wire  _T_716; // @[SRAM.scala 148:25:@62788.4]
  wire  _T_717; // @[SRAM.scala 148:15:@62789.4]
  wire  _T_718; // @[SRAM.scala 149:15:@62791.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@62790.4]
  reg  regs_4; // @[SRAM.scala 145:20:@62797.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@62798.4]
  wire  _T_725; // @[SRAM.scala 148:25:@62799.4]
  wire  _T_726; // @[SRAM.scala 148:15:@62800.4]
  wire  _T_727; // @[SRAM.scala 149:15:@62802.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@62801.4]
  reg  regs_5; // @[SRAM.scala 145:20:@62808.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@62809.4]
  wire  _T_734; // @[SRAM.scala 148:25:@62810.4]
  wire  _T_735; // @[SRAM.scala 148:15:@62811.4]
  wire  _T_736; // @[SRAM.scala 149:15:@62813.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@62812.4]
  reg  regs_6; // @[SRAM.scala 145:20:@62819.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@62820.4]
  wire  _T_743; // @[SRAM.scala 148:25:@62821.4]
  wire  _T_744; // @[SRAM.scala 148:15:@62822.4]
  wire  _T_745; // @[SRAM.scala 149:15:@62824.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@62823.4]
  reg  regs_7; // @[SRAM.scala 145:20:@62830.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@62831.4]
  wire  _T_752; // @[SRAM.scala 148:25:@62832.4]
  wire  _T_753; // @[SRAM.scala 148:15:@62833.4]
  wire  _T_754; // @[SRAM.scala 149:15:@62835.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@62834.4]
  reg  regs_8; // @[SRAM.scala 145:20:@62841.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@62842.4]
  wire  _T_761; // @[SRAM.scala 148:25:@62843.4]
  wire  _T_762; // @[SRAM.scala 148:15:@62844.4]
  wire  _T_763; // @[SRAM.scala 149:15:@62846.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@62845.4]
  reg  regs_9; // @[SRAM.scala 145:20:@62852.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@62853.4]
  wire  _T_770; // @[SRAM.scala 148:25:@62854.4]
  wire  _T_771; // @[SRAM.scala 148:15:@62855.4]
  wire  _T_772; // @[SRAM.scala 149:15:@62857.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@62856.4]
  reg  regs_10; // @[SRAM.scala 145:20:@62863.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@62864.4]
  wire  _T_779; // @[SRAM.scala 148:25:@62865.4]
  wire  _T_780; // @[SRAM.scala 148:15:@62866.4]
  wire  _T_781; // @[SRAM.scala 149:15:@62868.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@62867.4]
  reg  regs_11; // @[SRAM.scala 145:20:@62874.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@62875.4]
  wire  _T_788; // @[SRAM.scala 148:25:@62876.4]
  wire  _T_789; // @[SRAM.scala 148:15:@62877.4]
  wire  _T_790; // @[SRAM.scala 149:15:@62879.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@62878.4]
  reg  regs_12; // @[SRAM.scala 145:20:@62885.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@62886.4]
  wire  _T_797; // @[SRAM.scala 148:25:@62887.4]
  wire  _T_798; // @[SRAM.scala 148:15:@62888.4]
  wire  _T_799; // @[SRAM.scala 149:15:@62890.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@62889.4]
  reg  regs_13; // @[SRAM.scala 145:20:@62896.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@62897.4]
  wire  _T_806; // @[SRAM.scala 148:25:@62898.4]
  wire  _T_807; // @[SRAM.scala 148:15:@62899.4]
  wire  _T_808; // @[SRAM.scala 149:15:@62901.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@62900.4]
  reg  regs_14; // @[SRAM.scala 145:20:@62907.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@62908.4]
  wire  _T_815; // @[SRAM.scala 148:25:@62909.4]
  wire  _T_816; // @[SRAM.scala 148:15:@62910.4]
  wire  _T_817; // @[SRAM.scala 149:15:@62912.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@62911.4]
  reg  regs_15; // @[SRAM.scala 145:20:@62918.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@62919.4]
  wire  _T_824; // @[SRAM.scala 148:25:@62920.4]
  wire  _T_825; // @[SRAM.scala 148:15:@62921.4]
  wire  _T_826; // @[SRAM.scala 149:15:@62923.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@62922.4]
  reg  regs_16; // @[SRAM.scala 145:20:@62929.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@62930.4]
  wire  _T_833; // @[SRAM.scala 148:25:@62931.4]
  wire  _T_834; // @[SRAM.scala 148:15:@62932.4]
  wire  _T_835; // @[SRAM.scala 149:15:@62934.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@62933.4]
  reg  regs_17; // @[SRAM.scala 145:20:@62940.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@62941.4]
  wire  _T_842; // @[SRAM.scala 148:25:@62942.4]
  wire  _T_843; // @[SRAM.scala 148:15:@62943.4]
  wire  _T_844; // @[SRAM.scala 149:15:@62945.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@62944.4]
  reg  regs_18; // @[SRAM.scala 145:20:@62951.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@62952.4]
  wire  _T_851; // @[SRAM.scala 148:25:@62953.4]
  wire  _T_852; // @[SRAM.scala 148:15:@62954.4]
  wire  _T_853; // @[SRAM.scala 149:15:@62956.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@62955.4]
  reg  regs_19; // @[SRAM.scala 145:20:@62962.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@62963.4]
  wire  _T_860; // @[SRAM.scala 148:25:@62964.4]
  wire  _T_861; // @[SRAM.scala 148:15:@62965.4]
  wire  _T_862; // @[SRAM.scala 149:15:@62967.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@62966.4]
  reg  regs_20; // @[SRAM.scala 145:20:@62973.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@62974.4]
  wire  _T_869; // @[SRAM.scala 148:25:@62975.4]
  wire  _T_870; // @[SRAM.scala 148:15:@62976.4]
  wire  _T_871; // @[SRAM.scala 149:15:@62978.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@62977.4]
  reg  regs_21; // @[SRAM.scala 145:20:@62984.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@62985.4]
  wire  _T_878; // @[SRAM.scala 148:25:@62986.4]
  wire  _T_879; // @[SRAM.scala 148:15:@62987.4]
  wire  _T_880; // @[SRAM.scala 149:15:@62989.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@62988.4]
  reg  regs_22; // @[SRAM.scala 145:20:@62995.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@62996.4]
  wire  _T_887; // @[SRAM.scala 148:25:@62997.4]
  wire  _T_888; // @[SRAM.scala 148:15:@62998.4]
  wire  _T_889; // @[SRAM.scala 149:15:@63000.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@62999.4]
  reg  regs_23; // @[SRAM.scala 145:20:@63006.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@63007.4]
  wire  _T_896; // @[SRAM.scala 148:25:@63008.4]
  wire  _T_897; // @[SRAM.scala 148:15:@63009.4]
  wire  _T_898; // @[SRAM.scala 149:15:@63011.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@63010.4]
  reg  regs_24; // @[SRAM.scala 145:20:@63017.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@63018.4]
  wire  _T_905; // @[SRAM.scala 148:25:@63019.4]
  wire  _T_906; // @[SRAM.scala 148:15:@63020.4]
  wire  _T_907; // @[SRAM.scala 149:15:@63022.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@63021.4]
  reg  regs_25; // @[SRAM.scala 145:20:@63028.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@63029.4]
  wire  _T_914; // @[SRAM.scala 148:25:@63030.4]
  wire  _T_915; // @[SRAM.scala 148:15:@63031.4]
  wire  _T_916; // @[SRAM.scala 149:15:@63033.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@63032.4]
  reg  regs_26; // @[SRAM.scala 145:20:@63039.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@63040.4]
  wire  _T_923; // @[SRAM.scala 148:25:@63041.4]
  wire  _T_924; // @[SRAM.scala 148:15:@63042.4]
  wire  _T_925; // @[SRAM.scala 149:15:@63044.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@63043.4]
  reg  regs_27; // @[SRAM.scala 145:20:@63050.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@63051.4]
  wire  _T_932; // @[SRAM.scala 148:25:@63052.4]
  wire  _T_933; // @[SRAM.scala 148:15:@63053.4]
  wire  _T_934; // @[SRAM.scala 149:15:@63055.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@63054.4]
  reg  regs_28; // @[SRAM.scala 145:20:@63061.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@63062.4]
  wire  _T_941; // @[SRAM.scala 148:25:@63063.4]
  wire  _T_942; // @[SRAM.scala 148:15:@63064.4]
  wire  _T_943; // @[SRAM.scala 149:15:@63066.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@63065.4]
  reg  regs_29; // @[SRAM.scala 145:20:@63072.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@63073.4]
  wire  _T_950; // @[SRAM.scala 148:25:@63074.4]
  wire  _T_951; // @[SRAM.scala 148:15:@63075.4]
  wire  _T_952; // @[SRAM.scala 149:15:@63077.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@63076.4]
  reg  regs_30; // @[SRAM.scala 145:20:@63083.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@63084.4]
  wire  _T_959; // @[SRAM.scala 148:25:@63085.4]
  wire  _T_960; // @[SRAM.scala 148:15:@63086.4]
  wire  _T_961; // @[SRAM.scala 149:15:@63088.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@63087.4]
  reg  regs_31; // @[SRAM.scala 145:20:@63094.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@63095.4]
  wire  _T_968; // @[SRAM.scala 148:25:@63096.4]
  wire  _T_969; // @[SRAM.scala 148:15:@63097.4]
  wire  _T_970; // @[SRAM.scala 149:15:@63099.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@63098.4]
  reg  regs_32; // @[SRAM.scala 145:20:@63105.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@63106.4]
  wire  _T_977; // @[SRAM.scala 148:25:@63107.4]
  wire  _T_978; // @[SRAM.scala 148:15:@63108.4]
  wire  _T_979; // @[SRAM.scala 149:15:@63110.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@63109.4]
  reg  regs_33; // @[SRAM.scala 145:20:@63116.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@63117.4]
  wire  _T_986; // @[SRAM.scala 148:25:@63118.4]
  wire  _T_987; // @[SRAM.scala 148:15:@63119.4]
  wire  _T_988; // @[SRAM.scala 149:15:@63121.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@63120.4]
  reg  regs_34; // @[SRAM.scala 145:20:@63127.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@63128.4]
  wire  _T_995; // @[SRAM.scala 148:25:@63129.4]
  wire  _T_996; // @[SRAM.scala 148:15:@63130.4]
  wire  _T_997; // @[SRAM.scala 149:15:@63132.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@63131.4]
  reg  regs_35; // @[SRAM.scala 145:20:@63138.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@63139.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@63140.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@63141.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@63143.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@63142.4]
  reg  regs_36; // @[SRAM.scala 145:20:@63149.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@63150.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@63151.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@63152.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@63154.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@63153.4]
  reg  regs_37; // @[SRAM.scala 145:20:@63160.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@63161.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@63162.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@63163.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@63165.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@63164.4]
  reg  regs_38; // @[SRAM.scala 145:20:@63171.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@63172.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@63173.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@63174.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@63176.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@63175.4]
  reg  regs_39; // @[SRAM.scala 145:20:@63182.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@63183.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@63184.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@63185.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@63187.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@63186.4]
  reg  regs_40; // @[SRAM.scala 145:20:@63193.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@63194.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@63195.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@63196.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@63198.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@63197.4]
  reg  regs_41; // @[SRAM.scala 145:20:@63204.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@63205.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@63206.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@63207.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@63209.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@63208.4]
  reg  regs_42; // @[SRAM.scala 145:20:@63215.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@63216.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@63217.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@63218.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@63220.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@63219.4]
  reg  regs_43; // @[SRAM.scala 145:20:@63226.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@63227.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@63228.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@63229.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@63231.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@63230.4]
  reg  regs_44; // @[SRAM.scala 145:20:@63237.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@63238.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@63239.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@63240.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@63242.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@63241.4]
  reg  regs_45; // @[SRAM.scala 145:20:@63248.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@63249.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@63250.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@63251.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@63253.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@63252.4]
  reg  regs_46; // @[SRAM.scala 145:20:@63259.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@63260.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@63261.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@63262.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@63264.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@63263.4]
  reg  regs_47; // @[SRAM.scala 145:20:@63270.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@63271.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@63272.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@63273.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@63275.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@63274.4]
  reg  regs_48; // @[SRAM.scala 145:20:@63281.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@63282.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@63283.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@63284.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@63286.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@63285.4]
  reg  regs_49; // @[SRAM.scala 145:20:@63292.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@63293.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@63294.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@63295.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@63297.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@63296.4]
  reg  regs_50; // @[SRAM.scala 145:20:@63303.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@63304.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@63305.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@63306.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@63308.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@63307.4]
  reg  regs_51; // @[SRAM.scala 145:20:@63314.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@63315.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@63316.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@63317.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@63319.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@63318.4]
  reg  regs_52; // @[SRAM.scala 145:20:@63325.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@63326.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@63327.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@63328.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@63330.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@63329.4]
  reg  regs_53; // @[SRAM.scala 145:20:@63336.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@63337.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@63338.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@63339.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@63341.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@63340.4]
  reg  regs_54; // @[SRAM.scala 145:20:@63347.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@63348.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@63349.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@63350.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@63352.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@63351.4]
  reg  regs_55; // @[SRAM.scala 145:20:@63358.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@63359.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@63360.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@63361.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@63363.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@63362.4]
  reg  regs_56; // @[SRAM.scala 145:20:@63369.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@63370.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@63371.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@63372.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@63374.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@63373.4]
  reg  regs_57; // @[SRAM.scala 145:20:@63380.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@63381.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@63382.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@63383.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@63385.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@63384.4]
  reg  regs_58; // @[SRAM.scala 145:20:@63391.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@63392.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@63393.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@63394.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@63396.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@63395.4]
  reg  regs_59; // @[SRAM.scala 145:20:@63402.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@63403.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@63404.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@63405.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@63407.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@63406.4]
  reg  regs_60; // @[SRAM.scala 145:20:@63413.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@63414.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@63415.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@63416.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@63418.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@63417.4]
  reg  regs_61; // @[SRAM.scala 145:20:@63424.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@63425.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@63426.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@63427.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@63429.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@63428.4]
  reg  regs_62; // @[SRAM.scala 145:20:@63435.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@63436.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@63437.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@63438.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@63440.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@63439.4]
  reg  regs_63; // @[SRAM.scala 145:20:@63446.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@63447.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@63448.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@63449.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@63451.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@63450.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@63520.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@63520.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@62754.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@62755.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@62756.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62758.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@62757.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@62765.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@62766.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@62767.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62769.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@62768.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@62776.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@62777.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@62778.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62780.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@62779.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@62787.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@62788.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@62789.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62791.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@62790.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@62798.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@62799.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@62800.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62802.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@62801.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@62809.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@62810.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@62811.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62813.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@62812.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@62820.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@62821.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@62822.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62824.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@62823.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@62831.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@62832.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@62833.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62835.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@62834.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@62842.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@62843.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@62844.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62846.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@62845.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@62853.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@62854.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@62855.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62857.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@62856.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@62864.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@62865.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@62866.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62868.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@62867.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@62875.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@62876.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@62877.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62879.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@62878.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@62886.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@62887.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@62888.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62890.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@62889.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@62897.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@62898.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@62899.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62901.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@62900.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@62908.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@62909.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@62910.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62912.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@62911.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@62919.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@62920.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@62921.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62923.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@62922.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@62930.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@62931.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@62932.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62934.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@62933.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@62941.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@62942.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@62943.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62945.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@62944.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@62952.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@62953.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@62954.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62956.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@62955.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@62963.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@62964.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@62965.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62967.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@62966.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@62974.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@62975.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@62976.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62978.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@62977.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@62985.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@62986.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@62987.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62989.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@62988.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@62996.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@62997.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@62998.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63000.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@62999.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@63007.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@63008.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@63009.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63011.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@63010.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@63018.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@63019.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@63020.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63022.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@63021.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@63029.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@63030.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@63031.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63033.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@63032.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@63040.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@63041.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@63042.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63044.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@63043.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@63051.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@63052.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@63053.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63055.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@63054.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@63062.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@63063.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@63064.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63066.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@63065.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@63073.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@63074.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@63075.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63077.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@63076.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@63084.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@63085.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@63086.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63088.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@63087.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@63095.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@63096.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@63097.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63099.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@63098.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@63106.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@63107.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@63108.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63110.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@63109.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@63117.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@63118.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@63119.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63121.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@63120.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@63128.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@63129.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@63130.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63132.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@63131.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@63139.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@63140.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@63141.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63143.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@63142.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@63150.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@63151.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@63152.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63154.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@63153.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@63161.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@63162.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@63163.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63165.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@63164.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@63172.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@63173.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@63174.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63176.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@63175.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@63183.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@63184.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@63185.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63187.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@63186.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@63194.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@63195.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@63196.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63198.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@63197.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@63205.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@63206.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@63207.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63209.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@63208.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@63216.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@63217.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@63218.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63220.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@63219.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@63227.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@63228.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@63229.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63231.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@63230.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@63238.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@63239.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@63240.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63242.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@63241.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@63249.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@63250.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@63251.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63253.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@63252.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@63260.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@63261.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@63262.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63264.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@63263.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@63271.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@63272.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@63273.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63275.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@63274.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@63282.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@63283.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@63284.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63286.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@63285.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@63293.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@63294.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@63295.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63297.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@63296.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@63304.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@63305.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@63306.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63308.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@63307.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@63315.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@63316.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@63317.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63319.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@63318.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@63326.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@63327.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@63328.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63330.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@63329.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@63337.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@63338.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@63339.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63341.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@63340.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@63348.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@63349.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@63350.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63352.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@63351.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@63359.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@63360.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@63361.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63363.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@63362.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@63370.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@63371.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@63372.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63374.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@63373.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@63381.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@63382.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@63383.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63385.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@63384.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@63392.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@63393.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@63394.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63396.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@63395.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@63403.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@63404.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@63405.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63407.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@63406.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@63414.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@63415.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@63416.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63418.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@63417.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@63425.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@63426.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@63427.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63429.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@63428.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@63436.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@63437.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@63438.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63440.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@63439.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@63447.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@63448.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@63449.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@63451.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@63450.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@63520.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@63520.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@63520.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@63522.2]
  input   clock, // @[:@63523.4]
  input   reset, // @[:@63524.4]
  output  io_in_ready, // @[:@63525.4]
  input   io_in_valid, // @[:@63525.4]
  input   io_in_bits, // @[:@63525.4]
  input   io_out_ready, // @[:@63525.4]
  output  io_out_valid, // @[:@63525.4]
  output  io_out_bits, // @[:@63525.4]
  input   io_banks_0_wdata_valid, // @[:@63525.4]
  input   io_banks_0_wdata_bits, // @[:@63525.4]
  input   io_banks_1_wdata_valid, // @[:@63525.4]
  input   io_banks_1_wdata_bits, // @[:@63525.4]
  input   io_banks_2_wdata_valid, // @[:@63525.4]
  input   io_banks_2_wdata_bits, // @[:@63525.4]
  input   io_banks_3_wdata_valid, // @[:@63525.4]
  input   io_banks_3_wdata_bits, // @[:@63525.4]
  input   io_banks_4_wdata_valid, // @[:@63525.4]
  input   io_banks_4_wdata_bits, // @[:@63525.4]
  input   io_banks_5_wdata_valid, // @[:@63525.4]
  input   io_banks_5_wdata_bits, // @[:@63525.4]
  input   io_banks_6_wdata_valid, // @[:@63525.4]
  input   io_banks_6_wdata_bits, // @[:@63525.4]
  input   io_banks_7_wdata_valid, // @[:@63525.4]
  input   io_banks_7_wdata_bits, // @[:@63525.4]
  input   io_banks_8_wdata_valid, // @[:@63525.4]
  input   io_banks_8_wdata_bits, // @[:@63525.4]
  input   io_banks_9_wdata_valid, // @[:@63525.4]
  input   io_banks_9_wdata_bits, // @[:@63525.4]
  input   io_banks_10_wdata_valid, // @[:@63525.4]
  input   io_banks_10_wdata_bits, // @[:@63525.4]
  input   io_banks_11_wdata_valid, // @[:@63525.4]
  input   io_banks_11_wdata_bits, // @[:@63525.4]
  input   io_banks_12_wdata_valid, // @[:@63525.4]
  input   io_banks_12_wdata_bits, // @[:@63525.4]
  input   io_banks_13_wdata_valid, // @[:@63525.4]
  input   io_banks_13_wdata_bits, // @[:@63525.4]
  input   io_banks_14_wdata_valid, // @[:@63525.4]
  input   io_banks_14_wdata_bits, // @[:@63525.4]
  input   io_banks_15_wdata_valid, // @[:@63525.4]
  input   io_banks_15_wdata_bits, // @[:@63525.4]
  input   io_banks_16_wdata_valid, // @[:@63525.4]
  input   io_banks_16_wdata_bits, // @[:@63525.4]
  input   io_banks_17_wdata_valid, // @[:@63525.4]
  input   io_banks_17_wdata_bits, // @[:@63525.4]
  input   io_banks_18_wdata_valid, // @[:@63525.4]
  input   io_banks_18_wdata_bits, // @[:@63525.4]
  input   io_banks_19_wdata_valid, // @[:@63525.4]
  input   io_banks_19_wdata_bits, // @[:@63525.4]
  input   io_banks_20_wdata_valid, // @[:@63525.4]
  input   io_banks_20_wdata_bits, // @[:@63525.4]
  input   io_banks_21_wdata_valid, // @[:@63525.4]
  input   io_banks_21_wdata_bits, // @[:@63525.4]
  input   io_banks_22_wdata_valid, // @[:@63525.4]
  input   io_banks_22_wdata_bits, // @[:@63525.4]
  input   io_banks_23_wdata_valid, // @[:@63525.4]
  input   io_banks_23_wdata_bits, // @[:@63525.4]
  input   io_banks_24_wdata_valid, // @[:@63525.4]
  input   io_banks_24_wdata_bits, // @[:@63525.4]
  input   io_banks_25_wdata_valid, // @[:@63525.4]
  input   io_banks_25_wdata_bits, // @[:@63525.4]
  input   io_banks_26_wdata_valid, // @[:@63525.4]
  input   io_banks_26_wdata_bits, // @[:@63525.4]
  input   io_banks_27_wdata_valid, // @[:@63525.4]
  input   io_banks_27_wdata_bits, // @[:@63525.4]
  input   io_banks_28_wdata_valid, // @[:@63525.4]
  input   io_banks_28_wdata_bits, // @[:@63525.4]
  input   io_banks_29_wdata_valid, // @[:@63525.4]
  input   io_banks_29_wdata_bits, // @[:@63525.4]
  input   io_banks_30_wdata_valid, // @[:@63525.4]
  input   io_banks_30_wdata_bits, // @[:@63525.4]
  input   io_banks_31_wdata_valid, // @[:@63525.4]
  input   io_banks_31_wdata_bits, // @[:@63525.4]
  input   io_banks_32_wdata_valid, // @[:@63525.4]
  input   io_banks_32_wdata_bits, // @[:@63525.4]
  input   io_banks_33_wdata_valid, // @[:@63525.4]
  input   io_banks_33_wdata_bits, // @[:@63525.4]
  input   io_banks_34_wdata_valid, // @[:@63525.4]
  input   io_banks_34_wdata_bits, // @[:@63525.4]
  input   io_banks_35_wdata_valid, // @[:@63525.4]
  input   io_banks_35_wdata_bits, // @[:@63525.4]
  input   io_banks_36_wdata_valid, // @[:@63525.4]
  input   io_banks_36_wdata_bits, // @[:@63525.4]
  input   io_banks_37_wdata_valid, // @[:@63525.4]
  input   io_banks_37_wdata_bits, // @[:@63525.4]
  input   io_banks_38_wdata_valid, // @[:@63525.4]
  input   io_banks_38_wdata_bits, // @[:@63525.4]
  input   io_banks_39_wdata_valid, // @[:@63525.4]
  input   io_banks_39_wdata_bits, // @[:@63525.4]
  input   io_banks_40_wdata_valid, // @[:@63525.4]
  input   io_banks_40_wdata_bits, // @[:@63525.4]
  input   io_banks_41_wdata_valid, // @[:@63525.4]
  input   io_banks_41_wdata_bits, // @[:@63525.4]
  input   io_banks_42_wdata_valid, // @[:@63525.4]
  input   io_banks_42_wdata_bits, // @[:@63525.4]
  input   io_banks_43_wdata_valid, // @[:@63525.4]
  input   io_banks_43_wdata_bits, // @[:@63525.4]
  input   io_banks_44_wdata_valid, // @[:@63525.4]
  input   io_banks_44_wdata_bits, // @[:@63525.4]
  input   io_banks_45_wdata_valid, // @[:@63525.4]
  input   io_banks_45_wdata_bits, // @[:@63525.4]
  input   io_banks_46_wdata_valid, // @[:@63525.4]
  input   io_banks_46_wdata_bits, // @[:@63525.4]
  input   io_banks_47_wdata_valid, // @[:@63525.4]
  input   io_banks_47_wdata_bits, // @[:@63525.4]
  input   io_banks_48_wdata_valid, // @[:@63525.4]
  input   io_banks_48_wdata_bits, // @[:@63525.4]
  input   io_banks_49_wdata_valid, // @[:@63525.4]
  input   io_banks_49_wdata_bits, // @[:@63525.4]
  input   io_banks_50_wdata_valid, // @[:@63525.4]
  input   io_banks_50_wdata_bits, // @[:@63525.4]
  input   io_banks_51_wdata_valid, // @[:@63525.4]
  input   io_banks_51_wdata_bits, // @[:@63525.4]
  input   io_banks_52_wdata_valid, // @[:@63525.4]
  input   io_banks_52_wdata_bits, // @[:@63525.4]
  input   io_banks_53_wdata_valid, // @[:@63525.4]
  input   io_banks_53_wdata_bits, // @[:@63525.4]
  input   io_banks_54_wdata_valid, // @[:@63525.4]
  input   io_banks_54_wdata_bits, // @[:@63525.4]
  input   io_banks_55_wdata_valid, // @[:@63525.4]
  input   io_banks_55_wdata_bits, // @[:@63525.4]
  input   io_banks_56_wdata_valid, // @[:@63525.4]
  input   io_banks_56_wdata_bits, // @[:@63525.4]
  input   io_banks_57_wdata_valid, // @[:@63525.4]
  input   io_banks_57_wdata_bits, // @[:@63525.4]
  input   io_banks_58_wdata_valid, // @[:@63525.4]
  input   io_banks_58_wdata_bits, // @[:@63525.4]
  input   io_banks_59_wdata_valid, // @[:@63525.4]
  input   io_banks_59_wdata_bits, // @[:@63525.4]
  input   io_banks_60_wdata_valid, // @[:@63525.4]
  input   io_banks_60_wdata_bits, // @[:@63525.4]
  input   io_banks_61_wdata_valid, // @[:@63525.4]
  input   io_banks_61_wdata_bits, // @[:@63525.4]
  input   io_banks_62_wdata_valid, // @[:@63525.4]
  input   io_banks_62_wdata_bits, // @[:@63525.4]
  input   io_banks_63_wdata_valid, // @[:@63525.4]
  input   io_banks_63_wdata_bits // @[:@63525.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@63791.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@63791.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@63791.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@63791.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@63791.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@63801.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@63801.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@63801.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@63801.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@63801.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@63816.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@63816.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@63816.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@63816.4]
  wire  writeEn; // @[FIFO.scala 30:29:@63789.4]
  wire  readEn; // @[FIFO.scala 31:29:@63790.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@63811.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@63812.4]
  wire  _T_824; // @[FIFO.scala 45:27:@63813.4]
  wire  empty; // @[FIFO.scala 45:24:@63814.4]
  wire  full; // @[FIFO.scala 46:23:@63815.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@64982.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@64983.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@63791.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@63801.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@63816.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@63789.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@63790.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@63812.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@63813.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@63814.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@63815.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@64982.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@64983.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@64989.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@64987.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@64021.4]
  assign enqCounter_clock = clock; // @[:@63792.4]
  assign enqCounter_reset = reset; // @[:@63793.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@63799.4]
  assign deqCounter_clock = clock; // @[:@63802.4]
  assign deqCounter_reset = reset; // @[:@63803.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@63809.4]
  assign FFRAM_clock = clock; // @[:@63817.4]
  assign FFRAM_reset = reset; // @[:@63818.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@64017.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@64018.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@64019.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@64020.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@64023.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@64022.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@64026.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@64025.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@64029.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@64028.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@64032.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@64031.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@64035.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@64034.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@64038.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@64037.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@64041.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@64040.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@64044.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@64043.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@64047.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@64046.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@64050.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@64049.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@64053.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@64052.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@64056.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@64055.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@64059.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@64058.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@64062.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@64061.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@64065.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@64064.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@64068.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@64067.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@64071.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@64070.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@64074.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@64073.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@64077.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@64076.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@64080.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@64079.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@64083.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@64082.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@64086.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@64085.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@64089.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@64088.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@64092.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@64091.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@64095.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@64094.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@64098.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@64097.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@64101.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@64100.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@64104.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@64103.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@64107.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@64106.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@64110.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@64109.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@64113.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@64112.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@64116.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@64115.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@64119.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@64118.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@64122.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@64121.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@64125.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@64124.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@64128.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@64127.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@64131.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@64130.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@64134.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@64133.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@64137.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@64136.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@64140.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@64139.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@64143.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@64142.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@64146.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@64145.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@64149.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@64148.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@64152.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@64151.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@64155.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@64154.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@64158.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@64157.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@64161.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@64160.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@64164.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@64163.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@64167.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@64166.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@64170.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@64169.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@64173.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@64172.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@64176.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@64175.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@64179.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@64178.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@64182.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@64181.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@64185.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@64184.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@64188.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@64187.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@64191.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@64190.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@64194.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@64193.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@64197.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@64196.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@64200.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@64199.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@64203.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@64202.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@64206.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@64205.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@64209.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@64208.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@64212.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@64211.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@64991.2]
  input         clock, // @[:@64992.4]
  input         reset, // @[:@64993.4]
  input         io_dram_cmd_ready, // @[:@64994.4]
  output        io_dram_cmd_valid, // @[:@64994.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@64994.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@64994.4]
  input         io_dram_wdata_ready, // @[:@64994.4]
  output        io_dram_wdata_valid, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@64994.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@64994.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@64994.4]
  output        io_dram_wresp_ready, // @[:@64994.4]
  input         io_dram_wresp_valid, // @[:@64994.4]
  output        io_store_cmd_ready, // @[:@64994.4]
  input         io_store_cmd_valid, // @[:@64994.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@64994.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@64994.4]
  output        io_store_data_ready, // @[:@64994.4]
  input         io_store_data_valid, // @[:@64994.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@64994.4]
  input         io_store_data_bits_wstrb, // @[:@64994.4]
  input         io_store_wresp_ready, // @[:@64994.4]
  output        io_store_wresp_valid, // @[:@64994.4]
  output        io_store_wresp_bits // @[:@64994.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@65119.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@65119.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@65119.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@65119.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@65119.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@65119.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@65119.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@65119.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@65119.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@65119.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@65525.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@65525.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@65525.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@65525.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@65525.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@65525.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@65525.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@65525.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@65525.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@65766.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@65766.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@65522.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@65119.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@65525.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@65766.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@65522.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@65519.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@65520.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@65523.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@65555.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@65556.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@65557.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@65558.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@65559.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@65560.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@65561.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@65562.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@65563.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@65564.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@65565.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@65566.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@65567.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@65568.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@65569.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@65570.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@65571.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@65701.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@65702.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@65703.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@65704.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@65705.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@65706.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@65707.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@65708.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@65709.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@65710.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@65711.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@65712.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@65713.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@65714.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@65715.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@65716.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@65717.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@65718.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@65719.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@65720.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@65721.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@65722.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@65723.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@65724.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@65725.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@65726.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@65727.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@65728.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@65729.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@65730.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@65731.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@65732.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@65733.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@65734.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@65735.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@65736.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@65737.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@65738.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@65739.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@65740.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@65741.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@65742.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@65743.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@65744.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@65745.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@65746.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@65747.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@65748.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@65749.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@65750.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@65751.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@65752.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@65753.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@65754.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@65755.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@65756.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@65757.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@65758.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@65759.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@65760.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@65761.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@65762.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@65763.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@65764.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@66033.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@65517.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@65554.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@66034.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@66035.4]
  assign cmd_clock = clock; // @[:@65120.4]
  assign cmd_reset = reset; // @[:@65121.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@65514.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@65516.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@65515.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@65518.4]
  assign wdata_clock = clock; // @[:@65526.4]
  assign wdata_reset = reset; // @[:@65527.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@65551.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@65552.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@65553.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@65765.4]
  assign wresp_clock = clock; // @[:@65767.4]
  assign wresp_reset = reset; // @[:@65768.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@66031.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@66032.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@66036.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@66102.2]
  output        io_in_ready, // @[:@66105.4]
  input         io_in_valid, // @[:@66105.4]
  input  [63:0] io_in_bits_0_addr, // @[:@66105.4]
  input  [31:0] io_in_bits_0_size, // @[:@66105.4]
  input         io_in_bits_0_isWr, // @[:@66105.4]
  input  [31:0] io_in_bits_0_tag, // @[:@66105.4]
  input         io_out_ready, // @[:@66105.4]
  output        io_out_valid, // @[:@66105.4]
  output [63:0] io_out_bits_addr, // @[:@66105.4]
  output [31:0] io_out_bits_size, // @[:@66105.4]
  output        io_out_bits_isWr, // @[:@66105.4]
  output [31:0] io_out_bits_tag // @[:@66105.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@66107.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@66107.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@66116.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@66115.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@66121.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@66120.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@66118.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@66117.4]
endmodule
module MuxPipe_1( // @[:@66123.2]
  output        io_in_ready, // @[:@66126.4]
  input         io_in_valid, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@66126.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@66126.4]
  input         io_in_bits_0_wstrb_0, // @[:@66126.4]
  input         io_in_bits_0_wstrb_1, // @[:@66126.4]
  input         io_in_bits_0_wstrb_2, // @[:@66126.4]
  input         io_in_bits_0_wstrb_3, // @[:@66126.4]
  input         io_in_bits_0_wstrb_4, // @[:@66126.4]
  input         io_in_bits_0_wstrb_5, // @[:@66126.4]
  input         io_in_bits_0_wstrb_6, // @[:@66126.4]
  input         io_in_bits_0_wstrb_7, // @[:@66126.4]
  input         io_in_bits_0_wstrb_8, // @[:@66126.4]
  input         io_in_bits_0_wstrb_9, // @[:@66126.4]
  input         io_in_bits_0_wstrb_10, // @[:@66126.4]
  input         io_in_bits_0_wstrb_11, // @[:@66126.4]
  input         io_in_bits_0_wstrb_12, // @[:@66126.4]
  input         io_in_bits_0_wstrb_13, // @[:@66126.4]
  input         io_in_bits_0_wstrb_14, // @[:@66126.4]
  input         io_in_bits_0_wstrb_15, // @[:@66126.4]
  input         io_in_bits_0_wstrb_16, // @[:@66126.4]
  input         io_in_bits_0_wstrb_17, // @[:@66126.4]
  input         io_in_bits_0_wstrb_18, // @[:@66126.4]
  input         io_in_bits_0_wstrb_19, // @[:@66126.4]
  input         io_in_bits_0_wstrb_20, // @[:@66126.4]
  input         io_in_bits_0_wstrb_21, // @[:@66126.4]
  input         io_in_bits_0_wstrb_22, // @[:@66126.4]
  input         io_in_bits_0_wstrb_23, // @[:@66126.4]
  input         io_in_bits_0_wstrb_24, // @[:@66126.4]
  input         io_in_bits_0_wstrb_25, // @[:@66126.4]
  input         io_in_bits_0_wstrb_26, // @[:@66126.4]
  input         io_in_bits_0_wstrb_27, // @[:@66126.4]
  input         io_in_bits_0_wstrb_28, // @[:@66126.4]
  input         io_in_bits_0_wstrb_29, // @[:@66126.4]
  input         io_in_bits_0_wstrb_30, // @[:@66126.4]
  input         io_in_bits_0_wstrb_31, // @[:@66126.4]
  input         io_in_bits_0_wstrb_32, // @[:@66126.4]
  input         io_in_bits_0_wstrb_33, // @[:@66126.4]
  input         io_in_bits_0_wstrb_34, // @[:@66126.4]
  input         io_in_bits_0_wstrb_35, // @[:@66126.4]
  input         io_in_bits_0_wstrb_36, // @[:@66126.4]
  input         io_in_bits_0_wstrb_37, // @[:@66126.4]
  input         io_in_bits_0_wstrb_38, // @[:@66126.4]
  input         io_in_bits_0_wstrb_39, // @[:@66126.4]
  input         io_in_bits_0_wstrb_40, // @[:@66126.4]
  input         io_in_bits_0_wstrb_41, // @[:@66126.4]
  input         io_in_bits_0_wstrb_42, // @[:@66126.4]
  input         io_in_bits_0_wstrb_43, // @[:@66126.4]
  input         io_in_bits_0_wstrb_44, // @[:@66126.4]
  input         io_in_bits_0_wstrb_45, // @[:@66126.4]
  input         io_in_bits_0_wstrb_46, // @[:@66126.4]
  input         io_in_bits_0_wstrb_47, // @[:@66126.4]
  input         io_in_bits_0_wstrb_48, // @[:@66126.4]
  input         io_in_bits_0_wstrb_49, // @[:@66126.4]
  input         io_in_bits_0_wstrb_50, // @[:@66126.4]
  input         io_in_bits_0_wstrb_51, // @[:@66126.4]
  input         io_in_bits_0_wstrb_52, // @[:@66126.4]
  input         io_in_bits_0_wstrb_53, // @[:@66126.4]
  input         io_in_bits_0_wstrb_54, // @[:@66126.4]
  input         io_in_bits_0_wstrb_55, // @[:@66126.4]
  input         io_in_bits_0_wstrb_56, // @[:@66126.4]
  input         io_in_bits_0_wstrb_57, // @[:@66126.4]
  input         io_in_bits_0_wstrb_58, // @[:@66126.4]
  input         io_in_bits_0_wstrb_59, // @[:@66126.4]
  input         io_in_bits_0_wstrb_60, // @[:@66126.4]
  input         io_in_bits_0_wstrb_61, // @[:@66126.4]
  input         io_in_bits_0_wstrb_62, // @[:@66126.4]
  input         io_in_bits_0_wstrb_63, // @[:@66126.4]
  input         io_out_ready, // @[:@66126.4]
  output        io_out_valid, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_0, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_1, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_2, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_3, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_4, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_5, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_6, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_7, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_8, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_9, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_10, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_11, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_12, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_13, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_14, // @[:@66126.4]
  output [31:0] io_out_bits_wdata_15, // @[:@66126.4]
  output        io_out_bits_wstrb_0, // @[:@66126.4]
  output        io_out_bits_wstrb_1, // @[:@66126.4]
  output        io_out_bits_wstrb_2, // @[:@66126.4]
  output        io_out_bits_wstrb_3, // @[:@66126.4]
  output        io_out_bits_wstrb_4, // @[:@66126.4]
  output        io_out_bits_wstrb_5, // @[:@66126.4]
  output        io_out_bits_wstrb_6, // @[:@66126.4]
  output        io_out_bits_wstrb_7, // @[:@66126.4]
  output        io_out_bits_wstrb_8, // @[:@66126.4]
  output        io_out_bits_wstrb_9, // @[:@66126.4]
  output        io_out_bits_wstrb_10, // @[:@66126.4]
  output        io_out_bits_wstrb_11, // @[:@66126.4]
  output        io_out_bits_wstrb_12, // @[:@66126.4]
  output        io_out_bits_wstrb_13, // @[:@66126.4]
  output        io_out_bits_wstrb_14, // @[:@66126.4]
  output        io_out_bits_wstrb_15, // @[:@66126.4]
  output        io_out_bits_wstrb_16, // @[:@66126.4]
  output        io_out_bits_wstrb_17, // @[:@66126.4]
  output        io_out_bits_wstrb_18, // @[:@66126.4]
  output        io_out_bits_wstrb_19, // @[:@66126.4]
  output        io_out_bits_wstrb_20, // @[:@66126.4]
  output        io_out_bits_wstrb_21, // @[:@66126.4]
  output        io_out_bits_wstrb_22, // @[:@66126.4]
  output        io_out_bits_wstrb_23, // @[:@66126.4]
  output        io_out_bits_wstrb_24, // @[:@66126.4]
  output        io_out_bits_wstrb_25, // @[:@66126.4]
  output        io_out_bits_wstrb_26, // @[:@66126.4]
  output        io_out_bits_wstrb_27, // @[:@66126.4]
  output        io_out_bits_wstrb_28, // @[:@66126.4]
  output        io_out_bits_wstrb_29, // @[:@66126.4]
  output        io_out_bits_wstrb_30, // @[:@66126.4]
  output        io_out_bits_wstrb_31, // @[:@66126.4]
  output        io_out_bits_wstrb_32, // @[:@66126.4]
  output        io_out_bits_wstrb_33, // @[:@66126.4]
  output        io_out_bits_wstrb_34, // @[:@66126.4]
  output        io_out_bits_wstrb_35, // @[:@66126.4]
  output        io_out_bits_wstrb_36, // @[:@66126.4]
  output        io_out_bits_wstrb_37, // @[:@66126.4]
  output        io_out_bits_wstrb_38, // @[:@66126.4]
  output        io_out_bits_wstrb_39, // @[:@66126.4]
  output        io_out_bits_wstrb_40, // @[:@66126.4]
  output        io_out_bits_wstrb_41, // @[:@66126.4]
  output        io_out_bits_wstrb_42, // @[:@66126.4]
  output        io_out_bits_wstrb_43, // @[:@66126.4]
  output        io_out_bits_wstrb_44, // @[:@66126.4]
  output        io_out_bits_wstrb_45, // @[:@66126.4]
  output        io_out_bits_wstrb_46, // @[:@66126.4]
  output        io_out_bits_wstrb_47, // @[:@66126.4]
  output        io_out_bits_wstrb_48, // @[:@66126.4]
  output        io_out_bits_wstrb_49, // @[:@66126.4]
  output        io_out_bits_wstrb_50, // @[:@66126.4]
  output        io_out_bits_wstrb_51, // @[:@66126.4]
  output        io_out_bits_wstrb_52, // @[:@66126.4]
  output        io_out_bits_wstrb_53, // @[:@66126.4]
  output        io_out_bits_wstrb_54, // @[:@66126.4]
  output        io_out_bits_wstrb_55, // @[:@66126.4]
  output        io_out_bits_wstrb_56, // @[:@66126.4]
  output        io_out_bits_wstrb_57, // @[:@66126.4]
  output        io_out_bits_wstrb_58, // @[:@66126.4]
  output        io_out_bits_wstrb_59, // @[:@66126.4]
  output        io_out_bits_wstrb_60, // @[:@66126.4]
  output        io_out_bits_wstrb_61, // @[:@66126.4]
  output        io_out_bits_wstrb_62, // @[:@66126.4]
  output        io_out_bits_wstrb_63 // @[:@66126.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@66128.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@66128.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@66213.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@66212.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@66279.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@66280.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@66281.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@66282.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@66283.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@66284.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@66285.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@66286.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@66287.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@66288.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@66289.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@66290.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@66291.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@66292.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@66293.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@66294.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@66215.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@66216.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@66217.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@66218.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@66219.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@66220.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@66221.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@66222.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@66223.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@66224.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@66225.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@66226.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@66227.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@66228.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@66229.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@66230.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@66231.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@66232.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@66233.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@66234.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@66235.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@66236.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@66237.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@66238.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@66239.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@66240.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@66241.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@66242.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@66243.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@66244.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@66245.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@66246.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@66247.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@66248.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@66249.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@66250.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@66251.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@66252.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@66253.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@66254.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@66255.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@66256.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@66257.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@66258.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@66259.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@66260.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@66261.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@66262.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@66263.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@66264.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@66265.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@66266.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@66267.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@66268.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@66269.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@66270.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@66271.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@66272.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@66273.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@66274.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@66275.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@66276.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@66277.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@66278.4]
endmodule
module ElementCounter( // @[:@66296.2]
  input         clock, // @[:@66297.4]
  input         reset, // @[:@66298.4]
  input         io_reset, // @[:@66299.4]
  input         io_enable, // @[:@66299.4]
  output [31:0] io_out // @[:@66299.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@66301.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@66302.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@66303.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@66308.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@66304.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@66302.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@66303.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@66308.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@66304.4]
  assign io_out = count; // @[Counter.scala 47:10:@66311.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@66313.2]
  input         clock, // @[:@66314.4]
  input         reset, // @[:@66315.4]
  output        io_app_0_cmd_ready, // @[:@66316.4]
  input         io_app_0_cmd_valid, // @[:@66316.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@66316.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@66316.4]
  input         io_app_0_cmd_bits_isWr, // @[:@66316.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@66316.4]
  output        io_app_0_wdata_ready, // @[:@66316.4]
  input         io_app_0_wdata_valid, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@66316.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@66316.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@66316.4]
  input         io_app_0_rresp_ready, // @[:@66316.4]
  input         io_app_0_wresp_ready, // @[:@66316.4]
  output        io_app_0_wresp_valid, // @[:@66316.4]
  input         io_dram_cmd_ready, // @[:@66316.4]
  output        io_dram_cmd_valid, // @[:@66316.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@66316.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@66316.4]
  output        io_dram_cmd_bits_isWr, // @[:@66316.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@66316.4]
  input         io_dram_wdata_ready, // @[:@66316.4]
  output        io_dram_wdata_valid, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@66316.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@66316.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@66316.4]
  output        io_dram_rresp_ready, // @[:@66316.4]
  output        io_dram_wresp_ready, // @[:@66316.4]
  input         io_dram_wresp_valid, // @[:@66316.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@66316.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@66545.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@66545.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@66545.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@66545.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@66545.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@66552.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@66552.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@66552.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@66552.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@66552.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@66562.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@66562.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@66562.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@66562.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@66562.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@66562.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@66562.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@66562.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@66562.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@66562.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@66562.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@66562.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@66585.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@66585.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@66588.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@66588.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@66588.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@66588.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@66588.4]
  wire  _T_346; // @[package.scala 96:25:@66557.4 package.scala 96:25:@66558.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@66559.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@66561.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@66577.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@66579.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@66582.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@66591.4]
  wire [31:0] _T_365; // @[:@66595.4 :@66596.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@66597.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@66603.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@66606.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@66607.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@66794.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@66801.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@66806.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@66810.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@66811.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@66835.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@66545.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@66552.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@66562.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@66585.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@66588.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@66557.4 package.scala 96:25:@66558.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@66559.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@66561.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@66577.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@66579.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@66582.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@66591.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@66595.4 :@66596.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@66597.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@66603.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@66606.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@66607.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@66794.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@66801.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@66806.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@66810.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@66811.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@66835.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@66808.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@66814.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@66837.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@66697.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@66696.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@66695.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@66693.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@66692.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@66780.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@66764.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@66765.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@66766.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@66767.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@66768.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@66769.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@66770.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@66771.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@66772.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@66773.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@66774.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@66775.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@66776.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@66777.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@66778.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@66779.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@66700.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@66701.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@66702.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@66703.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@66704.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@66705.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@66706.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@66707.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@66708.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@66709.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@66710.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@66711.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@66712.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@66713.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@66714.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@66715.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@66716.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@66717.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@66718.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@66719.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@66720.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@66721.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@66722.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@66723.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@66724.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@66725.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@66726.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@66727.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@66728.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@66729.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@66730.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@66731.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@66732.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@66733.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@66734.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@66735.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@66736.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@66737.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@66738.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@66739.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@66740.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@66741.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@66742.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@66743.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@66744.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@66745.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@66746.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@66747.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@66748.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@66749.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@66750.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@66751.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@66752.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@66753.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@66754.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@66755.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@66756.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@66757.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@66758.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@66759.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@66760.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@66761.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@66762.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@66763.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@66841.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@66844.4]
  assign RetimeWrapper_clock = clock; // @[:@66546.4]
  assign RetimeWrapper_reset = reset; // @[:@66547.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@66549.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@66548.4]
  assign RetimeWrapper_1_clock = clock; // @[:@66553.4]
  assign RetimeWrapper_1_reset = reset; // @[:@66554.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@66556.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@66555.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@66565.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@66571.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@66570.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@66568.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@66567.4 FringeBundles.scala 115:32:@66584.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@66698.4 StreamArbiter.scala 57:23:@66804.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@66609.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@66676.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@66677.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@66678.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@66679.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@66680.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@66681.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@66682.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@66683.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@66684.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@66685.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@66686.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@66687.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@66688.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@66689.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@66690.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@66691.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@66612.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@66613.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@66614.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@66615.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@66616.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@66617.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@66618.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@66619.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@66620.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@66621.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@66622.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@66623.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@66624.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@66625.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@66626.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@66627.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@66628.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@66629.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@66630.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@66631.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@66632.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@66633.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@66634.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@66635.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@66636.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@66637.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@66638.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@66639.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@66640.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@66641.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@66642.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@66643.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@66644.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@66645.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@66646.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@66647.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@66648.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@66649.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@66650.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@66651.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@66652.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@66653.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@66654.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@66655.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@66656.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@66657.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@66658.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@66659.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@66660.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@66661.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@66662.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@66663.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@66664.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@66665.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@66666.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@66667.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@66668.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@66669.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@66670.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@66671.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@66672.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@66673.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@66674.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@66675.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@66781.4 StreamArbiter.scala 58:25:@66805.4]
  assign elementCtr_clock = clock; // @[:@66589.4]
  assign elementCtr_reset = reset; // @[:@66590.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@66593.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@66592.4]
endmodule
module Counter_72( // @[:@66846.2]
  input         clock, // @[:@66847.4]
  input         reset, // @[:@66848.4]
  input         io_reset, // @[:@66849.4]
  input         io_enable, // @[:@66849.4]
  input  [31:0] io_stride, // @[:@66849.4]
  output [31:0] io_out, // @[:@66849.4]
  output [31:0] io_next // @[:@66849.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@66851.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@66852.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@66853.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@66858.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@66854.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@66852.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@66853.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@66858.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@66854.4]
  assign io_out = count; // @[Counter.scala 25:10:@66861.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@66862.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@66864.2]
  input         clock, // @[:@66865.4]
  input         reset, // @[:@66866.4]
  output        io_in_cmd_ready, // @[:@66867.4]
  input         io_in_cmd_valid, // @[:@66867.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@66867.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@66867.4]
  input         io_in_cmd_bits_isWr, // @[:@66867.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@66867.4]
  output        io_in_wdata_ready, // @[:@66867.4]
  input         io_in_wdata_valid, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@66867.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@66867.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@66867.4]
  input         io_in_rresp_ready, // @[:@66867.4]
  input         io_in_wresp_ready, // @[:@66867.4]
  output        io_in_wresp_valid, // @[:@66867.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@66867.4]
  input         io_out_cmd_ready, // @[:@66867.4]
  output        io_out_cmd_valid, // @[:@66867.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@66867.4]
  output [31:0] io_out_cmd_bits_size, // @[:@66867.4]
  output        io_out_cmd_bits_isWr, // @[:@66867.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@66867.4]
  input         io_out_wdata_ready, // @[:@66867.4]
  output        io_out_wdata_valid, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@66867.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@66867.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@66867.4]
  output        io_out_rresp_ready, // @[:@66867.4]
  output        io_out_wresp_ready, // @[:@66867.4]
  input         io_out_wresp_valid, // @[:@66867.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@66867.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@66981.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@66981.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@66981.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@66981.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@66981.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@66981.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@66981.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@66984.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@66985.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@66986.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@66987.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@66990.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@66990.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@66991.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@66991.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@66992.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@66995.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@67002.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@67006.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@67009.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@67012.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@67023.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@66981.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@66984.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@66985.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@66986.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@66987.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@66990.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@66990.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@66991.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@66991.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@66992.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@66995.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@67002.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@67006.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@67009.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@67012.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@67023.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@66980.4 AXIProtocol.scala 38:19:@67014.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@66973.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@66870.4 AXIProtocol.scala 46:21:@67028.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@66869.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@66979.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@66978.4 AXIProtocol.scala 29:24:@66997.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@66977.4 AXIProtocol.scala 25:24:@66989.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@66975.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@66974.4 FringeBundles.scala 115:32:@67011.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@66972.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@66956.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@66957.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@66958.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@66959.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@66960.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@66961.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@66962.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@66963.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@66964.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@66965.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@66966.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@66967.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@66968.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@66969.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@66970.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@66971.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@66892.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@66893.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@66894.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@66895.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@66896.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@66897.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@66898.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@66899.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@66900.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@66901.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@66902.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@66903.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@66904.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@66905.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@66906.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@66907.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@66908.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@66909.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@66910.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@66911.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@66912.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@66913.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@66914.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@66915.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@66916.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@66917.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@66918.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@66919.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@66920.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@66921.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@66922.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@66923.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@66924.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@66925.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@66926.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@66927.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@66928.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@66929.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@66930.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@66931.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@66932.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@66933.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@66934.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@66935.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@66936.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@66937.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@66938.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@66939.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@66940.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@66941.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@66942.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@66943.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@66944.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@66945.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@66946.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@66947.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@66948.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@66949.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@66950.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@66951.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@66952.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@66953.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@66954.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@66955.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@66890.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@66871.4 AXIProtocol.scala 47:22:@67030.4]
  assign cmdSizeCounter_clock = clock; // @[:@66982.4]
  assign cmdSizeCounter_reset = reset; // @[:@66983.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@67015.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@67016.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@67017.4]
endmodule
module AXICmdIssue( // @[:@67050.2]
  input         clock, // @[:@67051.4]
  input         reset, // @[:@67052.4]
  output        io_in_cmd_ready, // @[:@67053.4]
  input         io_in_cmd_valid, // @[:@67053.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@67053.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@67053.4]
  input         io_in_cmd_bits_isWr, // @[:@67053.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@67053.4]
  output        io_in_wdata_ready, // @[:@67053.4]
  input         io_in_wdata_valid, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@67053.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@67053.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@67053.4]
  input         io_in_rresp_ready, // @[:@67053.4]
  input         io_in_wresp_ready, // @[:@67053.4]
  output        io_in_wresp_valid, // @[:@67053.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@67053.4]
  input         io_out_cmd_ready, // @[:@67053.4]
  output        io_out_cmd_valid, // @[:@67053.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@67053.4]
  output [31:0] io_out_cmd_bits_size, // @[:@67053.4]
  output        io_out_cmd_bits_isWr, // @[:@67053.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@67053.4]
  input         io_out_wdata_ready, // @[:@67053.4]
  output        io_out_wdata_valid, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@67053.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@67053.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@67053.4]
  output        io_out_wdata_bits_wlast, // @[:@67053.4]
  output        io_out_rresp_ready, // @[:@67053.4]
  output        io_out_wresp_ready, // @[:@67053.4]
  input         io_out_wresp_valid, // @[:@67053.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@67053.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@67167.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@67167.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@67167.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@67167.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@67167.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@67167.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@67167.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@67170.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@67171.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@67172.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@67173.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@67174.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@67180.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@67181.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@67176.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@67190.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@67191.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@67167.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@67171.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@67172.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@67173.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@67174.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@67180.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@67181.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@67176.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@67190.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@67191.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@67166.4 AXIProtocol.scala 81:19:@67188.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@67159.4 AXIProtocol.scala 82:21:@67189.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@67056.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@67055.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@67165.4 AXIProtocol.scala 84:20:@67193.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@67164.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@67163.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@67161.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@67160.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@67158.4 AXIProtocol.scala 86:22:@67195.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@67142.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@67143.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@67144.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@67145.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@67146.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@67147.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@67148.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@67149.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@67150.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@67151.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@67152.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@67153.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@67154.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@67155.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@67156.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@67157.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@67078.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@67079.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@67080.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@67081.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@67082.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@67083.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@67084.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@67085.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@67086.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@67087.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@67088.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@67089.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@67090.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@67091.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@67092.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@67093.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@67094.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@67095.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@67096.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@67097.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@67098.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@67099.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@67100.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@67101.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@67102.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@67103.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@67104.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@67105.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@67106.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@67107.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@67108.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@67109.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@67110.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@67111.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@67112.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@67113.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@67114.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@67115.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@67116.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@67117.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@67118.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@67119.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@67120.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@67121.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@67122.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@67123.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@67124.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@67125.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@67126.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@67127.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@67128.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@67129.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@67130.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@67131.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@67132.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@67133.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@67134.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@67135.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@67136.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@67137.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@67138.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@67139.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@67140.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@67141.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@67077.4 AXIProtocol.scala 87:27:@67196.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@67076.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@67057.4]
  assign wdataCounter_clock = clock; // @[:@67168.4]
  assign wdataCounter_reset = reset; // @[:@67169.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@67184.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@67185.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@67186.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@67198.2]
  input         clock, // @[:@67199.4]
  input         reset, // @[:@67200.4]
  input         io_enable, // @[:@67201.4]
  output        io_app_stores_0_cmd_ready, // @[:@67201.4]
  input         io_app_stores_0_cmd_valid, // @[:@67201.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@67201.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@67201.4]
  output        io_app_stores_0_data_ready, // @[:@67201.4]
  input         io_app_stores_0_data_valid, // @[:@67201.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@67201.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@67201.4]
  input         io_app_stores_0_wresp_ready, // @[:@67201.4]
  output        io_app_stores_0_wresp_valid, // @[:@67201.4]
  output        io_app_stores_0_wresp_bits, // @[:@67201.4]
  input         io_dram_cmd_ready, // @[:@67201.4]
  output        io_dram_cmd_valid, // @[:@67201.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@67201.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@67201.4]
  output        io_dram_cmd_bits_isWr, // @[:@67201.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@67201.4]
  input         io_dram_wdata_ready, // @[:@67201.4]
  output        io_dram_wdata_valid, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@67201.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@67201.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@67201.4]
  output        io_dram_wdata_bits_wlast, // @[:@67201.4]
  output        io_dram_rresp_ready, // @[:@67201.4]
  output        io_dram_wresp_ready, // @[:@67201.4]
  input         io_dram_wresp_valid, // @[:@67201.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@67201.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@68087.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@68101.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@68329.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@68444.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@68444.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@68087.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@68101.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@68329.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@68444.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@68100.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@68096.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@68091.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@68090.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@68669.4 DRAMArbiter.scala 100:23:@68672.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@68668.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@68667.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@68665.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@68664.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@68662.4 DRAMArbiter.scala 101:25:@68674.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@68646.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@68647.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@68648.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@68649.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@68650.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@68651.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@68652.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@68653.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@68654.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@68655.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@68656.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@68657.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@68658.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@68659.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@68660.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@68661.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@68582.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@68583.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@68584.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@68585.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@68586.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@68587.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@68588.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@68589.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@68590.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@68591.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@68592.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@68593.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@68594.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@68595.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@68596.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@68597.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@68598.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@68599.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@68600.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@68601.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@68602.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@68603.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@68604.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@68605.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@68606.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@68607.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@68608.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@68609.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@68610.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@68611.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@68612.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@68613.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@68614.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@68615.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@68616.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@68617.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@68618.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@68619.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@68620.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@68621.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@68622.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@68623.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@68624.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@68625.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@68626.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@68627.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@68628.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@68629.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@68630.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@68631.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@68632.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@68633.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@68634.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@68635.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@68636.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@68637.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@68638.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@68639.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@68640.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@68641.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@68642.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@68643.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@68644.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@68645.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@68581.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@68580.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@68561.4]
  assign StreamControllerStore_clock = clock; // @[:@68088.4]
  assign StreamControllerStore_reset = reset; // @[:@68089.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@68216.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@68209.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@68106.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@68099.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@68098.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@68097.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@68095.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@68094.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@68093.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@68092.4]
  assign StreamArbiter_clock = clock; // @[:@68102.4]
  assign StreamArbiter_reset = reset; // @[:@68103.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@68327.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@68326.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@68325.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@68323.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@68322.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@68320.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@68304.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@68305.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@68306.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@68307.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@68308.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@68309.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@68310.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@68311.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@68312.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@68313.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@68314.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@68315.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@68316.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@68317.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@68318.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@68319.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@68240.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@68241.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@68242.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@68243.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@68244.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@68245.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@68246.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@68247.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@68248.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@68249.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@68250.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@68251.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@68252.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@68253.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@68254.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@68255.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@68256.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@68257.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@68258.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@68259.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@68260.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@68261.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@68262.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@68263.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@68264.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@68265.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@68266.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@68267.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@68268.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@68269.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@68270.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@68271.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@68272.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@68273.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@68274.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@68275.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@68276.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@68277.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@68278.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@68279.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@68280.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@68281.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@68282.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@68283.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@68284.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@68285.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@68286.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@68287.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@68288.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@68289.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@68290.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@68291.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@68292.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@68293.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@68294.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@68295.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@68296.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@68297.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@68298.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@68299.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@68300.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@68301.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@68302.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@68303.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@68238.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@68219.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@68443.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@68436.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@68333.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@68332.4]
  assign AXICmdSplit_clock = clock; // @[:@68330.4]
  assign AXICmdSplit_reset = reset; // @[:@68331.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@68442.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@68441.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@68440.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@68438.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@68437.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@68435.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@68419.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@68420.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@68421.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@68422.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@68423.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@68424.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@68425.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@68426.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@68427.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@68428.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@68429.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@68430.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@68431.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@68432.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@68433.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@68434.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@68355.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@68356.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@68357.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@68358.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@68359.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@68360.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@68361.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@68362.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@68363.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@68364.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@68365.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@68366.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@68367.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@68368.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@68369.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@68370.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@68371.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@68372.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@68373.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@68374.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@68375.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@68376.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@68377.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@68378.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@68379.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@68380.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@68381.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@68382.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@68383.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@68384.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@68385.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@68386.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@68387.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@68388.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@68389.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@68390.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@68391.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@68392.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@68393.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@68394.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@68395.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@68396.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@68397.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@68398.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@68399.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@68400.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@68401.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@68402.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@68403.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@68404.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@68405.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@68406.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@68407.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@68408.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@68409.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@68410.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@68411.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@68412.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@68413.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@68414.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@68415.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@68416.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@68417.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@68418.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@68353.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@68334.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@68558.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@68551.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@68448.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@68447.4]
  assign AXICmdIssue_clock = clock; // @[:@68445.4]
  assign AXICmdIssue_reset = reset; // @[:@68446.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@68557.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@68556.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@68555.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@68553.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@68552.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@68550.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@68534.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@68535.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@68536.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@68537.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@68538.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@68539.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@68540.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@68541.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@68542.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@68543.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@68544.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@68545.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@68546.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@68547.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@68548.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@68549.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@68470.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@68471.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@68472.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@68473.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@68474.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@68475.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@68476.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@68477.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@68478.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@68479.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@68480.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@68481.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@68482.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@68483.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@68484.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@68485.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@68486.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@68487.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@68488.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@68489.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@68490.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@68491.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@68492.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@68493.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@68494.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@68495.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@68496.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@68497.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@68498.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@68499.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@68500.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@68501.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@68502.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@68503.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@68504.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@68505.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@68506.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@68507.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@68508.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@68509.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@68510.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@68511.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@68512.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@68513.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@68514.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@68515.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@68516.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@68517.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@68518.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@68519.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@68520.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@68521.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@68522.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@68523.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@68524.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@68525.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@68526.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@68527.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@68528.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@68529.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@68530.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@68531.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@68532.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@68533.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@68468.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@68449.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@68670.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@68663.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@68560.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@68559.4]
endmodule
module DRAMArbiter_1( // @[:@82899.2]
  input         clock, // @[:@82900.4]
  input         reset, // @[:@82901.4]
  input         io_enable, // @[:@82902.4]
  input         io_dram_cmd_ready, // @[:@82902.4]
  output        io_dram_cmd_valid, // @[:@82902.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@82902.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@82902.4]
  output        io_dram_cmd_bits_isWr, // @[:@82902.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@82902.4]
  input         io_dram_wdata_ready, // @[:@82902.4]
  output        io_dram_wdata_valid, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@82902.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@82902.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@82902.4]
  output        io_dram_wdata_bits_wlast, // @[:@82902.4]
  output        io_dram_rresp_ready, // @[:@82902.4]
  output        io_dram_wresp_ready, // @[:@82902.4]
  input         io_dram_wresp_valid, // @[:@82902.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@82902.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@83788.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@83802.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@84030.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@84145.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@84145.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@83788.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@83802.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@84030.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@84145.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@84370.4 DRAMArbiter.scala 100:23:@84373.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@84369.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@84368.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@84366.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@84365.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@84363.4 DRAMArbiter.scala 101:25:@84375.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@84347.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@84348.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@84349.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@84350.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@84351.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@84352.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@84353.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@84354.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@84355.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@84356.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@84357.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@84358.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@84359.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@84360.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@84361.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@84362.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@84283.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@84284.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@84285.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@84286.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@84287.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@84288.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@84289.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@84290.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@84291.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@84292.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@84293.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@84294.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@84295.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@84296.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@84297.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@84298.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@84299.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@84300.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@84301.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@84302.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@84303.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@84304.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@84305.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@84306.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@84307.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@84308.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@84309.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@84310.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@84311.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@84312.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@84313.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@84314.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@84315.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@84316.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@84317.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@84318.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@84319.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@84320.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@84321.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@84322.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@84323.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@84324.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@84325.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@84326.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@84327.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@84328.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@84329.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@84330.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@84331.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@84332.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@84333.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@84334.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@84335.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@84336.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@84337.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@84338.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@84339.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@84340.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@84341.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@84342.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@84343.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@84344.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@84345.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@84346.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@84282.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@84281.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@84262.4]
  assign StreamControllerStore_clock = clock; // @[:@83789.4]
  assign StreamControllerStore_reset = reset; // @[:@83790.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@83917.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@83910.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@83807.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@83800.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@83799.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@83798.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@83796.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@83795.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@83794.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@83793.4]
  assign StreamArbiter_clock = clock; // @[:@83803.4]
  assign StreamArbiter_reset = reset; // @[:@83804.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@84028.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@84027.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@84026.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@84024.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@84023.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@84021.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@84005.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@84006.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@84007.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@84008.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@84009.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@84010.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@84011.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@84012.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@84013.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@84014.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@84015.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@84016.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@84017.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@84018.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@84019.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@84020.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@83941.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@83942.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@83943.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@83944.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@83945.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@83946.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@83947.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@83948.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@83949.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@83950.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@83951.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@83952.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@83953.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@83954.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@83955.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@83956.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@83957.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@83958.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@83959.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@83960.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@83961.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@83962.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@83963.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@83964.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@83965.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@83966.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@83967.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@83968.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@83969.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@83970.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@83971.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@83972.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@83973.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@83974.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@83975.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@83976.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@83977.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@83978.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@83979.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@83980.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@83981.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@83982.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@83983.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@83984.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@83985.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@83986.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@83987.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@83988.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@83989.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@83990.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@83991.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@83992.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@83993.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@83994.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@83995.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@83996.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@83997.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@83998.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@83999.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@84000.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@84001.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@84002.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@84003.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@84004.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@83939.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@83920.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@84144.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@84137.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@84034.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@84033.4]
  assign AXICmdSplit_clock = clock; // @[:@84031.4]
  assign AXICmdSplit_reset = reset; // @[:@84032.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@84143.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@84142.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@84141.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@84139.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@84138.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@84136.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@84120.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@84121.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@84122.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@84123.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@84124.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@84125.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@84126.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@84127.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@84128.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@84129.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@84130.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@84131.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@84132.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@84133.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@84134.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@84135.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@84056.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@84057.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@84058.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@84059.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@84060.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@84061.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@84062.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@84063.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@84064.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@84065.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@84066.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@84067.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@84068.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@84069.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@84070.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@84071.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@84072.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@84073.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@84074.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@84075.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@84076.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@84077.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@84078.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@84079.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@84080.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@84081.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@84082.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@84083.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@84084.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@84085.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@84086.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@84087.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@84088.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@84089.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@84090.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@84091.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@84092.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@84093.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@84094.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@84095.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@84096.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@84097.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@84098.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@84099.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@84100.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@84101.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@84102.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@84103.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@84104.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@84105.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@84106.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@84107.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@84108.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@84109.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@84110.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@84111.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@84112.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@84113.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@84114.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@84115.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@84116.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@84117.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@84118.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@84119.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@84054.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@84035.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@84259.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@84252.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@84149.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@84148.4]
  assign AXICmdIssue_clock = clock; // @[:@84146.4]
  assign AXICmdIssue_reset = reset; // @[:@84147.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@84258.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@84257.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@84256.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@84254.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@84253.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@84251.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@84235.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@84236.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@84237.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@84238.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@84239.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@84240.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@84241.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@84242.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@84243.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@84244.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@84245.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@84246.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@84247.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@84248.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@84249.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@84250.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@84171.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@84172.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@84173.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@84174.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@84175.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@84176.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@84177.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@84178.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@84179.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@84180.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@84181.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@84182.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@84183.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@84184.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@84185.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@84186.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@84187.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@84188.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@84189.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@84190.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@84191.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@84192.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@84193.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@84194.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@84195.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@84196.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@84197.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@84198.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@84199.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@84200.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@84201.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@84202.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@84203.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@84204.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@84205.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@84206.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@84207.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@84208.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@84209.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@84210.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@84211.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@84212.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@84213.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@84214.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@84215.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@84216.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@84217.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@84218.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@84219.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@84220.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@84221.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@84222.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@84223.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@84224.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@84225.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@84226.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@84227.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@84228.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@84229.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@84230.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@84231.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@84232.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@84233.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@84234.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@84169.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@84150.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@84371.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@84364.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@84261.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@84260.4]
endmodule
module DRAMHeap( // @[:@115007.2]
  input         io_accel_0_req_valid, // @[:@115010.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@115010.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@115010.4]
  output        io_accel_0_resp_valid, // @[:@115010.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@115010.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@115010.4]
  output        io_host_0_req_valid, // @[:@115010.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@115010.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@115010.4]
  input         io_host_0_resp_valid, // @[:@115010.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@115010.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@115010.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@115017.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@115019.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@115018.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@115014.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@115013.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@115012.4]
endmodule
module RetimeWrapper_541( // @[:@115033.2]
  input         clock, // @[:@115034.4]
  input         reset, // @[:@115035.4]
  input         io_flow, // @[:@115036.4]
  input  [63:0] io_in, // @[:@115036.4]
  output [63:0] io_out // @[:@115036.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@115038.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@115038.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@115038.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@115038.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@115038.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@115038.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@115038.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@115051.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@115050.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@115049.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@115048.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@115047.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@115045.4]
endmodule
module FringeFF( // @[:@115053.2]
  input         clock, // @[:@115054.4]
  input         reset, // @[:@115055.4]
  input  [63:0] io_in, // @[:@115056.4]
  input         io_reset, // @[:@115056.4]
  output [63:0] io_out, // @[:@115056.4]
  input         io_enable // @[:@115056.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@115059.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@115059.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@115059.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@115059.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@115059.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@115064.4 package.scala 96:25:@115065.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@115070.6]
  RetimeWrapper_541 RetimeWrapper ( // @[package.scala 93:22:@115059.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@115064.4 package.scala 96:25:@115065.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@115070.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@115076.4]
  assign RetimeWrapper_clock = clock; // @[:@115060.4]
  assign RetimeWrapper_reset = reset; // @[:@115061.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@115063.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@115062.4]
endmodule
module MuxN( // @[:@143692.2]
  input  [63:0] io_ins_0, // @[:@143695.4]
  input  [63:0] io_ins_1, // @[:@143695.4]
  input  [63:0] io_ins_2, // @[:@143695.4]
  input  [63:0] io_ins_3, // @[:@143695.4]
  input  [63:0] io_ins_4, // @[:@143695.4]
  input  [63:0] io_ins_5, // @[:@143695.4]
  input  [63:0] io_ins_6, // @[:@143695.4]
  input  [63:0] io_ins_7, // @[:@143695.4]
  input  [63:0] io_ins_8, // @[:@143695.4]
  input  [63:0] io_ins_9, // @[:@143695.4]
  input  [63:0] io_ins_10, // @[:@143695.4]
  input  [63:0] io_ins_11, // @[:@143695.4]
  input  [63:0] io_ins_12, // @[:@143695.4]
  input  [63:0] io_ins_13, // @[:@143695.4]
  input  [63:0] io_ins_14, // @[:@143695.4]
  input  [63:0] io_ins_15, // @[:@143695.4]
  input  [63:0] io_ins_16, // @[:@143695.4]
  input  [63:0] io_ins_17, // @[:@143695.4]
  input  [63:0] io_ins_18, // @[:@143695.4]
  input  [63:0] io_ins_19, // @[:@143695.4]
  input  [63:0] io_ins_20, // @[:@143695.4]
  input  [63:0] io_ins_21, // @[:@143695.4]
  input  [63:0] io_ins_22, // @[:@143695.4]
  input  [63:0] io_ins_23, // @[:@143695.4]
  input  [63:0] io_ins_24, // @[:@143695.4]
  input  [63:0] io_ins_25, // @[:@143695.4]
  input  [63:0] io_ins_26, // @[:@143695.4]
  input  [63:0] io_ins_27, // @[:@143695.4]
  input  [63:0] io_ins_28, // @[:@143695.4]
  input  [63:0] io_ins_29, // @[:@143695.4]
  input  [63:0] io_ins_30, // @[:@143695.4]
  input  [63:0] io_ins_31, // @[:@143695.4]
  input  [63:0] io_ins_32, // @[:@143695.4]
  input  [63:0] io_ins_33, // @[:@143695.4]
  input  [63:0] io_ins_34, // @[:@143695.4]
  input  [63:0] io_ins_35, // @[:@143695.4]
  input  [63:0] io_ins_36, // @[:@143695.4]
  input  [63:0] io_ins_37, // @[:@143695.4]
  input  [63:0] io_ins_38, // @[:@143695.4]
  input  [63:0] io_ins_39, // @[:@143695.4]
  input  [63:0] io_ins_40, // @[:@143695.4]
  input  [63:0] io_ins_41, // @[:@143695.4]
  input  [63:0] io_ins_42, // @[:@143695.4]
  input  [63:0] io_ins_43, // @[:@143695.4]
  input  [63:0] io_ins_44, // @[:@143695.4]
  input  [63:0] io_ins_45, // @[:@143695.4]
  input  [63:0] io_ins_46, // @[:@143695.4]
  input  [63:0] io_ins_47, // @[:@143695.4]
  input  [63:0] io_ins_48, // @[:@143695.4]
  input  [63:0] io_ins_49, // @[:@143695.4]
  input  [63:0] io_ins_50, // @[:@143695.4]
  input  [63:0] io_ins_51, // @[:@143695.4]
  input  [63:0] io_ins_52, // @[:@143695.4]
  input  [63:0] io_ins_53, // @[:@143695.4]
  input  [63:0] io_ins_54, // @[:@143695.4]
  input  [63:0] io_ins_55, // @[:@143695.4]
  input  [63:0] io_ins_56, // @[:@143695.4]
  input  [63:0] io_ins_57, // @[:@143695.4]
  input  [63:0] io_ins_58, // @[:@143695.4]
  input  [63:0] io_ins_59, // @[:@143695.4]
  input  [63:0] io_ins_60, // @[:@143695.4]
  input  [63:0] io_ins_61, // @[:@143695.4]
  input  [63:0] io_ins_62, // @[:@143695.4]
  input  [63:0] io_ins_63, // @[:@143695.4]
  input  [63:0] io_ins_64, // @[:@143695.4]
  input  [63:0] io_ins_65, // @[:@143695.4]
  input  [63:0] io_ins_66, // @[:@143695.4]
  input  [63:0] io_ins_67, // @[:@143695.4]
  input  [63:0] io_ins_68, // @[:@143695.4]
  input  [63:0] io_ins_69, // @[:@143695.4]
  input  [63:0] io_ins_70, // @[:@143695.4]
  input  [63:0] io_ins_71, // @[:@143695.4]
  input  [63:0] io_ins_72, // @[:@143695.4]
  input  [63:0] io_ins_73, // @[:@143695.4]
  input  [63:0] io_ins_74, // @[:@143695.4]
  input  [63:0] io_ins_75, // @[:@143695.4]
  input  [63:0] io_ins_76, // @[:@143695.4]
  input  [63:0] io_ins_77, // @[:@143695.4]
  input  [63:0] io_ins_78, // @[:@143695.4]
  input  [63:0] io_ins_79, // @[:@143695.4]
  input  [63:0] io_ins_80, // @[:@143695.4]
  input  [63:0] io_ins_81, // @[:@143695.4]
  input  [63:0] io_ins_82, // @[:@143695.4]
  input  [63:0] io_ins_83, // @[:@143695.4]
  input  [63:0] io_ins_84, // @[:@143695.4]
  input  [63:0] io_ins_85, // @[:@143695.4]
  input  [63:0] io_ins_86, // @[:@143695.4]
  input  [63:0] io_ins_87, // @[:@143695.4]
  input  [63:0] io_ins_88, // @[:@143695.4]
  input  [63:0] io_ins_89, // @[:@143695.4]
  input  [63:0] io_ins_90, // @[:@143695.4]
  input  [63:0] io_ins_91, // @[:@143695.4]
  input  [63:0] io_ins_92, // @[:@143695.4]
  input  [63:0] io_ins_93, // @[:@143695.4]
  input  [63:0] io_ins_94, // @[:@143695.4]
  input  [63:0] io_ins_95, // @[:@143695.4]
  input  [63:0] io_ins_96, // @[:@143695.4]
  input  [63:0] io_ins_97, // @[:@143695.4]
  input  [63:0] io_ins_98, // @[:@143695.4]
  input  [63:0] io_ins_99, // @[:@143695.4]
  input  [63:0] io_ins_100, // @[:@143695.4]
  input  [63:0] io_ins_101, // @[:@143695.4]
  input  [63:0] io_ins_102, // @[:@143695.4]
  input  [63:0] io_ins_103, // @[:@143695.4]
  input  [63:0] io_ins_104, // @[:@143695.4]
  input  [63:0] io_ins_105, // @[:@143695.4]
  input  [63:0] io_ins_106, // @[:@143695.4]
  input  [63:0] io_ins_107, // @[:@143695.4]
  input  [63:0] io_ins_108, // @[:@143695.4]
  input  [63:0] io_ins_109, // @[:@143695.4]
  input  [63:0] io_ins_110, // @[:@143695.4]
  input  [63:0] io_ins_111, // @[:@143695.4]
  input  [63:0] io_ins_112, // @[:@143695.4]
  input  [63:0] io_ins_113, // @[:@143695.4]
  input  [63:0] io_ins_114, // @[:@143695.4]
  input  [63:0] io_ins_115, // @[:@143695.4]
  input  [63:0] io_ins_116, // @[:@143695.4]
  input  [63:0] io_ins_117, // @[:@143695.4]
  input  [63:0] io_ins_118, // @[:@143695.4]
  input  [63:0] io_ins_119, // @[:@143695.4]
  input  [63:0] io_ins_120, // @[:@143695.4]
  input  [63:0] io_ins_121, // @[:@143695.4]
  input  [63:0] io_ins_122, // @[:@143695.4]
  input  [63:0] io_ins_123, // @[:@143695.4]
  input  [63:0] io_ins_124, // @[:@143695.4]
  input  [63:0] io_ins_125, // @[:@143695.4]
  input  [63:0] io_ins_126, // @[:@143695.4]
  input  [63:0] io_ins_127, // @[:@143695.4]
  input  [63:0] io_ins_128, // @[:@143695.4]
  input  [63:0] io_ins_129, // @[:@143695.4]
  input  [63:0] io_ins_130, // @[:@143695.4]
  input  [63:0] io_ins_131, // @[:@143695.4]
  input  [63:0] io_ins_132, // @[:@143695.4]
  input  [63:0] io_ins_133, // @[:@143695.4]
  input  [63:0] io_ins_134, // @[:@143695.4]
  input  [63:0] io_ins_135, // @[:@143695.4]
  input  [63:0] io_ins_136, // @[:@143695.4]
  input  [63:0] io_ins_137, // @[:@143695.4]
  input  [63:0] io_ins_138, // @[:@143695.4]
  input  [63:0] io_ins_139, // @[:@143695.4]
  input  [63:0] io_ins_140, // @[:@143695.4]
  input  [63:0] io_ins_141, // @[:@143695.4]
  input  [63:0] io_ins_142, // @[:@143695.4]
  input  [63:0] io_ins_143, // @[:@143695.4]
  input  [63:0] io_ins_144, // @[:@143695.4]
  input  [63:0] io_ins_145, // @[:@143695.4]
  input  [63:0] io_ins_146, // @[:@143695.4]
  input  [63:0] io_ins_147, // @[:@143695.4]
  input  [63:0] io_ins_148, // @[:@143695.4]
  input  [63:0] io_ins_149, // @[:@143695.4]
  input  [63:0] io_ins_150, // @[:@143695.4]
  input  [63:0] io_ins_151, // @[:@143695.4]
  input  [63:0] io_ins_152, // @[:@143695.4]
  input  [63:0] io_ins_153, // @[:@143695.4]
  input  [63:0] io_ins_154, // @[:@143695.4]
  input  [63:0] io_ins_155, // @[:@143695.4]
  input  [63:0] io_ins_156, // @[:@143695.4]
  input  [63:0] io_ins_157, // @[:@143695.4]
  input  [63:0] io_ins_158, // @[:@143695.4]
  input  [63:0] io_ins_159, // @[:@143695.4]
  input  [63:0] io_ins_160, // @[:@143695.4]
  input  [63:0] io_ins_161, // @[:@143695.4]
  input  [63:0] io_ins_162, // @[:@143695.4]
  input  [63:0] io_ins_163, // @[:@143695.4]
  input  [63:0] io_ins_164, // @[:@143695.4]
  input  [63:0] io_ins_165, // @[:@143695.4]
  input  [63:0] io_ins_166, // @[:@143695.4]
  input  [63:0] io_ins_167, // @[:@143695.4]
  input  [63:0] io_ins_168, // @[:@143695.4]
  input  [63:0] io_ins_169, // @[:@143695.4]
  input  [63:0] io_ins_170, // @[:@143695.4]
  input  [63:0] io_ins_171, // @[:@143695.4]
  input  [63:0] io_ins_172, // @[:@143695.4]
  input  [63:0] io_ins_173, // @[:@143695.4]
  input  [63:0] io_ins_174, // @[:@143695.4]
  input  [63:0] io_ins_175, // @[:@143695.4]
  input  [63:0] io_ins_176, // @[:@143695.4]
  input  [63:0] io_ins_177, // @[:@143695.4]
  input  [63:0] io_ins_178, // @[:@143695.4]
  input  [63:0] io_ins_179, // @[:@143695.4]
  input  [63:0] io_ins_180, // @[:@143695.4]
  input  [63:0] io_ins_181, // @[:@143695.4]
  input  [63:0] io_ins_182, // @[:@143695.4]
  input  [63:0] io_ins_183, // @[:@143695.4]
  input  [63:0] io_ins_184, // @[:@143695.4]
  input  [63:0] io_ins_185, // @[:@143695.4]
  input  [63:0] io_ins_186, // @[:@143695.4]
  input  [63:0] io_ins_187, // @[:@143695.4]
  input  [63:0] io_ins_188, // @[:@143695.4]
  input  [63:0] io_ins_189, // @[:@143695.4]
  input  [63:0] io_ins_190, // @[:@143695.4]
  input  [63:0] io_ins_191, // @[:@143695.4]
  input  [63:0] io_ins_192, // @[:@143695.4]
  input  [63:0] io_ins_193, // @[:@143695.4]
  input  [63:0] io_ins_194, // @[:@143695.4]
  input  [63:0] io_ins_195, // @[:@143695.4]
  input  [63:0] io_ins_196, // @[:@143695.4]
  input  [63:0] io_ins_197, // @[:@143695.4]
  input  [63:0] io_ins_198, // @[:@143695.4]
  input  [63:0] io_ins_199, // @[:@143695.4]
  input  [63:0] io_ins_200, // @[:@143695.4]
  input  [63:0] io_ins_201, // @[:@143695.4]
  input  [63:0] io_ins_202, // @[:@143695.4]
  input  [63:0] io_ins_203, // @[:@143695.4]
  input  [63:0] io_ins_204, // @[:@143695.4]
  input  [63:0] io_ins_205, // @[:@143695.4]
  input  [63:0] io_ins_206, // @[:@143695.4]
  input  [63:0] io_ins_207, // @[:@143695.4]
  input  [63:0] io_ins_208, // @[:@143695.4]
  input  [63:0] io_ins_209, // @[:@143695.4]
  input  [63:0] io_ins_210, // @[:@143695.4]
  input  [63:0] io_ins_211, // @[:@143695.4]
  input  [63:0] io_ins_212, // @[:@143695.4]
  input  [63:0] io_ins_213, // @[:@143695.4]
  input  [63:0] io_ins_214, // @[:@143695.4]
  input  [63:0] io_ins_215, // @[:@143695.4]
  input  [63:0] io_ins_216, // @[:@143695.4]
  input  [63:0] io_ins_217, // @[:@143695.4]
  input  [63:0] io_ins_218, // @[:@143695.4]
  input  [63:0] io_ins_219, // @[:@143695.4]
  input  [63:0] io_ins_220, // @[:@143695.4]
  input  [63:0] io_ins_221, // @[:@143695.4]
  input  [63:0] io_ins_222, // @[:@143695.4]
  input  [63:0] io_ins_223, // @[:@143695.4]
  input  [63:0] io_ins_224, // @[:@143695.4]
  input  [63:0] io_ins_225, // @[:@143695.4]
  input  [63:0] io_ins_226, // @[:@143695.4]
  input  [63:0] io_ins_227, // @[:@143695.4]
  input  [63:0] io_ins_228, // @[:@143695.4]
  input  [63:0] io_ins_229, // @[:@143695.4]
  input  [63:0] io_ins_230, // @[:@143695.4]
  input  [63:0] io_ins_231, // @[:@143695.4]
  input  [63:0] io_ins_232, // @[:@143695.4]
  input  [63:0] io_ins_233, // @[:@143695.4]
  input  [63:0] io_ins_234, // @[:@143695.4]
  input  [63:0] io_ins_235, // @[:@143695.4]
  input  [63:0] io_ins_236, // @[:@143695.4]
  input  [63:0] io_ins_237, // @[:@143695.4]
  input  [63:0] io_ins_238, // @[:@143695.4]
  input  [63:0] io_ins_239, // @[:@143695.4]
  input  [63:0] io_ins_240, // @[:@143695.4]
  input  [63:0] io_ins_241, // @[:@143695.4]
  input  [63:0] io_ins_242, // @[:@143695.4]
  input  [63:0] io_ins_243, // @[:@143695.4]
  input  [63:0] io_ins_244, // @[:@143695.4]
  input  [63:0] io_ins_245, // @[:@143695.4]
  input  [63:0] io_ins_246, // @[:@143695.4]
  input  [63:0] io_ins_247, // @[:@143695.4]
  input  [63:0] io_ins_248, // @[:@143695.4]
  input  [63:0] io_ins_249, // @[:@143695.4]
  input  [63:0] io_ins_250, // @[:@143695.4]
  input  [63:0] io_ins_251, // @[:@143695.4]
  input  [63:0] io_ins_252, // @[:@143695.4]
  input  [63:0] io_ins_253, // @[:@143695.4]
  input  [63:0] io_ins_254, // @[:@143695.4]
  input  [63:0] io_ins_255, // @[:@143695.4]
  input  [63:0] io_ins_256, // @[:@143695.4]
  input  [63:0] io_ins_257, // @[:@143695.4]
  input  [63:0] io_ins_258, // @[:@143695.4]
  input  [63:0] io_ins_259, // @[:@143695.4]
  input  [63:0] io_ins_260, // @[:@143695.4]
  input  [63:0] io_ins_261, // @[:@143695.4]
  input  [63:0] io_ins_262, // @[:@143695.4]
  input  [63:0] io_ins_263, // @[:@143695.4]
  input  [63:0] io_ins_264, // @[:@143695.4]
  input  [63:0] io_ins_265, // @[:@143695.4]
  input  [63:0] io_ins_266, // @[:@143695.4]
  input  [63:0] io_ins_267, // @[:@143695.4]
  input  [63:0] io_ins_268, // @[:@143695.4]
  input  [63:0] io_ins_269, // @[:@143695.4]
  input  [63:0] io_ins_270, // @[:@143695.4]
  input  [63:0] io_ins_271, // @[:@143695.4]
  input  [63:0] io_ins_272, // @[:@143695.4]
  input  [63:0] io_ins_273, // @[:@143695.4]
  input  [63:0] io_ins_274, // @[:@143695.4]
  input  [63:0] io_ins_275, // @[:@143695.4]
  input  [63:0] io_ins_276, // @[:@143695.4]
  input  [63:0] io_ins_277, // @[:@143695.4]
  input  [63:0] io_ins_278, // @[:@143695.4]
  input  [63:0] io_ins_279, // @[:@143695.4]
  input  [63:0] io_ins_280, // @[:@143695.4]
  input  [63:0] io_ins_281, // @[:@143695.4]
  input  [63:0] io_ins_282, // @[:@143695.4]
  input  [63:0] io_ins_283, // @[:@143695.4]
  input  [63:0] io_ins_284, // @[:@143695.4]
  input  [63:0] io_ins_285, // @[:@143695.4]
  input  [63:0] io_ins_286, // @[:@143695.4]
  input  [63:0] io_ins_287, // @[:@143695.4]
  input  [63:0] io_ins_288, // @[:@143695.4]
  input  [63:0] io_ins_289, // @[:@143695.4]
  input  [63:0] io_ins_290, // @[:@143695.4]
  input  [63:0] io_ins_291, // @[:@143695.4]
  input  [63:0] io_ins_292, // @[:@143695.4]
  input  [63:0] io_ins_293, // @[:@143695.4]
  input  [63:0] io_ins_294, // @[:@143695.4]
  input  [63:0] io_ins_295, // @[:@143695.4]
  input  [63:0] io_ins_296, // @[:@143695.4]
  input  [63:0] io_ins_297, // @[:@143695.4]
  input  [63:0] io_ins_298, // @[:@143695.4]
  input  [63:0] io_ins_299, // @[:@143695.4]
  input  [63:0] io_ins_300, // @[:@143695.4]
  input  [63:0] io_ins_301, // @[:@143695.4]
  input  [63:0] io_ins_302, // @[:@143695.4]
  input  [63:0] io_ins_303, // @[:@143695.4]
  input  [63:0] io_ins_304, // @[:@143695.4]
  input  [63:0] io_ins_305, // @[:@143695.4]
  input  [63:0] io_ins_306, // @[:@143695.4]
  input  [63:0] io_ins_307, // @[:@143695.4]
  input  [63:0] io_ins_308, // @[:@143695.4]
  input  [63:0] io_ins_309, // @[:@143695.4]
  input  [63:0] io_ins_310, // @[:@143695.4]
  input  [63:0] io_ins_311, // @[:@143695.4]
  input  [63:0] io_ins_312, // @[:@143695.4]
  input  [63:0] io_ins_313, // @[:@143695.4]
  input  [63:0] io_ins_314, // @[:@143695.4]
  input  [63:0] io_ins_315, // @[:@143695.4]
  input  [63:0] io_ins_316, // @[:@143695.4]
  input  [63:0] io_ins_317, // @[:@143695.4]
  input  [63:0] io_ins_318, // @[:@143695.4]
  input  [63:0] io_ins_319, // @[:@143695.4]
  input  [63:0] io_ins_320, // @[:@143695.4]
  input  [63:0] io_ins_321, // @[:@143695.4]
  input  [63:0] io_ins_322, // @[:@143695.4]
  input  [63:0] io_ins_323, // @[:@143695.4]
  input  [63:0] io_ins_324, // @[:@143695.4]
  input  [63:0] io_ins_325, // @[:@143695.4]
  input  [63:0] io_ins_326, // @[:@143695.4]
  input  [63:0] io_ins_327, // @[:@143695.4]
  input  [63:0] io_ins_328, // @[:@143695.4]
  input  [63:0] io_ins_329, // @[:@143695.4]
  input  [63:0] io_ins_330, // @[:@143695.4]
  input  [63:0] io_ins_331, // @[:@143695.4]
  input  [63:0] io_ins_332, // @[:@143695.4]
  input  [63:0] io_ins_333, // @[:@143695.4]
  input  [63:0] io_ins_334, // @[:@143695.4]
  input  [63:0] io_ins_335, // @[:@143695.4]
  input  [63:0] io_ins_336, // @[:@143695.4]
  input  [63:0] io_ins_337, // @[:@143695.4]
  input  [63:0] io_ins_338, // @[:@143695.4]
  input  [63:0] io_ins_339, // @[:@143695.4]
  input  [63:0] io_ins_340, // @[:@143695.4]
  input  [63:0] io_ins_341, // @[:@143695.4]
  input  [63:0] io_ins_342, // @[:@143695.4]
  input  [63:0] io_ins_343, // @[:@143695.4]
  input  [63:0] io_ins_344, // @[:@143695.4]
  input  [63:0] io_ins_345, // @[:@143695.4]
  input  [63:0] io_ins_346, // @[:@143695.4]
  input  [63:0] io_ins_347, // @[:@143695.4]
  input  [63:0] io_ins_348, // @[:@143695.4]
  input  [63:0] io_ins_349, // @[:@143695.4]
  input  [63:0] io_ins_350, // @[:@143695.4]
  input  [63:0] io_ins_351, // @[:@143695.4]
  input  [63:0] io_ins_352, // @[:@143695.4]
  input  [63:0] io_ins_353, // @[:@143695.4]
  input  [63:0] io_ins_354, // @[:@143695.4]
  input  [63:0] io_ins_355, // @[:@143695.4]
  input  [63:0] io_ins_356, // @[:@143695.4]
  input  [63:0] io_ins_357, // @[:@143695.4]
  input  [63:0] io_ins_358, // @[:@143695.4]
  input  [63:0] io_ins_359, // @[:@143695.4]
  input  [63:0] io_ins_360, // @[:@143695.4]
  input  [63:0] io_ins_361, // @[:@143695.4]
  input  [63:0] io_ins_362, // @[:@143695.4]
  input  [63:0] io_ins_363, // @[:@143695.4]
  input  [63:0] io_ins_364, // @[:@143695.4]
  input  [63:0] io_ins_365, // @[:@143695.4]
  input  [63:0] io_ins_366, // @[:@143695.4]
  input  [63:0] io_ins_367, // @[:@143695.4]
  input  [63:0] io_ins_368, // @[:@143695.4]
  input  [63:0] io_ins_369, // @[:@143695.4]
  input  [63:0] io_ins_370, // @[:@143695.4]
  input  [63:0] io_ins_371, // @[:@143695.4]
  input  [63:0] io_ins_372, // @[:@143695.4]
  input  [63:0] io_ins_373, // @[:@143695.4]
  input  [63:0] io_ins_374, // @[:@143695.4]
  input  [63:0] io_ins_375, // @[:@143695.4]
  input  [63:0] io_ins_376, // @[:@143695.4]
  input  [63:0] io_ins_377, // @[:@143695.4]
  input  [63:0] io_ins_378, // @[:@143695.4]
  input  [63:0] io_ins_379, // @[:@143695.4]
  input  [63:0] io_ins_380, // @[:@143695.4]
  input  [63:0] io_ins_381, // @[:@143695.4]
  input  [63:0] io_ins_382, // @[:@143695.4]
  input  [63:0] io_ins_383, // @[:@143695.4]
  input  [63:0] io_ins_384, // @[:@143695.4]
  input  [63:0] io_ins_385, // @[:@143695.4]
  input  [63:0] io_ins_386, // @[:@143695.4]
  input  [63:0] io_ins_387, // @[:@143695.4]
  input  [63:0] io_ins_388, // @[:@143695.4]
  input  [63:0] io_ins_389, // @[:@143695.4]
  input  [63:0] io_ins_390, // @[:@143695.4]
  input  [63:0] io_ins_391, // @[:@143695.4]
  input  [63:0] io_ins_392, // @[:@143695.4]
  input  [63:0] io_ins_393, // @[:@143695.4]
  input  [63:0] io_ins_394, // @[:@143695.4]
  input  [63:0] io_ins_395, // @[:@143695.4]
  input  [63:0] io_ins_396, // @[:@143695.4]
  input  [63:0] io_ins_397, // @[:@143695.4]
  input  [63:0] io_ins_398, // @[:@143695.4]
  input  [63:0] io_ins_399, // @[:@143695.4]
  input  [63:0] io_ins_400, // @[:@143695.4]
  input  [63:0] io_ins_401, // @[:@143695.4]
  input  [63:0] io_ins_402, // @[:@143695.4]
  input  [63:0] io_ins_403, // @[:@143695.4]
  input  [63:0] io_ins_404, // @[:@143695.4]
  input  [63:0] io_ins_405, // @[:@143695.4]
  input  [63:0] io_ins_406, // @[:@143695.4]
  input  [63:0] io_ins_407, // @[:@143695.4]
  input  [63:0] io_ins_408, // @[:@143695.4]
  input  [63:0] io_ins_409, // @[:@143695.4]
  input  [63:0] io_ins_410, // @[:@143695.4]
  input  [63:0] io_ins_411, // @[:@143695.4]
  input  [63:0] io_ins_412, // @[:@143695.4]
  input  [63:0] io_ins_413, // @[:@143695.4]
  input  [63:0] io_ins_414, // @[:@143695.4]
  input  [63:0] io_ins_415, // @[:@143695.4]
  input  [63:0] io_ins_416, // @[:@143695.4]
  input  [63:0] io_ins_417, // @[:@143695.4]
  input  [63:0] io_ins_418, // @[:@143695.4]
  input  [63:0] io_ins_419, // @[:@143695.4]
  input  [63:0] io_ins_420, // @[:@143695.4]
  input  [63:0] io_ins_421, // @[:@143695.4]
  input  [63:0] io_ins_422, // @[:@143695.4]
  input  [63:0] io_ins_423, // @[:@143695.4]
  input  [63:0] io_ins_424, // @[:@143695.4]
  input  [63:0] io_ins_425, // @[:@143695.4]
  input  [63:0] io_ins_426, // @[:@143695.4]
  input  [63:0] io_ins_427, // @[:@143695.4]
  input  [63:0] io_ins_428, // @[:@143695.4]
  input  [63:0] io_ins_429, // @[:@143695.4]
  input  [63:0] io_ins_430, // @[:@143695.4]
  input  [63:0] io_ins_431, // @[:@143695.4]
  input  [63:0] io_ins_432, // @[:@143695.4]
  input  [63:0] io_ins_433, // @[:@143695.4]
  input  [63:0] io_ins_434, // @[:@143695.4]
  input  [63:0] io_ins_435, // @[:@143695.4]
  input  [63:0] io_ins_436, // @[:@143695.4]
  input  [63:0] io_ins_437, // @[:@143695.4]
  input  [63:0] io_ins_438, // @[:@143695.4]
  input  [63:0] io_ins_439, // @[:@143695.4]
  input  [63:0] io_ins_440, // @[:@143695.4]
  input  [63:0] io_ins_441, // @[:@143695.4]
  input  [63:0] io_ins_442, // @[:@143695.4]
  input  [63:0] io_ins_443, // @[:@143695.4]
  input  [63:0] io_ins_444, // @[:@143695.4]
  input  [63:0] io_ins_445, // @[:@143695.4]
  input  [63:0] io_ins_446, // @[:@143695.4]
  input  [63:0] io_ins_447, // @[:@143695.4]
  input  [63:0] io_ins_448, // @[:@143695.4]
  input  [63:0] io_ins_449, // @[:@143695.4]
  input  [63:0] io_ins_450, // @[:@143695.4]
  input  [63:0] io_ins_451, // @[:@143695.4]
  input  [63:0] io_ins_452, // @[:@143695.4]
  input  [63:0] io_ins_453, // @[:@143695.4]
  input  [63:0] io_ins_454, // @[:@143695.4]
  input  [63:0] io_ins_455, // @[:@143695.4]
  input  [63:0] io_ins_456, // @[:@143695.4]
  input  [63:0] io_ins_457, // @[:@143695.4]
  input  [63:0] io_ins_458, // @[:@143695.4]
  input  [63:0] io_ins_459, // @[:@143695.4]
  input  [63:0] io_ins_460, // @[:@143695.4]
  input  [63:0] io_ins_461, // @[:@143695.4]
  input  [63:0] io_ins_462, // @[:@143695.4]
  input  [63:0] io_ins_463, // @[:@143695.4]
  input  [63:0] io_ins_464, // @[:@143695.4]
  input  [63:0] io_ins_465, // @[:@143695.4]
  input  [63:0] io_ins_466, // @[:@143695.4]
  input  [63:0] io_ins_467, // @[:@143695.4]
  input  [63:0] io_ins_468, // @[:@143695.4]
  input  [63:0] io_ins_469, // @[:@143695.4]
  input  [63:0] io_ins_470, // @[:@143695.4]
  input  [63:0] io_ins_471, // @[:@143695.4]
  input  [63:0] io_ins_472, // @[:@143695.4]
  input  [63:0] io_ins_473, // @[:@143695.4]
  input  [63:0] io_ins_474, // @[:@143695.4]
  input  [63:0] io_ins_475, // @[:@143695.4]
  input  [63:0] io_ins_476, // @[:@143695.4]
  input  [63:0] io_ins_477, // @[:@143695.4]
  input  [63:0] io_ins_478, // @[:@143695.4]
  input  [63:0] io_ins_479, // @[:@143695.4]
  input  [63:0] io_ins_480, // @[:@143695.4]
  input  [63:0] io_ins_481, // @[:@143695.4]
  input  [63:0] io_ins_482, // @[:@143695.4]
  input  [63:0] io_ins_483, // @[:@143695.4]
  input  [63:0] io_ins_484, // @[:@143695.4]
  input  [63:0] io_ins_485, // @[:@143695.4]
  input  [63:0] io_ins_486, // @[:@143695.4]
  input  [63:0] io_ins_487, // @[:@143695.4]
  input  [63:0] io_ins_488, // @[:@143695.4]
  input  [63:0] io_ins_489, // @[:@143695.4]
  input  [63:0] io_ins_490, // @[:@143695.4]
  input  [63:0] io_ins_491, // @[:@143695.4]
  input  [63:0] io_ins_492, // @[:@143695.4]
  input  [63:0] io_ins_493, // @[:@143695.4]
  input  [63:0] io_ins_494, // @[:@143695.4]
  input  [63:0] io_ins_495, // @[:@143695.4]
  input  [63:0] io_ins_496, // @[:@143695.4]
  input  [63:0] io_ins_497, // @[:@143695.4]
  input  [63:0] io_ins_498, // @[:@143695.4]
  input  [63:0] io_ins_499, // @[:@143695.4]
  input  [63:0] io_ins_500, // @[:@143695.4]
  input  [63:0] io_ins_501, // @[:@143695.4]
  input  [63:0] io_ins_502, // @[:@143695.4]
  input  [8:0]  io_sel, // @[:@143695.4]
  output [63:0] io_out // @[:@143695.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@143697.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@143697.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@143697.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@143697.4]
endmodule
module RegFile( // @[:@143699.2]
  input         clock, // @[:@143700.4]
  input         reset, // @[:@143701.4]
  input  [31:0] io_raddr, // @[:@143702.4]
  input         io_wen, // @[:@143702.4]
  input  [31:0] io_waddr, // @[:@143702.4]
  input  [63:0] io_wdata, // @[:@143702.4]
  output [63:0] io_rdata, // @[:@143702.4]
  input         io_reset, // @[:@143702.4]
  output [63:0] io_argIns_0, // @[:@143702.4]
  output [63:0] io_argIns_1, // @[:@143702.4]
  output [63:0] io_argIns_2, // @[:@143702.4]
  output [63:0] io_argIns_3, // @[:@143702.4]
  input         io_argOuts_0_valid, // @[:@143702.4]
  input  [63:0] io_argOuts_0_bits, // @[:@143702.4]
  input         io_argOuts_1_valid, // @[:@143702.4]
  input  [63:0] io_argOuts_1_bits // @[:@143702.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@145712.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@145712.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@145712.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@145712.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@145712.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@145712.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@145724.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@145724.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@145724.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@145724.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@145724.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@145724.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@145743.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@145743.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@145743.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@145743.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@145743.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@145743.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@145755.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@145755.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@145767.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@145767.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@145767.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@145767.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@145767.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@145767.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@145781.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@145781.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@145781.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@145781.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@145781.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@145781.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@145795.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@145795.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@145795.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@145795.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@145795.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@145795.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@145809.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@145809.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@145809.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@145809.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@145809.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@145809.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@145823.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@145823.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@145823.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@145823.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@145823.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@145823.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@145837.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@145837.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@145837.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@145837.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@145837.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@145837.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@145851.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@145851.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@145851.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@145851.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@145851.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@145851.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@145865.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@145865.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@145865.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@145865.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@145865.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@145865.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@145879.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@145879.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@145879.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@145879.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@145879.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@145879.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@145893.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@145893.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@145893.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@145893.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@145893.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@145893.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@145907.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@145907.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@145907.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@145907.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@145907.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@145907.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@145921.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@145921.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@145921.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@145921.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@145921.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@145921.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@145935.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@145935.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@145935.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@145935.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@145935.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@145935.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@145949.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@145949.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@145949.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@145949.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@145949.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@145949.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@145963.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@145963.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@145963.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@145963.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@145963.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@145963.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@145977.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@145977.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@145977.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@145977.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@145977.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@145977.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@145991.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@145991.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@145991.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@145991.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@145991.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@145991.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@146005.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@146005.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@146005.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@146005.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@146005.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@146005.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@146019.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@146019.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@146019.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@146019.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@146019.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@146019.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@146033.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@146033.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@146033.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@146033.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@146033.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@146033.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@146047.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@146047.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@146047.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@146047.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@146047.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@146047.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@146061.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@146061.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@146061.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@146061.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@146061.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@146061.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@146075.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@146075.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@146075.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@146075.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@146075.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@146075.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@146089.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@146089.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@146089.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@146089.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@146089.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@146089.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@146103.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@146103.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@146103.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@146103.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@146103.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@146103.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@146117.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@146117.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@146117.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@146117.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@146117.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@146117.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@146131.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@146131.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@146131.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@146131.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@146131.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@146131.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@146145.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@146145.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@146145.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@146145.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@146145.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@146145.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@146159.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@146159.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@146159.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@146159.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@146159.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@146159.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@146173.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@146173.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@146173.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@146173.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@146173.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@146173.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@146187.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@146187.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@146187.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@146187.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@146187.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@146187.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@146201.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@146201.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@146201.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@146201.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@146201.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@146201.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@146215.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@146215.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@146215.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@146215.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@146215.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@146215.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@146229.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@146229.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@146229.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@146229.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@146229.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@146229.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@146243.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@146243.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@146243.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@146243.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@146243.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@146243.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@146257.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@146257.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@146257.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@146257.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@146257.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@146257.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@146271.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@146271.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@146271.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@146271.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@146271.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@146271.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@146285.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@146285.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@146285.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@146285.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@146285.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@146285.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@146299.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@146299.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@146299.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@146299.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@146299.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@146299.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@146313.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@146313.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@146313.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@146313.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@146313.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@146313.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@146327.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@146327.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@146327.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@146327.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@146327.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@146327.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@146341.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@146341.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@146341.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@146341.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@146341.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@146341.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@146355.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@146355.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@146355.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@146355.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@146355.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@146355.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@146369.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@146369.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@146369.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@146369.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@146369.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@146369.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@146383.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@146383.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@146383.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@146383.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@146383.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@146383.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@146397.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@146397.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@146397.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@146397.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@146397.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@146397.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@146411.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@146411.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@146411.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@146411.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@146411.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@146411.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@146425.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@146425.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@146425.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@146425.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@146425.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@146425.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@146439.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@146439.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@146439.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@146439.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@146439.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@146439.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@146453.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@146453.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@146453.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@146453.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@146453.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@146453.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@146467.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@146467.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@146467.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@146467.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@146467.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@146467.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@146481.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@146481.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@146481.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@146481.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@146481.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@146481.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@146495.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@146495.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@146495.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@146495.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@146495.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@146495.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@146509.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@146509.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@146509.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@146509.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@146509.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@146509.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@146523.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@146523.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@146523.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@146523.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@146523.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@146523.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@146537.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@146537.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@146537.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@146537.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@146537.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@146537.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@146551.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@146551.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@146551.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@146551.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@146551.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@146551.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@146565.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@146565.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@146565.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@146565.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@146565.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@146565.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@146579.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@146579.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@146579.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@146579.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@146579.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@146579.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@146593.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@146593.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@146593.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@146593.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@146593.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@146593.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@146607.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@146607.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@146607.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@146607.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@146607.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@146607.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@146621.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@146621.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@146621.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@146621.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@146621.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@146621.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@146635.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@146635.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@146635.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@146635.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@146635.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@146635.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@146649.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@146649.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@146649.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@146649.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@146649.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@146649.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@146663.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@146663.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@146663.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@146663.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@146663.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@146663.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@146677.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@146677.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@146677.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@146677.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@146677.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@146677.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@146691.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@146691.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@146691.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@146691.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@146691.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@146691.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@146705.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@146705.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@146705.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@146705.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@146705.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@146705.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@146719.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@146719.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@146719.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@146719.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@146719.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@146719.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@146733.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@146733.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@146733.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@146733.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@146733.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@146733.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@146747.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@146747.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@146747.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@146747.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@146747.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@146747.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@146761.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@146761.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@146761.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@146761.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@146761.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@146761.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@146775.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@146775.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@146775.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@146775.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@146775.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@146775.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@146789.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@146789.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@146789.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@146789.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@146789.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@146789.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@146803.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@146803.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@146803.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@146803.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@146803.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@146803.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@146817.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@146817.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@146817.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@146817.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@146817.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@146817.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@146831.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@146831.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@146831.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@146831.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@146831.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@146831.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@146845.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@146845.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@146845.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@146845.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@146845.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@146845.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@146859.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@146859.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@146859.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@146859.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@146859.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@146859.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@146873.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@146873.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@146873.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@146873.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@146873.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@146873.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@146887.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@146887.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@146887.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@146887.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@146887.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@146887.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@146901.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@146901.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@146901.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@146901.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@146901.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@146901.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@146915.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@146915.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@146915.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@146915.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@146915.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@146915.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@146929.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@146929.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@146929.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@146929.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@146929.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@146929.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@146943.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@146943.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@146943.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@146943.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@146943.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@146943.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@146957.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@146957.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@146957.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@146957.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@146957.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@146957.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@146971.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@146971.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@146971.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@146971.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@146971.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@146971.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@146985.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@146985.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@146985.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@146985.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@146985.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@146985.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@146999.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@146999.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@146999.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@146999.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@146999.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@146999.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@147013.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@147013.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@147013.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@147013.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@147013.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@147013.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@147027.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@147027.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@147027.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@147027.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@147027.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@147027.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@147041.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@147041.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@147041.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@147041.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@147041.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@147041.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@147055.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@147055.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@147055.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@147055.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@147055.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@147055.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@147069.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@147069.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@147069.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@147069.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@147069.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@147069.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@147083.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@147083.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@147083.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@147083.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@147083.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@147083.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@147097.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@147097.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@147097.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@147097.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@147097.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@147097.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@147111.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@147111.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@147111.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@147111.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@147111.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@147111.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@147125.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@147125.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@147125.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@147125.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@147125.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@147125.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@147139.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@147139.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@147139.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@147139.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@147139.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@147139.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@147153.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@147153.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@147153.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@147153.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@147153.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@147153.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@147167.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@147167.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@147167.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@147167.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@147167.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@147167.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@147181.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@147181.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@147181.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@147181.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@147181.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@147181.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@147195.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@147195.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@147195.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@147195.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@147195.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@147195.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@147209.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@147209.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@147209.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@147209.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@147209.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@147209.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@147223.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@147223.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@147223.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@147223.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@147223.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@147223.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@147237.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@147237.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@147237.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@147237.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@147237.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@147237.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@147251.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@147251.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@147251.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@147251.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@147251.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@147251.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@147265.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@147265.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@147265.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@147265.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@147265.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@147265.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@147279.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@147279.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@147279.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@147279.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@147279.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@147279.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@147293.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@147293.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@147293.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@147293.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@147293.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@147293.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@147307.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@147307.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@147307.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@147307.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@147307.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@147307.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@147321.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@147321.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@147321.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@147321.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@147321.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@147321.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@147335.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@147335.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@147335.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@147335.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@147335.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@147335.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@147349.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@147349.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@147349.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@147349.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@147349.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@147349.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@147363.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@147363.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@147363.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@147363.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@147363.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@147363.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@147377.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@147377.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@147377.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@147377.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@147377.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@147377.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@147391.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@147391.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@147391.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@147391.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@147391.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@147391.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@147405.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@147405.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@147405.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@147405.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@147405.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@147405.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@147419.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@147419.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@147419.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@147419.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@147419.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@147419.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@147433.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@147433.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@147433.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@147433.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@147433.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@147433.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@147447.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@147447.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@147447.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@147447.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@147447.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@147447.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@147461.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@147461.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@147461.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@147461.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@147461.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@147461.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@147475.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@147475.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@147475.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@147475.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@147475.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@147475.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@147489.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@147489.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@147489.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@147489.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@147489.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@147489.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@147503.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@147503.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@147503.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@147503.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@147503.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@147503.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@147517.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@147517.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@147517.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@147517.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@147517.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@147517.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@147531.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@147531.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@147531.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@147531.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@147531.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@147531.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@147545.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@147545.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@147545.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@147545.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@147545.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@147545.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@147559.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@147559.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@147559.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@147559.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@147559.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@147559.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@147573.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@147573.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@147573.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@147573.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@147573.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@147573.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@147587.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@147587.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@147587.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@147587.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@147587.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@147587.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@147601.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@147601.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@147601.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@147601.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@147601.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@147601.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@147615.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@147615.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@147615.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@147615.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@147615.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@147615.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@147629.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@147629.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@147629.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@147629.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@147629.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@147629.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@147643.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@147643.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@147643.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@147643.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@147643.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@147643.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@147657.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@147657.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@147657.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@147657.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@147657.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@147657.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@147671.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@147671.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@147671.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@147671.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@147671.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@147671.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@147685.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@147685.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@147685.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@147685.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@147685.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@147685.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@147699.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@147699.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@147699.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@147699.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@147699.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@147699.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@147713.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@147713.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@147713.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@147713.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@147713.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@147713.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@147727.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@147727.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@147727.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@147727.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@147727.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@147727.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@147741.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@147741.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@147741.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@147741.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@147741.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@147741.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@147755.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@147755.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@147755.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@147755.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@147755.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@147755.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@147769.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@147769.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@147769.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@147769.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@147769.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@147769.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@147783.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@147783.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@147783.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@147783.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@147783.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@147783.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@147797.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@147797.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@147797.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@147797.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@147797.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@147797.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@147811.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@147811.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@147811.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@147811.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@147811.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@147811.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@147825.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@147825.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@147825.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@147825.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@147825.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@147825.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@147839.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@147839.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@147839.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@147839.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@147839.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@147839.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@147853.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@147853.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@147853.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@147853.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@147853.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@147853.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@147867.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@147867.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@147867.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@147867.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@147867.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@147867.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@147881.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@147881.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@147881.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@147881.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@147881.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@147881.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@147895.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@147895.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@147895.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@147895.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@147895.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@147895.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@147909.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@147909.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@147909.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@147909.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@147909.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@147909.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@147923.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@147923.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@147923.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@147923.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@147923.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@147923.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@147937.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@147937.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@147937.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@147937.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@147937.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@147937.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@147951.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@147951.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@147951.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@147951.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@147951.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@147951.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@147965.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@147965.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@147965.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@147965.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@147965.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@147965.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@147979.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@147979.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@147979.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@147979.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@147979.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@147979.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@147993.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@147993.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@147993.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@147993.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@147993.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@147993.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@148007.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@148007.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@148007.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@148007.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@148007.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@148007.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@148021.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@148021.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@148021.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@148021.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@148021.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@148021.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@148035.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@148035.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@148035.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@148035.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@148035.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@148035.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@148049.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@148049.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@148049.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@148049.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@148049.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@148049.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@148063.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@148063.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@148063.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@148063.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@148063.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@148063.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@148077.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@148077.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@148077.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@148077.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@148077.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@148077.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@148091.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@148091.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@148091.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@148091.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@148091.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@148091.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@148105.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@148105.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@148105.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@148105.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@148105.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@148105.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@148119.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@148119.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@148119.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@148119.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@148119.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@148119.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@148133.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@148133.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@148133.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@148133.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@148133.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@148133.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@148147.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@148147.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@148147.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@148147.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@148147.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@148147.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@148161.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@148161.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@148161.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@148161.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@148161.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@148161.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@148175.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@148175.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@148175.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@148175.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@148175.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@148175.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@148189.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@148189.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@148189.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@148189.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@148189.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@148189.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@148203.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@148203.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@148203.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@148203.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@148203.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@148203.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@148217.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@148217.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@148217.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@148217.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@148217.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@148217.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@148231.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@148231.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@148231.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@148231.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@148231.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@148231.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@148245.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@148245.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@148245.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@148245.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@148245.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@148245.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@148259.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@148259.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@148259.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@148259.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@148259.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@148259.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@148273.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@148273.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@148273.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@148273.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@148273.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@148273.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@148287.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@148287.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@148287.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@148287.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@148287.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@148287.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@148301.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@148301.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@148301.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@148301.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@148301.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@148301.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@148315.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@148315.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@148315.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@148315.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@148315.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@148315.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@148329.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@148329.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@148329.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@148329.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@148329.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@148329.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@148343.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@148343.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@148343.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@148343.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@148343.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@148343.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@148357.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@148357.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@148357.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@148357.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@148357.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@148357.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@148371.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@148371.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@148371.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@148371.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@148371.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@148371.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@148385.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@148385.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@148385.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@148385.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@148385.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@148385.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@148399.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@148399.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@148399.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@148399.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@148399.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@148399.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@148413.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@148413.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@148413.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@148413.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@148413.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@148413.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@148427.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@148427.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@148427.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@148427.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@148427.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@148427.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@148441.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@148441.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@148441.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@148441.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@148441.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@148441.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@148455.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@148455.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@148455.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@148455.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@148455.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@148455.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@148469.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@148469.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@148469.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@148469.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@148469.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@148469.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@148483.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@148483.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@148483.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@148483.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@148483.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@148483.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@148497.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@148497.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@148497.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@148497.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@148497.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@148497.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@148511.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@148511.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@148511.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@148511.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@148511.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@148511.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@148525.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@148525.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@148525.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@148525.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@148525.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@148525.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@148539.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@148539.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@148539.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@148539.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@148539.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@148539.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@148553.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@148553.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@148553.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@148553.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@148553.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@148553.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@148567.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@148567.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@148567.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@148567.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@148567.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@148567.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@148581.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@148581.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@148581.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@148581.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@148581.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@148581.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@148595.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@148595.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@148595.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@148595.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@148595.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@148595.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@148609.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@148609.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@148609.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@148609.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@148609.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@148609.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@148623.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@148623.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@148623.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@148623.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@148623.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@148623.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@148637.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@148637.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@148637.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@148637.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@148637.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@148637.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@148651.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@148651.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@148651.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@148651.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@148651.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@148651.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@148665.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@148665.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@148665.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@148665.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@148665.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@148665.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@148679.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@148679.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@148679.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@148679.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@148679.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@148679.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@148693.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@148693.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@148693.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@148693.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@148693.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@148693.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@148707.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@148707.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@148707.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@148707.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@148707.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@148707.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@148721.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@148721.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@148721.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@148721.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@148721.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@148721.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@148735.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@148735.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@148735.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@148735.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@148735.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@148735.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@148749.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@148749.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@148749.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@148749.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@148749.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@148749.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@148763.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@148763.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@148763.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@148763.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@148763.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@148763.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@148777.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@148777.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@148777.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@148777.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@148777.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@148777.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@148791.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@148791.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@148791.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@148791.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@148791.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@148791.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@148805.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@148805.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@148805.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@148805.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@148805.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@148805.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@148819.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@148819.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@148819.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@148819.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@148819.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@148819.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@148833.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@148833.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@148833.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@148833.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@148833.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@148833.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@148847.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@148847.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@148847.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@148847.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@148847.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@148847.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@148861.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@148861.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@148861.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@148861.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@148861.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@148861.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@148875.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@148875.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@148875.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@148875.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@148875.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@148875.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@148889.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@148889.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@148889.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@148889.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@148889.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@148889.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@148903.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@148903.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@148903.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@148903.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@148903.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@148903.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@148917.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@148917.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@148917.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@148917.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@148917.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@148917.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@148931.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@148931.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@148931.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@148931.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@148931.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@148931.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@148945.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@148945.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@148945.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@148945.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@148945.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@148945.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@148959.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@148959.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@148959.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@148959.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@148959.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@148959.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@148973.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@148973.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@148973.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@148973.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@148973.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@148973.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@148987.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@148987.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@148987.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@148987.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@148987.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@148987.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@149001.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@149001.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@149001.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@149001.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@149001.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@149001.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@149015.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@149015.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@149015.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@149015.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@149015.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@149015.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@149029.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@149029.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@149029.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@149029.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@149029.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@149029.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@149043.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@149043.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@149043.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@149043.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@149043.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@149043.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@149057.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@149057.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@149057.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@149057.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@149057.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@149057.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@149071.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@149071.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@149071.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@149071.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@149071.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@149071.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@149085.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@149085.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@149085.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@149085.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@149085.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@149085.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@149099.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@149099.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@149099.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@149099.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@149099.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@149099.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@149113.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@149113.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@149113.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@149113.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@149113.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@149113.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@149127.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@149127.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@149127.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@149127.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@149127.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@149127.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@149141.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@149141.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@149141.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@149141.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@149141.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@149141.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@149155.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@149155.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@149155.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@149155.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@149155.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@149155.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@149169.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@149169.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@149169.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@149169.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@149169.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@149169.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@149183.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@149183.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@149183.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@149183.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@149183.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@149183.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@149197.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@149197.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@149197.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@149197.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@149197.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@149197.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@149211.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@149211.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@149211.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@149211.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@149211.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@149211.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@149225.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@149225.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@149225.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@149225.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@149225.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@149225.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@149239.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@149239.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@149239.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@149239.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@149239.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@149239.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@149253.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@149253.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@149253.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@149253.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@149253.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@149253.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@149267.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@149267.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@149267.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@149267.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@149267.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@149267.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@149281.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@149281.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@149281.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@149281.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@149281.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@149281.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@149295.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@149295.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@149295.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@149295.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@149295.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@149295.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@149309.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@149309.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@149309.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@149309.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@149309.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@149309.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@149323.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@149323.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@149323.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@149323.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@149323.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@149323.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@149337.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@149337.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@149337.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@149337.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@149337.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@149337.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@149351.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@149351.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@149351.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@149351.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@149351.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@149351.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@149365.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@149365.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@149365.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@149365.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@149365.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@149365.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@149379.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@149379.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@149379.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@149379.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@149379.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@149379.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@149393.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@149393.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@149393.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@149393.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@149393.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@149393.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@149407.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@149407.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@149407.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@149407.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@149407.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@149407.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@149421.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@149421.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@149421.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@149421.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@149421.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@149421.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@149435.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@149435.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@149435.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@149435.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@149435.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@149435.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@149449.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@149449.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@149449.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@149449.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@149449.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@149449.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@149463.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@149463.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@149463.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@149463.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@149463.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@149463.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@149477.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@149477.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@149477.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@149477.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@149477.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@149477.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@149491.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@149491.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@149491.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@149491.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@149491.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@149491.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@149505.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@149505.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@149505.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@149505.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@149505.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@149505.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@149519.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@149519.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@149519.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@149519.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@149519.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@149519.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@149533.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@149533.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@149533.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@149533.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@149533.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@149533.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@149547.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@149547.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@149547.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@149547.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@149547.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@149547.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@149561.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@149561.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@149561.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@149561.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@149561.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@149561.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@149575.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@149575.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@149575.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@149575.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@149575.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@149575.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@149589.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@149589.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@149589.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@149589.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@149589.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@149589.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@149603.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@149603.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@149603.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@149603.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@149603.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@149603.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@149617.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@149617.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@149617.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@149617.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@149617.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@149617.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@149631.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@149631.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@149631.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@149631.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@149631.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@149631.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@149645.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@149645.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@149645.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@149645.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@149645.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@149645.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@149659.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@149659.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@149659.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@149659.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@149659.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@149659.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@149673.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@149673.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@149673.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@149673.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@149673.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@149673.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@149687.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@149687.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@149687.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@149687.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@149687.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@149687.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@149701.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@149701.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@149701.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@149701.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@149701.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@149701.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@149715.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@149715.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@149715.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@149715.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@149715.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@149715.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@149729.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@149729.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@149729.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@149729.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@149729.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@149729.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@149743.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@149743.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@149743.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@149743.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@149743.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@149743.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@149757.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@149757.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@149757.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@149757.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@149757.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@149757.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@149771.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@149771.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@149771.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@149771.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@149771.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@149771.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@149785.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@149785.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@149785.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@149785.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@149785.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@149785.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@149799.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@149799.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@149799.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@149799.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@149799.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@149799.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@149813.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@149813.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@149813.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@149813.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@149813.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@149813.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@149827.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@149827.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@149827.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@149827.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@149827.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@149827.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@149841.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@149841.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@149841.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@149841.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@149841.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@149841.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@149855.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@149855.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@149855.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@149855.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@149855.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@149855.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@149869.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@149869.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@149869.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@149869.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@149869.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@149869.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@149883.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@149883.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@149883.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@149883.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@149883.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@149883.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@149897.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@149897.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@149897.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@149897.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@149897.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@149897.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@149911.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@149911.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@149911.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@149911.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@149911.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@149911.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@149925.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@149925.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@149925.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@149925.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@149925.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@149925.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@149939.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@149939.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@149939.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@149939.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@149939.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@149939.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@149953.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@149953.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@149953.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@149953.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@149953.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@149953.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@149967.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@149967.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@149967.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@149967.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@149967.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@149967.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@149981.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@149981.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@149981.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@149981.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@149981.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@149981.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@149995.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@149995.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@149995.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@149995.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@149995.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@149995.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@150009.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@150009.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@150009.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@150009.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@150009.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@150009.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@150023.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@150023.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@150023.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@150023.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@150023.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@150023.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@150037.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@150037.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@150037.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@150037.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@150037.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@150037.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@150051.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@150051.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@150051.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@150051.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@150051.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@150051.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@150065.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@150065.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@150065.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@150065.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@150065.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@150065.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@150079.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@150079.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@150079.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@150079.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@150079.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@150079.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@150093.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@150093.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@150093.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@150093.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@150093.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@150093.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@150107.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@150107.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@150107.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@150107.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@150107.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@150107.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@150121.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@150121.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@150121.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@150121.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@150121.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@150121.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@150135.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@150135.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@150135.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@150135.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@150135.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@150135.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@150149.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@150149.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@150149.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@150149.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@150149.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@150149.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@150163.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@150163.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@150163.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@150163.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@150163.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@150163.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@150177.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@150177.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@150177.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@150177.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@150177.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@150177.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@150191.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@150191.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@150191.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@150191.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@150191.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@150191.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@150205.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@150205.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@150205.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@150205.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@150205.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@150205.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@150219.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@150219.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@150219.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@150219.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@150219.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@150219.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@150233.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@150233.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@150233.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@150233.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@150233.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@150233.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@150247.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@150247.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@150247.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@150247.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@150247.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@150247.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@150261.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@150261.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@150261.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@150261.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@150261.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@150261.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@150275.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@150275.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@150275.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@150275.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@150275.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@150275.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@150289.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@150289.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@150289.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@150289.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@150289.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@150289.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@150303.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@150303.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@150303.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@150303.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@150303.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@150303.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@150317.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@150317.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@150317.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@150317.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@150317.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@150317.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@150331.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@150331.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@150331.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@150331.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@150331.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@150331.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@150345.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@150345.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@150345.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@150345.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@150345.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@150345.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@150359.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@150359.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@150359.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@150359.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@150359.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@150359.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@150373.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@150373.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@150373.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@150373.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@150373.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@150373.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@150387.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@150387.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@150387.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@150387.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@150387.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@150387.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@150401.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@150401.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@150401.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@150401.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@150401.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@150401.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@150415.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@150415.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@150415.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@150415.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@150415.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@150415.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@150429.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@150429.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@150429.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@150429.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@150429.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@150429.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@150443.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@150443.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@150443.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@150443.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@150443.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@150443.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@150457.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@150457.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@150457.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@150457.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@150457.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@150457.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@150471.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@150471.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@150471.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@150471.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@150471.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@150471.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@150485.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@150485.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@150485.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@150485.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@150485.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@150485.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@150499.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@150499.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@150499.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@150499.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@150499.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@150499.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@150513.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@150513.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@150513.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@150513.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@150513.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@150513.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@150527.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@150527.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@150527.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@150527.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@150527.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@150527.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@150541.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@150541.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@150541.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@150541.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@150541.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@150541.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@150555.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@150555.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@150555.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@150555.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@150555.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@150555.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@150569.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@150569.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@150569.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@150569.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@150569.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@150569.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@150583.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@150583.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@150583.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@150583.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@150583.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@150583.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@150597.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@150597.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@150597.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@150597.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@150597.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@150597.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@150611.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@150611.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@150611.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@150611.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@150611.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@150611.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@150625.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@150625.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@150625.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@150625.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@150625.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@150625.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@150639.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@150639.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@150639.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@150639.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@150639.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@150639.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@150653.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@150653.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@150653.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@150653.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@150653.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@150653.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@150667.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@150667.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@150667.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@150667.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@150667.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@150667.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@150681.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@150681.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@150681.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@150681.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@150681.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@150681.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@150695.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@150695.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@150695.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@150695.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@150695.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@150695.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@150709.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@150709.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@150709.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@150709.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@150709.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@150709.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@150723.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@150723.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@150723.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@150723.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@150723.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@150723.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@150737.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@150737.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@150737.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@150737.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@150737.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@150737.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@150751.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@150751.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@150751.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@150751.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@150751.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@150751.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@150765.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@150765.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@150765.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@150765.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@150765.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@150765.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@150779.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@150779.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@150779.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@150779.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@150779.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@150779.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@150793.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@150793.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@150793.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@150793.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@150793.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@150793.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@150807.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@150807.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@150807.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@150807.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@150807.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@150807.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@150821.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@150821.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@150821.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@150821.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@150821.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@150821.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@150835.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@150835.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@150835.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@150835.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@150835.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@150835.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@150849.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@150849.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@150849.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@150849.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@150849.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@150849.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@150863.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@150863.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@150863.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@150863.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@150863.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@150863.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@150877.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@150877.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@150877.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@150877.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@150877.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@150877.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@150891.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@150891.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@150891.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@150891.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@150891.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@150891.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@150905.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@150905.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@150905.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@150905.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@150905.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@150905.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@150919.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@150919.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@150919.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@150919.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@150919.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@150919.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@150933.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@150933.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@150933.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@150933.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@150933.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@150933.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@150947.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@150947.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@150947.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@150947.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@150947.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@150947.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@150961.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@150961.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@150961.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@150961.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@150961.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@150961.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@150975.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@150975.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@150975.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@150975.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@150975.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@150975.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@150989.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@150989.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@150989.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@150989.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@150989.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@150989.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@151003.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@151003.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@151003.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@151003.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@151003.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@151003.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@151017.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@151017.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@151017.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@151017.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@151017.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@151017.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@151031.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@151031.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@151031.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@151031.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@151031.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@151031.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@151045.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@151045.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@151045.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@151045.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@151045.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@151045.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@151059.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@151059.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@151059.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@151059.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@151059.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@151059.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@151073.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@151073.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@151073.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@151073.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@151073.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@151073.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@151087.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@151087.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@151087.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@151087.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@151087.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@151087.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@151101.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@151101.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@151101.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@151101.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@151101.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@151101.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@151115.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@151115.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@151115.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@151115.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@151115.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@151115.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@151129.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@151129.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@151129.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@151129.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@151129.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@151129.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@151143.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@151143.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@151143.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@151143.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@151143.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@151143.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@151157.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@151157.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@151157.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@151157.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@151157.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@151157.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@151171.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@151171.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@151171.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@151171.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@151171.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@151171.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@151185.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@151185.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@151185.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@151185.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@151185.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@151185.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@151199.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@151199.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@151199.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@151199.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@151199.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@151199.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@151213.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@151213.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@151213.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@151213.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@151213.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@151213.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@151227.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@151227.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@151227.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@151227.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@151227.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@151227.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@151241.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@151241.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@151241.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@151241.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@151241.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@151241.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@151255.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@151255.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@151255.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@151255.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@151255.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@151255.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@151269.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@151269.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@151269.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@151269.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@151269.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@151269.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@151283.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@151283.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@151283.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@151283.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@151283.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@151283.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@151297.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@151297.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@151297.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@151297.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@151297.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@151297.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@151311.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@151311.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@151311.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@151311.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@151311.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@151311.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@151325.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@151325.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@151325.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@151325.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@151325.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@151325.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@151339.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@151339.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@151339.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@151339.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@151339.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@151339.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@151353.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@151353.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@151353.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@151353.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@151353.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@151353.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@151367.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@151367.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@151367.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@151367.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@151367.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@151367.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@151381.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@151381.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@151381.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@151381.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@151381.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@151381.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@151395.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@151395.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@151395.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@151395.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@151395.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@151395.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@151409.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@151409.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@151409.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@151409.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@151409.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@151409.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@151423.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@151423.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@151423.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@151423.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@151423.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@151423.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@151437.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@151437.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@151437.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@151437.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@151437.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@151437.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@151451.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@151451.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@151451.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@151451.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@151451.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@151451.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@151465.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@151465.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@151465.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@151465.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@151465.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@151465.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@151479.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@151479.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@151479.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@151479.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@151479.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@151479.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@151493.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@151493.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@151493.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@151493.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@151493.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@151493.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@151507.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@151507.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@151507.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@151507.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@151507.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@151507.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@151521.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@151521.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@151521.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@151521.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@151521.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@151521.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@151535.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@151535.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@151535.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@151535.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@151535.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@151535.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@151549.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@151549.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@151549.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@151549.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@151549.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@151549.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@151563.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@151563.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@151563.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@151563.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@151563.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@151563.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@151577.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@151577.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@151577.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@151577.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@151577.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@151577.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@151591.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@151591.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@151591.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@151591.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@151591.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@151591.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@151605.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@151605.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@151605.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@151605.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@151605.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@151605.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@151619.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@151619.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@151619.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@151619.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@151619.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@151619.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@151633.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@151633.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@151633.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@151633.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@151633.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@151633.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@151647.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@151647.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@151647.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@151647.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@151647.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@151647.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@151661.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@151661.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@151661.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@151661.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@151661.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@151661.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@151675.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@151675.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@151675.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@151675.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@151675.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@151675.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@151689.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@151689.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@151689.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@151689.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@151689.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@151689.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@151703.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@151703.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@151703.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@151703.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@151703.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@151703.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@151717.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@151717.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@151717.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@151717.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@151717.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@151717.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@151731.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@151731.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@151731.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@151731.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@151731.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@151731.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@151745.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@151745.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@151745.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@151745.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@151745.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@151745.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@151759.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@151759.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@151759.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@151759.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@151759.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@151759.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@151773.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@151773.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@151773.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@151773.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@151773.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@151773.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@151787.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@151787.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@151787.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@151787.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@151787.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@151787.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@151801.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@151801.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@151801.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@151801.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@151801.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@151801.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@151815.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@151815.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@151815.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@151815.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@151815.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@151815.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@151829.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@151829.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@151829.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@151829.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@151829.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@151829.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@151843.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@151843.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@151843.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@151843.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@151843.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@151843.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@151857.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@151857.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@151857.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@151857.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@151857.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@151857.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@151871.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@151871.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@151871.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@151871.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@151871.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@151871.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@151885.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@151885.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@151885.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@151885.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@151885.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@151885.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@151899.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@151899.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@151899.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@151899.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@151899.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@151899.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@151913.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@151913.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@151913.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@151913.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@151913.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@151913.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@151927.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@151927.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@151927.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@151927.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@151927.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@151927.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@151941.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@151941.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@151941.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@151941.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@151941.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@151941.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@151955.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@151955.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@151955.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@151955.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@151955.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@151955.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@151969.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@151969.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@151969.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@151969.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@151969.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@151969.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@151983.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@151983.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@151983.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@151983.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@151983.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@151983.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@151997.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@151997.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@151997.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@151997.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@151997.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@151997.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@152011.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@152011.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@152011.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@152011.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@152011.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@152011.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@152025.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@152025.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@152025.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@152025.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@152025.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@152025.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@152039.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@152039.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@152039.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@152039.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@152039.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@152039.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@152053.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@152053.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@152053.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@152053.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@152053.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@152053.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@152067.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@152067.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@152067.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@152067.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@152067.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@152067.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@152081.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@152081.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@152081.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@152081.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@152081.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@152081.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@152095.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@152095.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@152095.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@152095.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@152095.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@152095.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@152109.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@152109.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@152109.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@152109.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@152109.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@152109.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@152123.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@152123.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@152123.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@152123.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@152123.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@152123.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@152137.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@152137.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@152137.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@152137.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@152137.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@152137.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@152151.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@152151.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@152151.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@152151.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@152151.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@152151.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@152165.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@152165.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@152165.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@152165.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@152165.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@152165.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@152179.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@152179.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@152179.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@152179.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@152179.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@152179.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@152193.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@152193.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@152193.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@152193.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@152193.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@152193.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@152207.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@152207.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@152207.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@152207.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@152207.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@152207.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@152221.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@152221.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@152221.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@152221.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@152221.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@152221.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@152235.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@152235.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@152235.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@152235.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@152235.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@152235.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@152249.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@152249.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@152249.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@152249.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@152249.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@152249.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@152263.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@152263.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@152263.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@152263.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@152263.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@152263.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@152277.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@152277.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@152277.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@152277.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@152277.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@152277.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@152291.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@152291.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@152291.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@152291.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@152291.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@152291.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@152305.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@152305.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@152305.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@152305.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@152305.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@152305.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@152319.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@152319.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@152319.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@152319.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@152319.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@152319.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@152333.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@152333.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@152333.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@152333.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@152333.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@152333.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@152347.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@152347.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@152347.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@152347.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@152347.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@152347.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@152361.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@152361.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@152361.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@152361.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@152361.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@152361.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@152375.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@152375.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@152375.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@152375.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@152375.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@152375.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@152389.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@152389.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@152389.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@152389.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@152389.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@152389.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@152403.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@152403.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@152403.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@152403.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@152403.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@152403.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@152417.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@152417.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@152417.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@152417.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@152417.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@152417.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@152431.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@152431.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@152431.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@152431.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@152431.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@152431.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@152445.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@152445.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@152445.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@152445.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@152445.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@152445.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@152459.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@152459.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@152459.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@152459.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@152459.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@152459.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@152473.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@152473.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@152473.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@152473.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@152473.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@152473.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@152487.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@152487.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@152487.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@152487.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@152487.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@152487.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@152501.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@152501.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@152501.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@152501.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@152501.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@152501.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@152515.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@152515.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@152515.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@152515.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@152515.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@152515.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@152529.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@152529.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@152529.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@152529.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@152529.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@152529.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@152543.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@152543.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@152543.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@152543.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@152543.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@152543.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@152557.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@152557.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@152557.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@152557.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@152557.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@152557.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@152571.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@152571.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@152571.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@152571.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@152571.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@152571.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@152585.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@152585.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@152585.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@152585.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@152585.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@152585.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@152599.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@152599.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@152599.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@152599.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@152599.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@152599.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@152613.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@152613.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@152613.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@152613.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@152613.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@152613.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@152627.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@152627.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@152627.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@152627.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@152627.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@152627.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@152641.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@152641.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@152641.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@152641.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@152641.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@152641.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@152655.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@152655.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@152655.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@152655.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@152655.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@152655.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@152669.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@152669.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@152669.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@152669.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@152669.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@152669.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@152683.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@152683.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@152683.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@152683.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@152683.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@152683.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@152697.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@152697.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@152697.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@152697.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@152697.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@152697.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@152711.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@152711.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@152711.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@152711.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@152711.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@152711.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@152725.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@152725.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@152725.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@152725.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@152725.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@152725.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@152739.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@152739.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@152739.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@152739.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@152739.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@152739.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@152753.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@152753.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@152753.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@145715.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@145727.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@145728.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@145746.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@145758.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@145770.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@145771.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@145712.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@145724.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@145743.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@145755.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@145767.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@145781.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@145795.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@145809.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@145823.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@145837.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@145851.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@145865.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@145879.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@145893.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@145907.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@145921.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@145935.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@145949.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@145963.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@145977.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@145991.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@146005.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@146019.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@146033.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@146047.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@146061.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@146075.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@146089.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@146103.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@146117.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@146131.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@146145.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@146159.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@146173.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@146187.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@146201.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@146215.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@146229.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@146243.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@146257.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@146271.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@146285.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@146299.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@146313.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@146327.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@146341.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@146355.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@146369.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@146383.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@146397.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@146411.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@146425.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@146439.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@146453.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@146467.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@146481.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@146495.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@146509.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@146523.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@146537.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@146551.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@146565.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@146579.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@146593.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@146607.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@146621.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@146635.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@146649.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@146663.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@146677.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@146691.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@146705.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@146719.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@146733.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@146747.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@146761.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@146775.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@146789.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@146803.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@146817.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@146831.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@146845.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@146859.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@146873.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@146887.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@146901.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@146915.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@146929.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@146943.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@146957.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@146971.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@146985.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@146999.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@147013.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@147027.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@147041.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@147055.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@147069.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@147083.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@147097.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@147111.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@147125.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@147139.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@147153.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@147167.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@147181.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@147195.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@147209.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@147223.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@147237.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@147251.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@147265.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@147279.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@147293.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@147307.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@147321.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@147335.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@147349.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@147363.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@147377.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@147391.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@147405.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@147419.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@147433.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@147447.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@147461.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@147475.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@147489.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@147503.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@147517.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@147531.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@147545.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@147559.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@147573.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@147587.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@147601.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@147615.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@147629.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@147643.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@147657.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@147671.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@147685.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@147699.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@147713.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@147727.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@147741.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@147755.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@147769.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@147783.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@147797.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@147811.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@147825.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@147839.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@147853.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@147867.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@147881.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@147895.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@147909.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@147923.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@147937.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@147951.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@147965.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@147979.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@147993.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@148007.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@148021.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@148035.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@148049.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@148063.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@148077.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@148091.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@148105.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@148119.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@148133.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@148147.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@148161.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@148175.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@148189.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@148203.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@148217.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@148231.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@148245.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@148259.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@148273.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@148287.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@148301.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@148315.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@148329.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@148343.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@148357.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@148371.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@148385.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@148399.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@148413.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@148427.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@148441.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@148455.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@148469.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@148483.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@148497.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@148511.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@148525.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@148539.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@148553.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@148567.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@148581.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@148595.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@148609.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@148623.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@148637.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@148651.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@148665.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@148679.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@148693.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@148707.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@148721.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@148735.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@148749.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@148763.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@148777.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@148791.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@148805.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@148819.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@148833.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@148847.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@148861.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@148875.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@148889.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@148903.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@148917.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@148931.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@148945.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@148959.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@148973.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@148987.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@149001.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@149015.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@149029.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@149043.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@149057.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@149071.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@149085.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@149099.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@149113.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@149127.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@149141.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@149155.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@149169.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@149183.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@149197.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@149211.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@149225.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@149239.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@149253.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@149267.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@149281.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@149295.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@149309.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@149323.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@149337.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@149351.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@149365.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@149379.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@149393.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@149407.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@149421.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@149435.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@149449.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@149463.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@149477.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@149491.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@149505.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@149519.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@149533.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@149547.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@149561.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@149575.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@149589.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@149603.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@149617.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@149631.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@149645.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@149659.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@149673.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@149687.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@149701.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@149715.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@149729.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@149743.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@149757.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@149771.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@149785.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@149799.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@149813.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@149827.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@149841.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@149855.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@149869.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@149883.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@149897.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@149911.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@149925.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@149939.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@149953.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@149967.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@149981.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@149995.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@150009.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@150023.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@150037.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@150051.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@150065.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@150079.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@150093.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@150107.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@150121.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@150135.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@150149.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@150163.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@150177.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@150191.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@150205.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@150219.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@150233.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@150247.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@150261.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@150275.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@150289.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@150303.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@150317.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@150331.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@150345.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@150359.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@150373.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@150387.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@150401.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@150415.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@150429.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@150443.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@150457.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@150471.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@150485.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@150499.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@150513.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@150527.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@150541.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@150555.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@150569.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@150583.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@150597.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@150611.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@150625.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@150639.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@150653.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@150667.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@150681.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@150695.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@150709.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@150723.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@150737.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@150751.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@150765.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@150779.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@150793.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@150807.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@150821.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@150835.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@150849.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@150863.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@150877.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@150891.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@150905.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@150919.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@150933.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@150947.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@150961.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@150975.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@150989.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@151003.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@151017.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@151031.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@151045.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@151059.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@151073.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@151087.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@151101.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@151115.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@151129.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@151143.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@151157.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@151171.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@151185.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@151199.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@151213.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@151227.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@151241.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@151255.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@151269.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@151283.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@151297.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@151311.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@151325.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@151339.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@151353.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@151367.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@151381.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@151395.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@151409.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@151423.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@151437.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@151451.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@151465.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@151479.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@151493.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@151507.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@151521.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@151535.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@151549.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@151563.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@151577.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@151591.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@151605.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@151619.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@151633.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@151647.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@151661.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@151675.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@151689.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@151703.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@151717.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@151731.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@151745.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@151759.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@151773.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@151787.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@151801.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@151815.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@151829.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@151843.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@151857.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@151871.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@151885.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@151899.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@151913.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@151927.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@151941.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@151955.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@151969.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@151983.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@151997.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@152011.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@152025.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@152039.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@152053.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@152067.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@152081.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@152095.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@152109.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@152123.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@152137.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@152151.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@152165.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@152179.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@152193.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@152207.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@152221.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@152235.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@152249.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@152263.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@152277.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@152291.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@152305.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@152319.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@152333.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@152347.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@152361.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@152375.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@152389.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@152403.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@152417.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@152431.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@152445.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@152459.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@152473.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@152487.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@152501.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@152515.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@152529.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@152543.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@152557.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@152571.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@152585.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@152599.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@152613.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@152627.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@152641.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@152655.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@152669.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@152683.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@152697.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@152711.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@152725.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@152739.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@152753.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@145715.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@145727.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@145728.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@145746.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@145758.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@145770.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@145771.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@153764.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@153770.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@153771.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@153772.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@153773.4]
  assign regs_0_clock = clock; // @[:@145713.4]
  assign regs_0_reset = reset; // @[:@145714.4 RegFile.scala 82:16:@145720.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@145718.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@145722.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@145717.4]
  assign regs_1_clock = clock; // @[:@145725.4]
  assign regs_1_reset = reset; // @[:@145726.4 RegFile.scala 70:16:@145738.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@145736.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@145741.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@145732.4]
  assign regs_2_clock = clock; // @[:@145744.4]
  assign regs_2_reset = reset; // @[:@145745.4 RegFile.scala 82:16:@145751.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@145749.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@145753.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@145748.4]
  assign regs_3_clock = clock; // @[:@145756.4]
  assign regs_3_reset = reset; // @[:@145757.4 RegFile.scala 82:16:@145763.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@145761.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@145765.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@145760.4]
  assign regs_4_clock = clock; // @[:@145768.4]
  assign regs_4_reset = io_reset; // @[:@145769.4 RegFile.scala 76:16:@145776.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@145775.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@145779.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@145773.4]
  assign regs_5_clock = clock; // @[:@145782.4]
  assign regs_5_reset = io_reset; // @[:@145783.4 RegFile.scala 76:16:@145790.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@145789.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@145793.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@145787.4]
  assign regs_6_clock = clock; // @[:@145796.4]
  assign regs_6_reset = io_reset; // @[:@145797.4 RegFile.scala 76:16:@145804.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@145803.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@145807.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@145801.4]
  assign regs_7_clock = clock; // @[:@145810.4]
  assign regs_7_reset = io_reset; // @[:@145811.4 RegFile.scala 76:16:@145818.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@145817.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@145821.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@145815.4]
  assign regs_8_clock = clock; // @[:@145824.4]
  assign regs_8_reset = io_reset; // @[:@145825.4 RegFile.scala 76:16:@145832.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@145831.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@145835.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@145829.4]
  assign regs_9_clock = clock; // @[:@145838.4]
  assign regs_9_reset = io_reset; // @[:@145839.4 RegFile.scala 76:16:@145846.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@145845.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@145849.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@145843.4]
  assign regs_10_clock = clock; // @[:@145852.4]
  assign regs_10_reset = io_reset; // @[:@145853.4 RegFile.scala 76:16:@145860.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@145859.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@145863.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@145857.4]
  assign regs_11_clock = clock; // @[:@145866.4]
  assign regs_11_reset = io_reset; // @[:@145867.4 RegFile.scala 76:16:@145874.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@145873.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@145877.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@145871.4]
  assign regs_12_clock = clock; // @[:@145880.4]
  assign regs_12_reset = io_reset; // @[:@145881.4 RegFile.scala 76:16:@145888.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@145887.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@145891.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@145885.4]
  assign regs_13_clock = clock; // @[:@145894.4]
  assign regs_13_reset = io_reset; // @[:@145895.4 RegFile.scala 76:16:@145902.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@145901.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@145905.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@145899.4]
  assign regs_14_clock = clock; // @[:@145908.4]
  assign regs_14_reset = io_reset; // @[:@145909.4 RegFile.scala 76:16:@145916.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@145915.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@145919.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@145913.4]
  assign regs_15_clock = clock; // @[:@145922.4]
  assign regs_15_reset = io_reset; // @[:@145923.4 RegFile.scala 76:16:@145930.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@145929.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@145933.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@145927.4]
  assign regs_16_clock = clock; // @[:@145936.4]
  assign regs_16_reset = io_reset; // @[:@145937.4 RegFile.scala 76:16:@145944.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@145943.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@145947.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@145941.4]
  assign regs_17_clock = clock; // @[:@145950.4]
  assign regs_17_reset = io_reset; // @[:@145951.4 RegFile.scala 76:16:@145958.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@145957.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@145961.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@145955.4]
  assign regs_18_clock = clock; // @[:@145964.4]
  assign regs_18_reset = io_reset; // @[:@145965.4 RegFile.scala 76:16:@145972.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@145971.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@145975.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@145969.4]
  assign regs_19_clock = clock; // @[:@145978.4]
  assign regs_19_reset = io_reset; // @[:@145979.4 RegFile.scala 76:16:@145986.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@145985.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@145989.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@145983.4]
  assign regs_20_clock = clock; // @[:@145992.4]
  assign regs_20_reset = io_reset; // @[:@145993.4 RegFile.scala 76:16:@146000.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@145999.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@146003.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@145997.4]
  assign regs_21_clock = clock; // @[:@146006.4]
  assign regs_21_reset = io_reset; // @[:@146007.4 RegFile.scala 76:16:@146014.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@146013.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@146017.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@146011.4]
  assign regs_22_clock = clock; // @[:@146020.4]
  assign regs_22_reset = io_reset; // @[:@146021.4 RegFile.scala 76:16:@146028.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@146027.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@146031.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@146025.4]
  assign regs_23_clock = clock; // @[:@146034.4]
  assign regs_23_reset = io_reset; // @[:@146035.4 RegFile.scala 76:16:@146042.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@146041.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@146045.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@146039.4]
  assign regs_24_clock = clock; // @[:@146048.4]
  assign regs_24_reset = io_reset; // @[:@146049.4 RegFile.scala 76:16:@146056.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@146055.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@146059.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@146053.4]
  assign regs_25_clock = clock; // @[:@146062.4]
  assign regs_25_reset = io_reset; // @[:@146063.4 RegFile.scala 76:16:@146070.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@146069.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@146073.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@146067.4]
  assign regs_26_clock = clock; // @[:@146076.4]
  assign regs_26_reset = io_reset; // @[:@146077.4 RegFile.scala 76:16:@146084.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@146083.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@146087.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@146081.4]
  assign regs_27_clock = clock; // @[:@146090.4]
  assign regs_27_reset = io_reset; // @[:@146091.4 RegFile.scala 76:16:@146098.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@146097.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@146101.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@146095.4]
  assign regs_28_clock = clock; // @[:@146104.4]
  assign regs_28_reset = io_reset; // @[:@146105.4 RegFile.scala 76:16:@146112.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@146111.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@146115.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@146109.4]
  assign regs_29_clock = clock; // @[:@146118.4]
  assign regs_29_reset = io_reset; // @[:@146119.4 RegFile.scala 76:16:@146126.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@146125.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@146129.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@146123.4]
  assign regs_30_clock = clock; // @[:@146132.4]
  assign regs_30_reset = io_reset; // @[:@146133.4 RegFile.scala 76:16:@146140.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@146139.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@146143.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@146137.4]
  assign regs_31_clock = clock; // @[:@146146.4]
  assign regs_31_reset = io_reset; // @[:@146147.4 RegFile.scala 76:16:@146154.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@146153.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@146157.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@146151.4]
  assign regs_32_clock = clock; // @[:@146160.4]
  assign regs_32_reset = io_reset; // @[:@146161.4 RegFile.scala 76:16:@146168.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@146167.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@146171.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@146165.4]
  assign regs_33_clock = clock; // @[:@146174.4]
  assign regs_33_reset = io_reset; // @[:@146175.4 RegFile.scala 76:16:@146182.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@146181.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@146185.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@146179.4]
  assign regs_34_clock = clock; // @[:@146188.4]
  assign regs_34_reset = io_reset; // @[:@146189.4 RegFile.scala 76:16:@146196.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@146195.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@146199.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@146193.4]
  assign regs_35_clock = clock; // @[:@146202.4]
  assign regs_35_reset = io_reset; // @[:@146203.4 RegFile.scala 76:16:@146210.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@146209.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@146213.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@146207.4]
  assign regs_36_clock = clock; // @[:@146216.4]
  assign regs_36_reset = io_reset; // @[:@146217.4 RegFile.scala 76:16:@146224.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@146223.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@146227.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@146221.4]
  assign regs_37_clock = clock; // @[:@146230.4]
  assign regs_37_reset = io_reset; // @[:@146231.4 RegFile.scala 76:16:@146238.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@146237.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@146241.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@146235.4]
  assign regs_38_clock = clock; // @[:@146244.4]
  assign regs_38_reset = io_reset; // @[:@146245.4 RegFile.scala 76:16:@146252.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@146251.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@146255.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@146249.4]
  assign regs_39_clock = clock; // @[:@146258.4]
  assign regs_39_reset = io_reset; // @[:@146259.4 RegFile.scala 76:16:@146266.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@146265.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@146269.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@146263.4]
  assign regs_40_clock = clock; // @[:@146272.4]
  assign regs_40_reset = io_reset; // @[:@146273.4 RegFile.scala 76:16:@146280.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@146279.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@146283.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@146277.4]
  assign regs_41_clock = clock; // @[:@146286.4]
  assign regs_41_reset = io_reset; // @[:@146287.4 RegFile.scala 76:16:@146294.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@146293.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@146297.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@146291.4]
  assign regs_42_clock = clock; // @[:@146300.4]
  assign regs_42_reset = io_reset; // @[:@146301.4 RegFile.scala 76:16:@146308.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@146307.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@146311.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@146305.4]
  assign regs_43_clock = clock; // @[:@146314.4]
  assign regs_43_reset = io_reset; // @[:@146315.4 RegFile.scala 76:16:@146322.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@146321.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@146325.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@146319.4]
  assign regs_44_clock = clock; // @[:@146328.4]
  assign regs_44_reset = io_reset; // @[:@146329.4 RegFile.scala 76:16:@146336.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@146335.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@146339.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@146333.4]
  assign regs_45_clock = clock; // @[:@146342.4]
  assign regs_45_reset = io_reset; // @[:@146343.4 RegFile.scala 76:16:@146350.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@146349.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@146353.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@146347.4]
  assign regs_46_clock = clock; // @[:@146356.4]
  assign regs_46_reset = io_reset; // @[:@146357.4 RegFile.scala 76:16:@146364.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@146363.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@146367.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@146361.4]
  assign regs_47_clock = clock; // @[:@146370.4]
  assign regs_47_reset = io_reset; // @[:@146371.4 RegFile.scala 76:16:@146378.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@146377.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@146381.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@146375.4]
  assign regs_48_clock = clock; // @[:@146384.4]
  assign regs_48_reset = io_reset; // @[:@146385.4 RegFile.scala 76:16:@146392.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@146391.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@146395.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@146389.4]
  assign regs_49_clock = clock; // @[:@146398.4]
  assign regs_49_reset = io_reset; // @[:@146399.4 RegFile.scala 76:16:@146406.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@146405.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@146409.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@146403.4]
  assign regs_50_clock = clock; // @[:@146412.4]
  assign regs_50_reset = io_reset; // @[:@146413.4 RegFile.scala 76:16:@146420.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@146419.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@146423.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@146417.4]
  assign regs_51_clock = clock; // @[:@146426.4]
  assign regs_51_reset = io_reset; // @[:@146427.4 RegFile.scala 76:16:@146434.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@146433.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@146437.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@146431.4]
  assign regs_52_clock = clock; // @[:@146440.4]
  assign regs_52_reset = io_reset; // @[:@146441.4 RegFile.scala 76:16:@146448.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@146447.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@146451.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@146445.4]
  assign regs_53_clock = clock; // @[:@146454.4]
  assign regs_53_reset = io_reset; // @[:@146455.4 RegFile.scala 76:16:@146462.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@146461.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@146465.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@146459.4]
  assign regs_54_clock = clock; // @[:@146468.4]
  assign regs_54_reset = io_reset; // @[:@146469.4 RegFile.scala 76:16:@146476.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@146475.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@146479.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@146473.4]
  assign regs_55_clock = clock; // @[:@146482.4]
  assign regs_55_reset = io_reset; // @[:@146483.4 RegFile.scala 76:16:@146490.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@146489.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@146493.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@146487.4]
  assign regs_56_clock = clock; // @[:@146496.4]
  assign regs_56_reset = io_reset; // @[:@146497.4 RegFile.scala 76:16:@146504.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@146503.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@146507.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@146501.4]
  assign regs_57_clock = clock; // @[:@146510.4]
  assign regs_57_reset = io_reset; // @[:@146511.4 RegFile.scala 76:16:@146518.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@146517.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@146521.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@146515.4]
  assign regs_58_clock = clock; // @[:@146524.4]
  assign regs_58_reset = io_reset; // @[:@146525.4 RegFile.scala 76:16:@146532.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@146531.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@146535.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@146529.4]
  assign regs_59_clock = clock; // @[:@146538.4]
  assign regs_59_reset = io_reset; // @[:@146539.4 RegFile.scala 76:16:@146546.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@146545.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@146549.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@146543.4]
  assign regs_60_clock = clock; // @[:@146552.4]
  assign regs_60_reset = io_reset; // @[:@146553.4 RegFile.scala 76:16:@146560.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@146559.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@146563.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@146557.4]
  assign regs_61_clock = clock; // @[:@146566.4]
  assign regs_61_reset = io_reset; // @[:@146567.4 RegFile.scala 76:16:@146574.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@146573.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@146577.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@146571.4]
  assign regs_62_clock = clock; // @[:@146580.4]
  assign regs_62_reset = io_reset; // @[:@146581.4 RegFile.scala 76:16:@146588.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@146587.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@146591.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@146585.4]
  assign regs_63_clock = clock; // @[:@146594.4]
  assign regs_63_reset = io_reset; // @[:@146595.4 RegFile.scala 76:16:@146602.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@146601.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@146605.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@146599.4]
  assign regs_64_clock = clock; // @[:@146608.4]
  assign regs_64_reset = io_reset; // @[:@146609.4 RegFile.scala 76:16:@146616.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@146615.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@146619.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@146613.4]
  assign regs_65_clock = clock; // @[:@146622.4]
  assign regs_65_reset = io_reset; // @[:@146623.4 RegFile.scala 76:16:@146630.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@146629.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@146633.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@146627.4]
  assign regs_66_clock = clock; // @[:@146636.4]
  assign regs_66_reset = io_reset; // @[:@146637.4 RegFile.scala 76:16:@146644.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@146643.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@146647.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@146641.4]
  assign regs_67_clock = clock; // @[:@146650.4]
  assign regs_67_reset = io_reset; // @[:@146651.4 RegFile.scala 76:16:@146658.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@146657.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@146661.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@146655.4]
  assign regs_68_clock = clock; // @[:@146664.4]
  assign regs_68_reset = io_reset; // @[:@146665.4 RegFile.scala 76:16:@146672.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@146671.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@146675.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@146669.4]
  assign regs_69_clock = clock; // @[:@146678.4]
  assign regs_69_reset = io_reset; // @[:@146679.4 RegFile.scala 76:16:@146686.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@146685.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@146689.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@146683.4]
  assign regs_70_clock = clock; // @[:@146692.4]
  assign regs_70_reset = io_reset; // @[:@146693.4 RegFile.scala 76:16:@146700.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@146699.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@146703.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@146697.4]
  assign regs_71_clock = clock; // @[:@146706.4]
  assign regs_71_reset = io_reset; // @[:@146707.4 RegFile.scala 76:16:@146714.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@146713.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@146717.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@146711.4]
  assign regs_72_clock = clock; // @[:@146720.4]
  assign regs_72_reset = io_reset; // @[:@146721.4 RegFile.scala 76:16:@146728.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@146727.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@146731.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@146725.4]
  assign regs_73_clock = clock; // @[:@146734.4]
  assign regs_73_reset = io_reset; // @[:@146735.4 RegFile.scala 76:16:@146742.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@146741.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@146745.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@146739.4]
  assign regs_74_clock = clock; // @[:@146748.4]
  assign regs_74_reset = io_reset; // @[:@146749.4 RegFile.scala 76:16:@146756.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@146755.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@146759.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@146753.4]
  assign regs_75_clock = clock; // @[:@146762.4]
  assign regs_75_reset = io_reset; // @[:@146763.4 RegFile.scala 76:16:@146770.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@146769.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@146773.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@146767.4]
  assign regs_76_clock = clock; // @[:@146776.4]
  assign regs_76_reset = io_reset; // @[:@146777.4 RegFile.scala 76:16:@146784.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@146783.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@146787.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@146781.4]
  assign regs_77_clock = clock; // @[:@146790.4]
  assign regs_77_reset = io_reset; // @[:@146791.4 RegFile.scala 76:16:@146798.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@146797.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@146801.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@146795.4]
  assign regs_78_clock = clock; // @[:@146804.4]
  assign regs_78_reset = io_reset; // @[:@146805.4 RegFile.scala 76:16:@146812.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@146811.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@146815.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@146809.4]
  assign regs_79_clock = clock; // @[:@146818.4]
  assign regs_79_reset = io_reset; // @[:@146819.4 RegFile.scala 76:16:@146826.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@146825.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@146829.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@146823.4]
  assign regs_80_clock = clock; // @[:@146832.4]
  assign regs_80_reset = io_reset; // @[:@146833.4 RegFile.scala 76:16:@146840.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@146839.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@146843.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@146837.4]
  assign regs_81_clock = clock; // @[:@146846.4]
  assign regs_81_reset = io_reset; // @[:@146847.4 RegFile.scala 76:16:@146854.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@146853.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@146857.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@146851.4]
  assign regs_82_clock = clock; // @[:@146860.4]
  assign regs_82_reset = io_reset; // @[:@146861.4 RegFile.scala 76:16:@146868.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@146867.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@146871.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@146865.4]
  assign regs_83_clock = clock; // @[:@146874.4]
  assign regs_83_reset = io_reset; // @[:@146875.4 RegFile.scala 76:16:@146882.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@146881.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@146885.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@146879.4]
  assign regs_84_clock = clock; // @[:@146888.4]
  assign regs_84_reset = io_reset; // @[:@146889.4 RegFile.scala 76:16:@146896.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@146895.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@146899.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@146893.4]
  assign regs_85_clock = clock; // @[:@146902.4]
  assign regs_85_reset = io_reset; // @[:@146903.4 RegFile.scala 76:16:@146910.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@146909.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@146913.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@146907.4]
  assign regs_86_clock = clock; // @[:@146916.4]
  assign regs_86_reset = io_reset; // @[:@146917.4 RegFile.scala 76:16:@146924.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@146923.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@146927.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@146921.4]
  assign regs_87_clock = clock; // @[:@146930.4]
  assign regs_87_reset = io_reset; // @[:@146931.4 RegFile.scala 76:16:@146938.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@146937.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@146941.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@146935.4]
  assign regs_88_clock = clock; // @[:@146944.4]
  assign regs_88_reset = io_reset; // @[:@146945.4 RegFile.scala 76:16:@146952.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@146951.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@146955.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@146949.4]
  assign regs_89_clock = clock; // @[:@146958.4]
  assign regs_89_reset = io_reset; // @[:@146959.4 RegFile.scala 76:16:@146966.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@146965.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@146969.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@146963.4]
  assign regs_90_clock = clock; // @[:@146972.4]
  assign regs_90_reset = io_reset; // @[:@146973.4 RegFile.scala 76:16:@146980.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@146979.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@146983.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@146977.4]
  assign regs_91_clock = clock; // @[:@146986.4]
  assign regs_91_reset = io_reset; // @[:@146987.4 RegFile.scala 76:16:@146994.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@146993.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@146997.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@146991.4]
  assign regs_92_clock = clock; // @[:@147000.4]
  assign regs_92_reset = io_reset; // @[:@147001.4 RegFile.scala 76:16:@147008.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@147007.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@147011.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@147005.4]
  assign regs_93_clock = clock; // @[:@147014.4]
  assign regs_93_reset = io_reset; // @[:@147015.4 RegFile.scala 76:16:@147022.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@147021.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@147025.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@147019.4]
  assign regs_94_clock = clock; // @[:@147028.4]
  assign regs_94_reset = io_reset; // @[:@147029.4 RegFile.scala 76:16:@147036.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@147035.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@147039.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@147033.4]
  assign regs_95_clock = clock; // @[:@147042.4]
  assign regs_95_reset = io_reset; // @[:@147043.4 RegFile.scala 76:16:@147050.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@147049.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@147053.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@147047.4]
  assign regs_96_clock = clock; // @[:@147056.4]
  assign regs_96_reset = io_reset; // @[:@147057.4 RegFile.scala 76:16:@147064.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@147063.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@147067.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@147061.4]
  assign regs_97_clock = clock; // @[:@147070.4]
  assign regs_97_reset = io_reset; // @[:@147071.4 RegFile.scala 76:16:@147078.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@147077.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@147081.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@147075.4]
  assign regs_98_clock = clock; // @[:@147084.4]
  assign regs_98_reset = io_reset; // @[:@147085.4 RegFile.scala 76:16:@147092.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@147091.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@147095.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@147089.4]
  assign regs_99_clock = clock; // @[:@147098.4]
  assign regs_99_reset = io_reset; // @[:@147099.4 RegFile.scala 76:16:@147106.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@147105.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@147109.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@147103.4]
  assign regs_100_clock = clock; // @[:@147112.4]
  assign regs_100_reset = io_reset; // @[:@147113.4 RegFile.scala 76:16:@147120.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@147119.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@147123.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@147117.4]
  assign regs_101_clock = clock; // @[:@147126.4]
  assign regs_101_reset = io_reset; // @[:@147127.4 RegFile.scala 76:16:@147134.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@147133.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@147137.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@147131.4]
  assign regs_102_clock = clock; // @[:@147140.4]
  assign regs_102_reset = io_reset; // @[:@147141.4 RegFile.scala 76:16:@147148.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@147147.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@147151.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@147145.4]
  assign regs_103_clock = clock; // @[:@147154.4]
  assign regs_103_reset = io_reset; // @[:@147155.4 RegFile.scala 76:16:@147162.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@147161.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@147165.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@147159.4]
  assign regs_104_clock = clock; // @[:@147168.4]
  assign regs_104_reset = io_reset; // @[:@147169.4 RegFile.scala 76:16:@147176.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@147175.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@147179.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@147173.4]
  assign regs_105_clock = clock; // @[:@147182.4]
  assign regs_105_reset = io_reset; // @[:@147183.4 RegFile.scala 76:16:@147190.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@147189.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@147193.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@147187.4]
  assign regs_106_clock = clock; // @[:@147196.4]
  assign regs_106_reset = io_reset; // @[:@147197.4 RegFile.scala 76:16:@147204.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@147203.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@147207.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@147201.4]
  assign regs_107_clock = clock; // @[:@147210.4]
  assign regs_107_reset = io_reset; // @[:@147211.4 RegFile.scala 76:16:@147218.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@147217.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@147221.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@147215.4]
  assign regs_108_clock = clock; // @[:@147224.4]
  assign regs_108_reset = io_reset; // @[:@147225.4 RegFile.scala 76:16:@147232.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@147231.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@147235.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@147229.4]
  assign regs_109_clock = clock; // @[:@147238.4]
  assign regs_109_reset = io_reset; // @[:@147239.4 RegFile.scala 76:16:@147246.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@147245.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@147249.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@147243.4]
  assign regs_110_clock = clock; // @[:@147252.4]
  assign regs_110_reset = io_reset; // @[:@147253.4 RegFile.scala 76:16:@147260.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@147259.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@147263.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@147257.4]
  assign regs_111_clock = clock; // @[:@147266.4]
  assign regs_111_reset = io_reset; // @[:@147267.4 RegFile.scala 76:16:@147274.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@147273.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@147277.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@147271.4]
  assign regs_112_clock = clock; // @[:@147280.4]
  assign regs_112_reset = io_reset; // @[:@147281.4 RegFile.scala 76:16:@147288.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@147287.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@147291.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@147285.4]
  assign regs_113_clock = clock; // @[:@147294.4]
  assign regs_113_reset = io_reset; // @[:@147295.4 RegFile.scala 76:16:@147302.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@147301.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@147305.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@147299.4]
  assign regs_114_clock = clock; // @[:@147308.4]
  assign regs_114_reset = io_reset; // @[:@147309.4 RegFile.scala 76:16:@147316.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@147315.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@147319.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@147313.4]
  assign regs_115_clock = clock; // @[:@147322.4]
  assign regs_115_reset = io_reset; // @[:@147323.4 RegFile.scala 76:16:@147330.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@147329.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@147333.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@147327.4]
  assign regs_116_clock = clock; // @[:@147336.4]
  assign regs_116_reset = io_reset; // @[:@147337.4 RegFile.scala 76:16:@147344.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@147343.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@147347.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@147341.4]
  assign regs_117_clock = clock; // @[:@147350.4]
  assign regs_117_reset = io_reset; // @[:@147351.4 RegFile.scala 76:16:@147358.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@147357.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@147361.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@147355.4]
  assign regs_118_clock = clock; // @[:@147364.4]
  assign regs_118_reset = io_reset; // @[:@147365.4 RegFile.scala 76:16:@147372.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@147371.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@147375.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@147369.4]
  assign regs_119_clock = clock; // @[:@147378.4]
  assign regs_119_reset = io_reset; // @[:@147379.4 RegFile.scala 76:16:@147386.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@147385.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@147389.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@147383.4]
  assign regs_120_clock = clock; // @[:@147392.4]
  assign regs_120_reset = io_reset; // @[:@147393.4 RegFile.scala 76:16:@147400.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@147399.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@147403.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@147397.4]
  assign regs_121_clock = clock; // @[:@147406.4]
  assign regs_121_reset = io_reset; // @[:@147407.4 RegFile.scala 76:16:@147414.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@147413.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@147417.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@147411.4]
  assign regs_122_clock = clock; // @[:@147420.4]
  assign regs_122_reset = io_reset; // @[:@147421.4 RegFile.scala 76:16:@147428.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@147427.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@147431.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@147425.4]
  assign regs_123_clock = clock; // @[:@147434.4]
  assign regs_123_reset = io_reset; // @[:@147435.4 RegFile.scala 76:16:@147442.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@147441.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@147445.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@147439.4]
  assign regs_124_clock = clock; // @[:@147448.4]
  assign regs_124_reset = io_reset; // @[:@147449.4 RegFile.scala 76:16:@147456.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@147455.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@147459.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@147453.4]
  assign regs_125_clock = clock; // @[:@147462.4]
  assign regs_125_reset = io_reset; // @[:@147463.4 RegFile.scala 76:16:@147470.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@147469.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@147473.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@147467.4]
  assign regs_126_clock = clock; // @[:@147476.4]
  assign regs_126_reset = io_reset; // @[:@147477.4 RegFile.scala 76:16:@147484.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@147483.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@147487.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@147481.4]
  assign regs_127_clock = clock; // @[:@147490.4]
  assign regs_127_reset = io_reset; // @[:@147491.4 RegFile.scala 76:16:@147498.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@147497.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@147501.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@147495.4]
  assign regs_128_clock = clock; // @[:@147504.4]
  assign regs_128_reset = io_reset; // @[:@147505.4 RegFile.scala 76:16:@147512.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@147511.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@147515.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@147509.4]
  assign regs_129_clock = clock; // @[:@147518.4]
  assign regs_129_reset = io_reset; // @[:@147519.4 RegFile.scala 76:16:@147526.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@147525.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@147529.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@147523.4]
  assign regs_130_clock = clock; // @[:@147532.4]
  assign regs_130_reset = io_reset; // @[:@147533.4 RegFile.scala 76:16:@147540.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@147539.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@147543.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@147537.4]
  assign regs_131_clock = clock; // @[:@147546.4]
  assign regs_131_reset = io_reset; // @[:@147547.4 RegFile.scala 76:16:@147554.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@147553.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@147557.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@147551.4]
  assign regs_132_clock = clock; // @[:@147560.4]
  assign regs_132_reset = io_reset; // @[:@147561.4 RegFile.scala 76:16:@147568.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@147567.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@147571.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@147565.4]
  assign regs_133_clock = clock; // @[:@147574.4]
  assign regs_133_reset = io_reset; // @[:@147575.4 RegFile.scala 76:16:@147582.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@147581.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@147585.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@147579.4]
  assign regs_134_clock = clock; // @[:@147588.4]
  assign regs_134_reset = io_reset; // @[:@147589.4 RegFile.scala 76:16:@147596.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@147595.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@147599.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@147593.4]
  assign regs_135_clock = clock; // @[:@147602.4]
  assign regs_135_reset = io_reset; // @[:@147603.4 RegFile.scala 76:16:@147610.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@147609.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@147613.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@147607.4]
  assign regs_136_clock = clock; // @[:@147616.4]
  assign regs_136_reset = io_reset; // @[:@147617.4 RegFile.scala 76:16:@147624.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@147623.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@147627.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@147621.4]
  assign regs_137_clock = clock; // @[:@147630.4]
  assign regs_137_reset = io_reset; // @[:@147631.4 RegFile.scala 76:16:@147638.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@147637.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@147641.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@147635.4]
  assign regs_138_clock = clock; // @[:@147644.4]
  assign regs_138_reset = io_reset; // @[:@147645.4 RegFile.scala 76:16:@147652.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@147651.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@147655.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@147649.4]
  assign regs_139_clock = clock; // @[:@147658.4]
  assign regs_139_reset = io_reset; // @[:@147659.4 RegFile.scala 76:16:@147666.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@147665.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@147669.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@147663.4]
  assign regs_140_clock = clock; // @[:@147672.4]
  assign regs_140_reset = io_reset; // @[:@147673.4 RegFile.scala 76:16:@147680.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@147679.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@147683.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@147677.4]
  assign regs_141_clock = clock; // @[:@147686.4]
  assign regs_141_reset = io_reset; // @[:@147687.4 RegFile.scala 76:16:@147694.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@147693.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@147697.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@147691.4]
  assign regs_142_clock = clock; // @[:@147700.4]
  assign regs_142_reset = io_reset; // @[:@147701.4 RegFile.scala 76:16:@147708.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@147707.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@147711.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@147705.4]
  assign regs_143_clock = clock; // @[:@147714.4]
  assign regs_143_reset = io_reset; // @[:@147715.4 RegFile.scala 76:16:@147722.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@147721.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@147725.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@147719.4]
  assign regs_144_clock = clock; // @[:@147728.4]
  assign regs_144_reset = io_reset; // @[:@147729.4 RegFile.scala 76:16:@147736.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@147735.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@147739.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@147733.4]
  assign regs_145_clock = clock; // @[:@147742.4]
  assign regs_145_reset = io_reset; // @[:@147743.4 RegFile.scala 76:16:@147750.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@147749.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@147753.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@147747.4]
  assign regs_146_clock = clock; // @[:@147756.4]
  assign regs_146_reset = io_reset; // @[:@147757.4 RegFile.scala 76:16:@147764.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@147763.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@147767.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@147761.4]
  assign regs_147_clock = clock; // @[:@147770.4]
  assign regs_147_reset = io_reset; // @[:@147771.4 RegFile.scala 76:16:@147778.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@147777.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@147781.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@147775.4]
  assign regs_148_clock = clock; // @[:@147784.4]
  assign regs_148_reset = io_reset; // @[:@147785.4 RegFile.scala 76:16:@147792.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@147791.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@147795.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@147789.4]
  assign regs_149_clock = clock; // @[:@147798.4]
  assign regs_149_reset = io_reset; // @[:@147799.4 RegFile.scala 76:16:@147806.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@147805.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@147809.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@147803.4]
  assign regs_150_clock = clock; // @[:@147812.4]
  assign regs_150_reset = io_reset; // @[:@147813.4 RegFile.scala 76:16:@147820.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@147819.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@147823.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@147817.4]
  assign regs_151_clock = clock; // @[:@147826.4]
  assign regs_151_reset = io_reset; // @[:@147827.4 RegFile.scala 76:16:@147834.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@147833.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@147837.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@147831.4]
  assign regs_152_clock = clock; // @[:@147840.4]
  assign regs_152_reset = io_reset; // @[:@147841.4 RegFile.scala 76:16:@147848.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@147847.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@147851.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@147845.4]
  assign regs_153_clock = clock; // @[:@147854.4]
  assign regs_153_reset = io_reset; // @[:@147855.4 RegFile.scala 76:16:@147862.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@147861.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@147865.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@147859.4]
  assign regs_154_clock = clock; // @[:@147868.4]
  assign regs_154_reset = io_reset; // @[:@147869.4 RegFile.scala 76:16:@147876.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@147875.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@147879.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@147873.4]
  assign regs_155_clock = clock; // @[:@147882.4]
  assign regs_155_reset = io_reset; // @[:@147883.4 RegFile.scala 76:16:@147890.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@147889.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@147893.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@147887.4]
  assign regs_156_clock = clock; // @[:@147896.4]
  assign regs_156_reset = io_reset; // @[:@147897.4 RegFile.scala 76:16:@147904.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@147903.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@147907.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@147901.4]
  assign regs_157_clock = clock; // @[:@147910.4]
  assign regs_157_reset = io_reset; // @[:@147911.4 RegFile.scala 76:16:@147918.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@147917.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@147921.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@147915.4]
  assign regs_158_clock = clock; // @[:@147924.4]
  assign regs_158_reset = io_reset; // @[:@147925.4 RegFile.scala 76:16:@147932.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@147931.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@147935.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@147929.4]
  assign regs_159_clock = clock; // @[:@147938.4]
  assign regs_159_reset = io_reset; // @[:@147939.4 RegFile.scala 76:16:@147946.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@147945.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@147949.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@147943.4]
  assign regs_160_clock = clock; // @[:@147952.4]
  assign regs_160_reset = io_reset; // @[:@147953.4 RegFile.scala 76:16:@147960.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@147959.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@147963.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@147957.4]
  assign regs_161_clock = clock; // @[:@147966.4]
  assign regs_161_reset = io_reset; // @[:@147967.4 RegFile.scala 76:16:@147974.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@147973.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@147977.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@147971.4]
  assign regs_162_clock = clock; // @[:@147980.4]
  assign regs_162_reset = io_reset; // @[:@147981.4 RegFile.scala 76:16:@147988.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@147987.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@147991.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@147985.4]
  assign regs_163_clock = clock; // @[:@147994.4]
  assign regs_163_reset = io_reset; // @[:@147995.4 RegFile.scala 76:16:@148002.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@148001.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@148005.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@147999.4]
  assign regs_164_clock = clock; // @[:@148008.4]
  assign regs_164_reset = io_reset; // @[:@148009.4 RegFile.scala 76:16:@148016.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@148015.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@148019.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@148013.4]
  assign regs_165_clock = clock; // @[:@148022.4]
  assign regs_165_reset = io_reset; // @[:@148023.4 RegFile.scala 76:16:@148030.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@148029.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@148033.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@148027.4]
  assign regs_166_clock = clock; // @[:@148036.4]
  assign regs_166_reset = io_reset; // @[:@148037.4 RegFile.scala 76:16:@148044.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@148043.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@148047.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@148041.4]
  assign regs_167_clock = clock; // @[:@148050.4]
  assign regs_167_reset = io_reset; // @[:@148051.4 RegFile.scala 76:16:@148058.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@148057.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@148061.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@148055.4]
  assign regs_168_clock = clock; // @[:@148064.4]
  assign regs_168_reset = io_reset; // @[:@148065.4 RegFile.scala 76:16:@148072.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@148071.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@148075.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@148069.4]
  assign regs_169_clock = clock; // @[:@148078.4]
  assign regs_169_reset = io_reset; // @[:@148079.4 RegFile.scala 76:16:@148086.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@148085.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@148089.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@148083.4]
  assign regs_170_clock = clock; // @[:@148092.4]
  assign regs_170_reset = io_reset; // @[:@148093.4 RegFile.scala 76:16:@148100.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@148099.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@148103.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@148097.4]
  assign regs_171_clock = clock; // @[:@148106.4]
  assign regs_171_reset = io_reset; // @[:@148107.4 RegFile.scala 76:16:@148114.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@148113.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@148117.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@148111.4]
  assign regs_172_clock = clock; // @[:@148120.4]
  assign regs_172_reset = io_reset; // @[:@148121.4 RegFile.scala 76:16:@148128.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@148127.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@148131.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@148125.4]
  assign regs_173_clock = clock; // @[:@148134.4]
  assign regs_173_reset = io_reset; // @[:@148135.4 RegFile.scala 76:16:@148142.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@148141.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@148145.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@148139.4]
  assign regs_174_clock = clock; // @[:@148148.4]
  assign regs_174_reset = io_reset; // @[:@148149.4 RegFile.scala 76:16:@148156.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@148155.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@148159.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@148153.4]
  assign regs_175_clock = clock; // @[:@148162.4]
  assign regs_175_reset = io_reset; // @[:@148163.4 RegFile.scala 76:16:@148170.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@148169.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@148173.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@148167.4]
  assign regs_176_clock = clock; // @[:@148176.4]
  assign regs_176_reset = io_reset; // @[:@148177.4 RegFile.scala 76:16:@148184.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@148183.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@148187.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@148181.4]
  assign regs_177_clock = clock; // @[:@148190.4]
  assign regs_177_reset = io_reset; // @[:@148191.4 RegFile.scala 76:16:@148198.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@148197.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@148201.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@148195.4]
  assign regs_178_clock = clock; // @[:@148204.4]
  assign regs_178_reset = io_reset; // @[:@148205.4 RegFile.scala 76:16:@148212.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@148211.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@148215.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@148209.4]
  assign regs_179_clock = clock; // @[:@148218.4]
  assign regs_179_reset = io_reset; // @[:@148219.4 RegFile.scala 76:16:@148226.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@148225.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@148229.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@148223.4]
  assign regs_180_clock = clock; // @[:@148232.4]
  assign regs_180_reset = io_reset; // @[:@148233.4 RegFile.scala 76:16:@148240.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@148239.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@148243.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@148237.4]
  assign regs_181_clock = clock; // @[:@148246.4]
  assign regs_181_reset = io_reset; // @[:@148247.4 RegFile.scala 76:16:@148254.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@148253.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@148257.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@148251.4]
  assign regs_182_clock = clock; // @[:@148260.4]
  assign regs_182_reset = io_reset; // @[:@148261.4 RegFile.scala 76:16:@148268.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@148267.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@148271.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@148265.4]
  assign regs_183_clock = clock; // @[:@148274.4]
  assign regs_183_reset = io_reset; // @[:@148275.4 RegFile.scala 76:16:@148282.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@148281.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@148285.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@148279.4]
  assign regs_184_clock = clock; // @[:@148288.4]
  assign regs_184_reset = io_reset; // @[:@148289.4 RegFile.scala 76:16:@148296.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@148295.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@148299.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@148293.4]
  assign regs_185_clock = clock; // @[:@148302.4]
  assign regs_185_reset = io_reset; // @[:@148303.4 RegFile.scala 76:16:@148310.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@148309.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@148313.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@148307.4]
  assign regs_186_clock = clock; // @[:@148316.4]
  assign regs_186_reset = io_reset; // @[:@148317.4 RegFile.scala 76:16:@148324.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@148323.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@148327.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@148321.4]
  assign regs_187_clock = clock; // @[:@148330.4]
  assign regs_187_reset = io_reset; // @[:@148331.4 RegFile.scala 76:16:@148338.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@148337.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@148341.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@148335.4]
  assign regs_188_clock = clock; // @[:@148344.4]
  assign regs_188_reset = io_reset; // @[:@148345.4 RegFile.scala 76:16:@148352.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@148351.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@148355.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@148349.4]
  assign regs_189_clock = clock; // @[:@148358.4]
  assign regs_189_reset = io_reset; // @[:@148359.4 RegFile.scala 76:16:@148366.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@148365.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@148369.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@148363.4]
  assign regs_190_clock = clock; // @[:@148372.4]
  assign regs_190_reset = io_reset; // @[:@148373.4 RegFile.scala 76:16:@148380.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@148379.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@148383.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@148377.4]
  assign regs_191_clock = clock; // @[:@148386.4]
  assign regs_191_reset = io_reset; // @[:@148387.4 RegFile.scala 76:16:@148394.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@148393.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@148397.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@148391.4]
  assign regs_192_clock = clock; // @[:@148400.4]
  assign regs_192_reset = io_reset; // @[:@148401.4 RegFile.scala 76:16:@148408.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@148407.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@148411.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@148405.4]
  assign regs_193_clock = clock; // @[:@148414.4]
  assign regs_193_reset = io_reset; // @[:@148415.4 RegFile.scala 76:16:@148422.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@148421.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@148425.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@148419.4]
  assign regs_194_clock = clock; // @[:@148428.4]
  assign regs_194_reset = io_reset; // @[:@148429.4 RegFile.scala 76:16:@148436.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@148435.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@148439.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@148433.4]
  assign regs_195_clock = clock; // @[:@148442.4]
  assign regs_195_reset = io_reset; // @[:@148443.4 RegFile.scala 76:16:@148450.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@148449.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@148453.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@148447.4]
  assign regs_196_clock = clock; // @[:@148456.4]
  assign regs_196_reset = io_reset; // @[:@148457.4 RegFile.scala 76:16:@148464.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@148463.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@148467.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@148461.4]
  assign regs_197_clock = clock; // @[:@148470.4]
  assign regs_197_reset = io_reset; // @[:@148471.4 RegFile.scala 76:16:@148478.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@148477.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@148481.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@148475.4]
  assign regs_198_clock = clock; // @[:@148484.4]
  assign regs_198_reset = io_reset; // @[:@148485.4 RegFile.scala 76:16:@148492.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@148491.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@148495.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@148489.4]
  assign regs_199_clock = clock; // @[:@148498.4]
  assign regs_199_reset = io_reset; // @[:@148499.4 RegFile.scala 76:16:@148506.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@148505.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@148509.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@148503.4]
  assign regs_200_clock = clock; // @[:@148512.4]
  assign regs_200_reset = io_reset; // @[:@148513.4 RegFile.scala 76:16:@148520.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@148519.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@148523.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@148517.4]
  assign regs_201_clock = clock; // @[:@148526.4]
  assign regs_201_reset = io_reset; // @[:@148527.4 RegFile.scala 76:16:@148534.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@148533.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@148537.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@148531.4]
  assign regs_202_clock = clock; // @[:@148540.4]
  assign regs_202_reset = io_reset; // @[:@148541.4 RegFile.scala 76:16:@148548.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@148547.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@148551.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@148545.4]
  assign regs_203_clock = clock; // @[:@148554.4]
  assign regs_203_reset = io_reset; // @[:@148555.4 RegFile.scala 76:16:@148562.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@148561.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@148565.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@148559.4]
  assign regs_204_clock = clock; // @[:@148568.4]
  assign regs_204_reset = io_reset; // @[:@148569.4 RegFile.scala 76:16:@148576.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@148575.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@148579.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@148573.4]
  assign regs_205_clock = clock; // @[:@148582.4]
  assign regs_205_reset = io_reset; // @[:@148583.4 RegFile.scala 76:16:@148590.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@148589.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@148593.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@148587.4]
  assign regs_206_clock = clock; // @[:@148596.4]
  assign regs_206_reset = io_reset; // @[:@148597.4 RegFile.scala 76:16:@148604.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@148603.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@148607.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@148601.4]
  assign regs_207_clock = clock; // @[:@148610.4]
  assign regs_207_reset = io_reset; // @[:@148611.4 RegFile.scala 76:16:@148618.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@148617.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@148621.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@148615.4]
  assign regs_208_clock = clock; // @[:@148624.4]
  assign regs_208_reset = io_reset; // @[:@148625.4 RegFile.scala 76:16:@148632.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@148631.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@148635.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@148629.4]
  assign regs_209_clock = clock; // @[:@148638.4]
  assign regs_209_reset = io_reset; // @[:@148639.4 RegFile.scala 76:16:@148646.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@148645.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@148649.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@148643.4]
  assign regs_210_clock = clock; // @[:@148652.4]
  assign regs_210_reset = io_reset; // @[:@148653.4 RegFile.scala 76:16:@148660.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@148659.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@148663.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@148657.4]
  assign regs_211_clock = clock; // @[:@148666.4]
  assign regs_211_reset = io_reset; // @[:@148667.4 RegFile.scala 76:16:@148674.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@148673.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@148677.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@148671.4]
  assign regs_212_clock = clock; // @[:@148680.4]
  assign regs_212_reset = io_reset; // @[:@148681.4 RegFile.scala 76:16:@148688.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@148687.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@148691.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@148685.4]
  assign regs_213_clock = clock; // @[:@148694.4]
  assign regs_213_reset = io_reset; // @[:@148695.4 RegFile.scala 76:16:@148702.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@148701.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@148705.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@148699.4]
  assign regs_214_clock = clock; // @[:@148708.4]
  assign regs_214_reset = io_reset; // @[:@148709.4 RegFile.scala 76:16:@148716.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@148715.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@148719.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@148713.4]
  assign regs_215_clock = clock; // @[:@148722.4]
  assign regs_215_reset = io_reset; // @[:@148723.4 RegFile.scala 76:16:@148730.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@148729.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@148733.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@148727.4]
  assign regs_216_clock = clock; // @[:@148736.4]
  assign regs_216_reset = io_reset; // @[:@148737.4 RegFile.scala 76:16:@148744.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@148743.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@148747.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@148741.4]
  assign regs_217_clock = clock; // @[:@148750.4]
  assign regs_217_reset = io_reset; // @[:@148751.4 RegFile.scala 76:16:@148758.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@148757.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@148761.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@148755.4]
  assign regs_218_clock = clock; // @[:@148764.4]
  assign regs_218_reset = io_reset; // @[:@148765.4 RegFile.scala 76:16:@148772.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@148771.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@148775.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@148769.4]
  assign regs_219_clock = clock; // @[:@148778.4]
  assign regs_219_reset = io_reset; // @[:@148779.4 RegFile.scala 76:16:@148786.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@148785.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@148789.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@148783.4]
  assign regs_220_clock = clock; // @[:@148792.4]
  assign regs_220_reset = io_reset; // @[:@148793.4 RegFile.scala 76:16:@148800.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@148799.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@148803.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@148797.4]
  assign regs_221_clock = clock; // @[:@148806.4]
  assign regs_221_reset = io_reset; // @[:@148807.4 RegFile.scala 76:16:@148814.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@148813.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@148817.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@148811.4]
  assign regs_222_clock = clock; // @[:@148820.4]
  assign regs_222_reset = io_reset; // @[:@148821.4 RegFile.scala 76:16:@148828.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@148827.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@148831.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@148825.4]
  assign regs_223_clock = clock; // @[:@148834.4]
  assign regs_223_reset = io_reset; // @[:@148835.4 RegFile.scala 76:16:@148842.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@148841.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@148845.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@148839.4]
  assign regs_224_clock = clock; // @[:@148848.4]
  assign regs_224_reset = io_reset; // @[:@148849.4 RegFile.scala 76:16:@148856.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@148855.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@148859.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@148853.4]
  assign regs_225_clock = clock; // @[:@148862.4]
  assign regs_225_reset = io_reset; // @[:@148863.4 RegFile.scala 76:16:@148870.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@148869.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@148873.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@148867.4]
  assign regs_226_clock = clock; // @[:@148876.4]
  assign regs_226_reset = io_reset; // @[:@148877.4 RegFile.scala 76:16:@148884.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@148883.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@148887.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@148881.4]
  assign regs_227_clock = clock; // @[:@148890.4]
  assign regs_227_reset = io_reset; // @[:@148891.4 RegFile.scala 76:16:@148898.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@148897.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@148901.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@148895.4]
  assign regs_228_clock = clock; // @[:@148904.4]
  assign regs_228_reset = io_reset; // @[:@148905.4 RegFile.scala 76:16:@148912.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@148911.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@148915.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@148909.4]
  assign regs_229_clock = clock; // @[:@148918.4]
  assign regs_229_reset = io_reset; // @[:@148919.4 RegFile.scala 76:16:@148926.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@148925.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@148929.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@148923.4]
  assign regs_230_clock = clock; // @[:@148932.4]
  assign regs_230_reset = io_reset; // @[:@148933.4 RegFile.scala 76:16:@148940.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@148939.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@148943.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@148937.4]
  assign regs_231_clock = clock; // @[:@148946.4]
  assign regs_231_reset = io_reset; // @[:@148947.4 RegFile.scala 76:16:@148954.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@148953.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@148957.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@148951.4]
  assign regs_232_clock = clock; // @[:@148960.4]
  assign regs_232_reset = io_reset; // @[:@148961.4 RegFile.scala 76:16:@148968.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@148967.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@148971.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@148965.4]
  assign regs_233_clock = clock; // @[:@148974.4]
  assign regs_233_reset = io_reset; // @[:@148975.4 RegFile.scala 76:16:@148982.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@148981.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@148985.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@148979.4]
  assign regs_234_clock = clock; // @[:@148988.4]
  assign regs_234_reset = io_reset; // @[:@148989.4 RegFile.scala 76:16:@148996.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@148995.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@148999.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@148993.4]
  assign regs_235_clock = clock; // @[:@149002.4]
  assign regs_235_reset = io_reset; // @[:@149003.4 RegFile.scala 76:16:@149010.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@149009.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@149013.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@149007.4]
  assign regs_236_clock = clock; // @[:@149016.4]
  assign regs_236_reset = io_reset; // @[:@149017.4 RegFile.scala 76:16:@149024.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@149023.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@149027.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@149021.4]
  assign regs_237_clock = clock; // @[:@149030.4]
  assign regs_237_reset = io_reset; // @[:@149031.4 RegFile.scala 76:16:@149038.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@149037.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@149041.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@149035.4]
  assign regs_238_clock = clock; // @[:@149044.4]
  assign regs_238_reset = io_reset; // @[:@149045.4 RegFile.scala 76:16:@149052.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@149051.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@149055.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@149049.4]
  assign regs_239_clock = clock; // @[:@149058.4]
  assign regs_239_reset = io_reset; // @[:@149059.4 RegFile.scala 76:16:@149066.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@149065.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@149069.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@149063.4]
  assign regs_240_clock = clock; // @[:@149072.4]
  assign regs_240_reset = io_reset; // @[:@149073.4 RegFile.scala 76:16:@149080.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@149079.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@149083.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@149077.4]
  assign regs_241_clock = clock; // @[:@149086.4]
  assign regs_241_reset = io_reset; // @[:@149087.4 RegFile.scala 76:16:@149094.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@149093.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@149097.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@149091.4]
  assign regs_242_clock = clock; // @[:@149100.4]
  assign regs_242_reset = io_reset; // @[:@149101.4 RegFile.scala 76:16:@149108.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@149107.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@149111.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@149105.4]
  assign regs_243_clock = clock; // @[:@149114.4]
  assign regs_243_reset = io_reset; // @[:@149115.4 RegFile.scala 76:16:@149122.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@149121.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@149125.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@149119.4]
  assign regs_244_clock = clock; // @[:@149128.4]
  assign regs_244_reset = io_reset; // @[:@149129.4 RegFile.scala 76:16:@149136.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@149135.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@149139.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@149133.4]
  assign regs_245_clock = clock; // @[:@149142.4]
  assign regs_245_reset = io_reset; // @[:@149143.4 RegFile.scala 76:16:@149150.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@149149.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@149153.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@149147.4]
  assign regs_246_clock = clock; // @[:@149156.4]
  assign regs_246_reset = io_reset; // @[:@149157.4 RegFile.scala 76:16:@149164.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@149163.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@149167.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@149161.4]
  assign regs_247_clock = clock; // @[:@149170.4]
  assign regs_247_reset = io_reset; // @[:@149171.4 RegFile.scala 76:16:@149178.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@149177.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@149181.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@149175.4]
  assign regs_248_clock = clock; // @[:@149184.4]
  assign regs_248_reset = io_reset; // @[:@149185.4 RegFile.scala 76:16:@149192.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@149191.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@149195.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@149189.4]
  assign regs_249_clock = clock; // @[:@149198.4]
  assign regs_249_reset = io_reset; // @[:@149199.4 RegFile.scala 76:16:@149206.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@149205.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@149209.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@149203.4]
  assign regs_250_clock = clock; // @[:@149212.4]
  assign regs_250_reset = io_reset; // @[:@149213.4 RegFile.scala 76:16:@149220.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@149219.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@149223.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@149217.4]
  assign regs_251_clock = clock; // @[:@149226.4]
  assign regs_251_reset = io_reset; // @[:@149227.4 RegFile.scala 76:16:@149234.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@149233.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@149237.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@149231.4]
  assign regs_252_clock = clock; // @[:@149240.4]
  assign regs_252_reset = io_reset; // @[:@149241.4 RegFile.scala 76:16:@149248.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@149247.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@149251.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@149245.4]
  assign regs_253_clock = clock; // @[:@149254.4]
  assign regs_253_reset = io_reset; // @[:@149255.4 RegFile.scala 76:16:@149262.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@149261.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@149265.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@149259.4]
  assign regs_254_clock = clock; // @[:@149268.4]
  assign regs_254_reset = io_reset; // @[:@149269.4 RegFile.scala 76:16:@149276.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@149275.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@149279.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@149273.4]
  assign regs_255_clock = clock; // @[:@149282.4]
  assign regs_255_reset = io_reset; // @[:@149283.4 RegFile.scala 76:16:@149290.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@149289.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@149293.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@149287.4]
  assign regs_256_clock = clock; // @[:@149296.4]
  assign regs_256_reset = io_reset; // @[:@149297.4 RegFile.scala 76:16:@149304.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@149303.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@149307.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@149301.4]
  assign regs_257_clock = clock; // @[:@149310.4]
  assign regs_257_reset = io_reset; // @[:@149311.4 RegFile.scala 76:16:@149318.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@149317.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@149321.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@149315.4]
  assign regs_258_clock = clock; // @[:@149324.4]
  assign regs_258_reset = io_reset; // @[:@149325.4 RegFile.scala 76:16:@149332.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@149331.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@149335.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@149329.4]
  assign regs_259_clock = clock; // @[:@149338.4]
  assign regs_259_reset = io_reset; // @[:@149339.4 RegFile.scala 76:16:@149346.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@149345.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@149349.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@149343.4]
  assign regs_260_clock = clock; // @[:@149352.4]
  assign regs_260_reset = io_reset; // @[:@149353.4 RegFile.scala 76:16:@149360.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@149359.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@149363.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@149357.4]
  assign regs_261_clock = clock; // @[:@149366.4]
  assign regs_261_reset = io_reset; // @[:@149367.4 RegFile.scala 76:16:@149374.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@149373.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@149377.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@149371.4]
  assign regs_262_clock = clock; // @[:@149380.4]
  assign regs_262_reset = io_reset; // @[:@149381.4 RegFile.scala 76:16:@149388.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@149387.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@149391.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@149385.4]
  assign regs_263_clock = clock; // @[:@149394.4]
  assign regs_263_reset = io_reset; // @[:@149395.4 RegFile.scala 76:16:@149402.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@149401.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@149405.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@149399.4]
  assign regs_264_clock = clock; // @[:@149408.4]
  assign regs_264_reset = io_reset; // @[:@149409.4 RegFile.scala 76:16:@149416.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@149415.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@149419.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@149413.4]
  assign regs_265_clock = clock; // @[:@149422.4]
  assign regs_265_reset = io_reset; // @[:@149423.4 RegFile.scala 76:16:@149430.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@149429.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@149433.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@149427.4]
  assign regs_266_clock = clock; // @[:@149436.4]
  assign regs_266_reset = io_reset; // @[:@149437.4 RegFile.scala 76:16:@149444.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@149443.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@149447.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@149441.4]
  assign regs_267_clock = clock; // @[:@149450.4]
  assign regs_267_reset = io_reset; // @[:@149451.4 RegFile.scala 76:16:@149458.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@149457.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@149461.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@149455.4]
  assign regs_268_clock = clock; // @[:@149464.4]
  assign regs_268_reset = io_reset; // @[:@149465.4 RegFile.scala 76:16:@149472.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@149471.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@149475.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@149469.4]
  assign regs_269_clock = clock; // @[:@149478.4]
  assign regs_269_reset = io_reset; // @[:@149479.4 RegFile.scala 76:16:@149486.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@149485.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@149489.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@149483.4]
  assign regs_270_clock = clock; // @[:@149492.4]
  assign regs_270_reset = io_reset; // @[:@149493.4 RegFile.scala 76:16:@149500.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@149499.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@149503.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@149497.4]
  assign regs_271_clock = clock; // @[:@149506.4]
  assign regs_271_reset = io_reset; // @[:@149507.4 RegFile.scala 76:16:@149514.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@149513.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@149517.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@149511.4]
  assign regs_272_clock = clock; // @[:@149520.4]
  assign regs_272_reset = io_reset; // @[:@149521.4 RegFile.scala 76:16:@149528.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@149527.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@149531.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@149525.4]
  assign regs_273_clock = clock; // @[:@149534.4]
  assign regs_273_reset = io_reset; // @[:@149535.4 RegFile.scala 76:16:@149542.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@149541.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@149545.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@149539.4]
  assign regs_274_clock = clock; // @[:@149548.4]
  assign regs_274_reset = io_reset; // @[:@149549.4 RegFile.scala 76:16:@149556.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@149555.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@149559.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@149553.4]
  assign regs_275_clock = clock; // @[:@149562.4]
  assign regs_275_reset = io_reset; // @[:@149563.4 RegFile.scala 76:16:@149570.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@149569.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@149573.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@149567.4]
  assign regs_276_clock = clock; // @[:@149576.4]
  assign regs_276_reset = io_reset; // @[:@149577.4 RegFile.scala 76:16:@149584.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@149583.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@149587.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@149581.4]
  assign regs_277_clock = clock; // @[:@149590.4]
  assign regs_277_reset = io_reset; // @[:@149591.4 RegFile.scala 76:16:@149598.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@149597.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@149601.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@149595.4]
  assign regs_278_clock = clock; // @[:@149604.4]
  assign regs_278_reset = io_reset; // @[:@149605.4 RegFile.scala 76:16:@149612.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@149611.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@149615.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@149609.4]
  assign regs_279_clock = clock; // @[:@149618.4]
  assign regs_279_reset = io_reset; // @[:@149619.4 RegFile.scala 76:16:@149626.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@149625.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@149629.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@149623.4]
  assign regs_280_clock = clock; // @[:@149632.4]
  assign regs_280_reset = io_reset; // @[:@149633.4 RegFile.scala 76:16:@149640.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@149639.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@149643.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@149637.4]
  assign regs_281_clock = clock; // @[:@149646.4]
  assign regs_281_reset = io_reset; // @[:@149647.4 RegFile.scala 76:16:@149654.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@149653.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@149657.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@149651.4]
  assign regs_282_clock = clock; // @[:@149660.4]
  assign regs_282_reset = io_reset; // @[:@149661.4 RegFile.scala 76:16:@149668.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@149667.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@149671.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@149665.4]
  assign regs_283_clock = clock; // @[:@149674.4]
  assign regs_283_reset = io_reset; // @[:@149675.4 RegFile.scala 76:16:@149682.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@149681.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@149685.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@149679.4]
  assign regs_284_clock = clock; // @[:@149688.4]
  assign regs_284_reset = io_reset; // @[:@149689.4 RegFile.scala 76:16:@149696.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@149695.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@149699.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@149693.4]
  assign regs_285_clock = clock; // @[:@149702.4]
  assign regs_285_reset = io_reset; // @[:@149703.4 RegFile.scala 76:16:@149710.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@149709.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@149713.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@149707.4]
  assign regs_286_clock = clock; // @[:@149716.4]
  assign regs_286_reset = io_reset; // @[:@149717.4 RegFile.scala 76:16:@149724.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@149723.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@149727.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@149721.4]
  assign regs_287_clock = clock; // @[:@149730.4]
  assign regs_287_reset = io_reset; // @[:@149731.4 RegFile.scala 76:16:@149738.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@149737.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@149741.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@149735.4]
  assign regs_288_clock = clock; // @[:@149744.4]
  assign regs_288_reset = io_reset; // @[:@149745.4 RegFile.scala 76:16:@149752.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@149751.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@149755.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@149749.4]
  assign regs_289_clock = clock; // @[:@149758.4]
  assign regs_289_reset = io_reset; // @[:@149759.4 RegFile.scala 76:16:@149766.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@149765.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@149769.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@149763.4]
  assign regs_290_clock = clock; // @[:@149772.4]
  assign regs_290_reset = io_reset; // @[:@149773.4 RegFile.scala 76:16:@149780.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@149779.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@149783.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@149777.4]
  assign regs_291_clock = clock; // @[:@149786.4]
  assign regs_291_reset = io_reset; // @[:@149787.4 RegFile.scala 76:16:@149794.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@149793.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@149797.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@149791.4]
  assign regs_292_clock = clock; // @[:@149800.4]
  assign regs_292_reset = io_reset; // @[:@149801.4 RegFile.scala 76:16:@149808.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@149807.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@149811.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@149805.4]
  assign regs_293_clock = clock; // @[:@149814.4]
  assign regs_293_reset = io_reset; // @[:@149815.4 RegFile.scala 76:16:@149822.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@149821.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@149825.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@149819.4]
  assign regs_294_clock = clock; // @[:@149828.4]
  assign regs_294_reset = io_reset; // @[:@149829.4 RegFile.scala 76:16:@149836.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@149835.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@149839.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@149833.4]
  assign regs_295_clock = clock; // @[:@149842.4]
  assign regs_295_reset = io_reset; // @[:@149843.4 RegFile.scala 76:16:@149850.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@149849.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@149853.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@149847.4]
  assign regs_296_clock = clock; // @[:@149856.4]
  assign regs_296_reset = io_reset; // @[:@149857.4 RegFile.scala 76:16:@149864.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@149863.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@149867.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@149861.4]
  assign regs_297_clock = clock; // @[:@149870.4]
  assign regs_297_reset = io_reset; // @[:@149871.4 RegFile.scala 76:16:@149878.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@149877.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@149881.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@149875.4]
  assign regs_298_clock = clock; // @[:@149884.4]
  assign regs_298_reset = io_reset; // @[:@149885.4 RegFile.scala 76:16:@149892.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@149891.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@149895.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@149889.4]
  assign regs_299_clock = clock; // @[:@149898.4]
  assign regs_299_reset = io_reset; // @[:@149899.4 RegFile.scala 76:16:@149906.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@149905.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@149909.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@149903.4]
  assign regs_300_clock = clock; // @[:@149912.4]
  assign regs_300_reset = io_reset; // @[:@149913.4 RegFile.scala 76:16:@149920.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@149919.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@149923.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@149917.4]
  assign regs_301_clock = clock; // @[:@149926.4]
  assign regs_301_reset = io_reset; // @[:@149927.4 RegFile.scala 76:16:@149934.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@149933.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@149937.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@149931.4]
  assign regs_302_clock = clock; // @[:@149940.4]
  assign regs_302_reset = io_reset; // @[:@149941.4 RegFile.scala 76:16:@149948.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@149947.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@149951.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@149945.4]
  assign regs_303_clock = clock; // @[:@149954.4]
  assign regs_303_reset = io_reset; // @[:@149955.4 RegFile.scala 76:16:@149962.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@149961.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@149965.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@149959.4]
  assign regs_304_clock = clock; // @[:@149968.4]
  assign regs_304_reset = io_reset; // @[:@149969.4 RegFile.scala 76:16:@149976.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@149975.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@149979.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@149973.4]
  assign regs_305_clock = clock; // @[:@149982.4]
  assign regs_305_reset = io_reset; // @[:@149983.4 RegFile.scala 76:16:@149990.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@149989.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@149993.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@149987.4]
  assign regs_306_clock = clock; // @[:@149996.4]
  assign regs_306_reset = io_reset; // @[:@149997.4 RegFile.scala 76:16:@150004.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@150003.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@150007.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@150001.4]
  assign regs_307_clock = clock; // @[:@150010.4]
  assign regs_307_reset = io_reset; // @[:@150011.4 RegFile.scala 76:16:@150018.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@150017.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@150021.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@150015.4]
  assign regs_308_clock = clock; // @[:@150024.4]
  assign regs_308_reset = io_reset; // @[:@150025.4 RegFile.scala 76:16:@150032.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@150031.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@150035.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@150029.4]
  assign regs_309_clock = clock; // @[:@150038.4]
  assign regs_309_reset = io_reset; // @[:@150039.4 RegFile.scala 76:16:@150046.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@150045.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@150049.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@150043.4]
  assign regs_310_clock = clock; // @[:@150052.4]
  assign regs_310_reset = io_reset; // @[:@150053.4 RegFile.scala 76:16:@150060.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@150059.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@150063.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@150057.4]
  assign regs_311_clock = clock; // @[:@150066.4]
  assign regs_311_reset = io_reset; // @[:@150067.4 RegFile.scala 76:16:@150074.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@150073.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@150077.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@150071.4]
  assign regs_312_clock = clock; // @[:@150080.4]
  assign regs_312_reset = io_reset; // @[:@150081.4 RegFile.scala 76:16:@150088.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@150087.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@150091.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@150085.4]
  assign regs_313_clock = clock; // @[:@150094.4]
  assign regs_313_reset = io_reset; // @[:@150095.4 RegFile.scala 76:16:@150102.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@150101.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@150105.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@150099.4]
  assign regs_314_clock = clock; // @[:@150108.4]
  assign regs_314_reset = io_reset; // @[:@150109.4 RegFile.scala 76:16:@150116.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@150115.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@150119.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@150113.4]
  assign regs_315_clock = clock; // @[:@150122.4]
  assign regs_315_reset = io_reset; // @[:@150123.4 RegFile.scala 76:16:@150130.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@150129.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@150133.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@150127.4]
  assign regs_316_clock = clock; // @[:@150136.4]
  assign regs_316_reset = io_reset; // @[:@150137.4 RegFile.scala 76:16:@150144.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@150143.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@150147.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@150141.4]
  assign regs_317_clock = clock; // @[:@150150.4]
  assign regs_317_reset = io_reset; // @[:@150151.4 RegFile.scala 76:16:@150158.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@150157.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@150161.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@150155.4]
  assign regs_318_clock = clock; // @[:@150164.4]
  assign regs_318_reset = io_reset; // @[:@150165.4 RegFile.scala 76:16:@150172.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@150171.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@150175.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@150169.4]
  assign regs_319_clock = clock; // @[:@150178.4]
  assign regs_319_reset = io_reset; // @[:@150179.4 RegFile.scala 76:16:@150186.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@150185.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@150189.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@150183.4]
  assign regs_320_clock = clock; // @[:@150192.4]
  assign regs_320_reset = io_reset; // @[:@150193.4 RegFile.scala 76:16:@150200.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@150199.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@150203.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@150197.4]
  assign regs_321_clock = clock; // @[:@150206.4]
  assign regs_321_reset = io_reset; // @[:@150207.4 RegFile.scala 76:16:@150214.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@150213.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@150217.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@150211.4]
  assign regs_322_clock = clock; // @[:@150220.4]
  assign regs_322_reset = io_reset; // @[:@150221.4 RegFile.scala 76:16:@150228.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@150227.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@150231.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@150225.4]
  assign regs_323_clock = clock; // @[:@150234.4]
  assign regs_323_reset = io_reset; // @[:@150235.4 RegFile.scala 76:16:@150242.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@150241.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@150245.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@150239.4]
  assign regs_324_clock = clock; // @[:@150248.4]
  assign regs_324_reset = io_reset; // @[:@150249.4 RegFile.scala 76:16:@150256.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@150255.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@150259.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@150253.4]
  assign regs_325_clock = clock; // @[:@150262.4]
  assign regs_325_reset = io_reset; // @[:@150263.4 RegFile.scala 76:16:@150270.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@150269.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@150273.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@150267.4]
  assign regs_326_clock = clock; // @[:@150276.4]
  assign regs_326_reset = io_reset; // @[:@150277.4 RegFile.scala 76:16:@150284.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@150283.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@150287.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@150281.4]
  assign regs_327_clock = clock; // @[:@150290.4]
  assign regs_327_reset = io_reset; // @[:@150291.4 RegFile.scala 76:16:@150298.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@150297.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@150301.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@150295.4]
  assign regs_328_clock = clock; // @[:@150304.4]
  assign regs_328_reset = io_reset; // @[:@150305.4 RegFile.scala 76:16:@150312.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@150311.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@150315.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@150309.4]
  assign regs_329_clock = clock; // @[:@150318.4]
  assign regs_329_reset = io_reset; // @[:@150319.4 RegFile.scala 76:16:@150326.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@150325.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@150329.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@150323.4]
  assign regs_330_clock = clock; // @[:@150332.4]
  assign regs_330_reset = io_reset; // @[:@150333.4 RegFile.scala 76:16:@150340.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@150339.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@150343.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@150337.4]
  assign regs_331_clock = clock; // @[:@150346.4]
  assign regs_331_reset = io_reset; // @[:@150347.4 RegFile.scala 76:16:@150354.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@150353.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@150357.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@150351.4]
  assign regs_332_clock = clock; // @[:@150360.4]
  assign regs_332_reset = io_reset; // @[:@150361.4 RegFile.scala 76:16:@150368.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@150367.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@150371.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@150365.4]
  assign regs_333_clock = clock; // @[:@150374.4]
  assign regs_333_reset = io_reset; // @[:@150375.4 RegFile.scala 76:16:@150382.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@150381.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@150385.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@150379.4]
  assign regs_334_clock = clock; // @[:@150388.4]
  assign regs_334_reset = io_reset; // @[:@150389.4 RegFile.scala 76:16:@150396.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@150395.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@150399.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@150393.4]
  assign regs_335_clock = clock; // @[:@150402.4]
  assign regs_335_reset = io_reset; // @[:@150403.4 RegFile.scala 76:16:@150410.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@150409.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@150413.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@150407.4]
  assign regs_336_clock = clock; // @[:@150416.4]
  assign regs_336_reset = io_reset; // @[:@150417.4 RegFile.scala 76:16:@150424.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@150423.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@150427.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@150421.4]
  assign regs_337_clock = clock; // @[:@150430.4]
  assign regs_337_reset = io_reset; // @[:@150431.4 RegFile.scala 76:16:@150438.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@150437.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@150441.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@150435.4]
  assign regs_338_clock = clock; // @[:@150444.4]
  assign regs_338_reset = io_reset; // @[:@150445.4 RegFile.scala 76:16:@150452.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@150451.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@150455.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@150449.4]
  assign regs_339_clock = clock; // @[:@150458.4]
  assign regs_339_reset = io_reset; // @[:@150459.4 RegFile.scala 76:16:@150466.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@150465.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@150469.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@150463.4]
  assign regs_340_clock = clock; // @[:@150472.4]
  assign regs_340_reset = io_reset; // @[:@150473.4 RegFile.scala 76:16:@150480.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@150479.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@150483.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@150477.4]
  assign regs_341_clock = clock; // @[:@150486.4]
  assign regs_341_reset = io_reset; // @[:@150487.4 RegFile.scala 76:16:@150494.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@150493.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@150497.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@150491.4]
  assign regs_342_clock = clock; // @[:@150500.4]
  assign regs_342_reset = io_reset; // @[:@150501.4 RegFile.scala 76:16:@150508.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@150507.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@150511.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@150505.4]
  assign regs_343_clock = clock; // @[:@150514.4]
  assign regs_343_reset = io_reset; // @[:@150515.4 RegFile.scala 76:16:@150522.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@150521.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@150525.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@150519.4]
  assign regs_344_clock = clock; // @[:@150528.4]
  assign regs_344_reset = io_reset; // @[:@150529.4 RegFile.scala 76:16:@150536.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@150535.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@150539.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@150533.4]
  assign regs_345_clock = clock; // @[:@150542.4]
  assign regs_345_reset = io_reset; // @[:@150543.4 RegFile.scala 76:16:@150550.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@150549.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@150553.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@150547.4]
  assign regs_346_clock = clock; // @[:@150556.4]
  assign regs_346_reset = io_reset; // @[:@150557.4 RegFile.scala 76:16:@150564.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@150563.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@150567.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@150561.4]
  assign regs_347_clock = clock; // @[:@150570.4]
  assign regs_347_reset = io_reset; // @[:@150571.4 RegFile.scala 76:16:@150578.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@150577.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@150581.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@150575.4]
  assign regs_348_clock = clock; // @[:@150584.4]
  assign regs_348_reset = io_reset; // @[:@150585.4 RegFile.scala 76:16:@150592.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@150591.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@150595.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@150589.4]
  assign regs_349_clock = clock; // @[:@150598.4]
  assign regs_349_reset = io_reset; // @[:@150599.4 RegFile.scala 76:16:@150606.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@150605.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@150609.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@150603.4]
  assign regs_350_clock = clock; // @[:@150612.4]
  assign regs_350_reset = io_reset; // @[:@150613.4 RegFile.scala 76:16:@150620.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@150619.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@150623.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@150617.4]
  assign regs_351_clock = clock; // @[:@150626.4]
  assign regs_351_reset = io_reset; // @[:@150627.4 RegFile.scala 76:16:@150634.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@150633.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@150637.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@150631.4]
  assign regs_352_clock = clock; // @[:@150640.4]
  assign regs_352_reset = io_reset; // @[:@150641.4 RegFile.scala 76:16:@150648.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@150647.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@150651.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@150645.4]
  assign regs_353_clock = clock; // @[:@150654.4]
  assign regs_353_reset = io_reset; // @[:@150655.4 RegFile.scala 76:16:@150662.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@150661.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@150665.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@150659.4]
  assign regs_354_clock = clock; // @[:@150668.4]
  assign regs_354_reset = io_reset; // @[:@150669.4 RegFile.scala 76:16:@150676.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@150675.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@150679.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@150673.4]
  assign regs_355_clock = clock; // @[:@150682.4]
  assign regs_355_reset = io_reset; // @[:@150683.4 RegFile.scala 76:16:@150690.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@150689.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@150693.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@150687.4]
  assign regs_356_clock = clock; // @[:@150696.4]
  assign regs_356_reset = io_reset; // @[:@150697.4 RegFile.scala 76:16:@150704.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@150703.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@150707.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@150701.4]
  assign regs_357_clock = clock; // @[:@150710.4]
  assign regs_357_reset = io_reset; // @[:@150711.4 RegFile.scala 76:16:@150718.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@150717.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@150721.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@150715.4]
  assign regs_358_clock = clock; // @[:@150724.4]
  assign regs_358_reset = io_reset; // @[:@150725.4 RegFile.scala 76:16:@150732.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@150731.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@150735.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@150729.4]
  assign regs_359_clock = clock; // @[:@150738.4]
  assign regs_359_reset = io_reset; // @[:@150739.4 RegFile.scala 76:16:@150746.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@150745.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@150749.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@150743.4]
  assign regs_360_clock = clock; // @[:@150752.4]
  assign regs_360_reset = io_reset; // @[:@150753.4 RegFile.scala 76:16:@150760.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@150759.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@150763.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@150757.4]
  assign regs_361_clock = clock; // @[:@150766.4]
  assign regs_361_reset = io_reset; // @[:@150767.4 RegFile.scala 76:16:@150774.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@150773.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@150777.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@150771.4]
  assign regs_362_clock = clock; // @[:@150780.4]
  assign regs_362_reset = io_reset; // @[:@150781.4 RegFile.scala 76:16:@150788.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@150787.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@150791.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@150785.4]
  assign regs_363_clock = clock; // @[:@150794.4]
  assign regs_363_reset = io_reset; // @[:@150795.4 RegFile.scala 76:16:@150802.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@150801.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@150805.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@150799.4]
  assign regs_364_clock = clock; // @[:@150808.4]
  assign regs_364_reset = io_reset; // @[:@150809.4 RegFile.scala 76:16:@150816.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@150815.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@150819.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@150813.4]
  assign regs_365_clock = clock; // @[:@150822.4]
  assign regs_365_reset = io_reset; // @[:@150823.4 RegFile.scala 76:16:@150830.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@150829.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@150833.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@150827.4]
  assign regs_366_clock = clock; // @[:@150836.4]
  assign regs_366_reset = io_reset; // @[:@150837.4 RegFile.scala 76:16:@150844.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@150843.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@150847.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@150841.4]
  assign regs_367_clock = clock; // @[:@150850.4]
  assign regs_367_reset = io_reset; // @[:@150851.4 RegFile.scala 76:16:@150858.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@150857.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@150861.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@150855.4]
  assign regs_368_clock = clock; // @[:@150864.4]
  assign regs_368_reset = io_reset; // @[:@150865.4 RegFile.scala 76:16:@150872.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@150871.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@150875.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@150869.4]
  assign regs_369_clock = clock; // @[:@150878.4]
  assign regs_369_reset = io_reset; // @[:@150879.4 RegFile.scala 76:16:@150886.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@150885.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@150889.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@150883.4]
  assign regs_370_clock = clock; // @[:@150892.4]
  assign regs_370_reset = io_reset; // @[:@150893.4 RegFile.scala 76:16:@150900.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@150899.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@150903.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@150897.4]
  assign regs_371_clock = clock; // @[:@150906.4]
  assign regs_371_reset = io_reset; // @[:@150907.4 RegFile.scala 76:16:@150914.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@150913.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@150917.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@150911.4]
  assign regs_372_clock = clock; // @[:@150920.4]
  assign regs_372_reset = io_reset; // @[:@150921.4 RegFile.scala 76:16:@150928.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@150927.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@150931.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@150925.4]
  assign regs_373_clock = clock; // @[:@150934.4]
  assign regs_373_reset = io_reset; // @[:@150935.4 RegFile.scala 76:16:@150942.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@150941.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@150945.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@150939.4]
  assign regs_374_clock = clock; // @[:@150948.4]
  assign regs_374_reset = io_reset; // @[:@150949.4 RegFile.scala 76:16:@150956.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@150955.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@150959.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@150953.4]
  assign regs_375_clock = clock; // @[:@150962.4]
  assign regs_375_reset = io_reset; // @[:@150963.4 RegFile.scala 76:16:@150970.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@150969.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@150973.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@150967.4]
  assign regs_376_clock = clock; // @[:@150976.4]
  assign regs_376_reset = io_reset; // @[:@150977.4 RegFile.scala 76:16:@150984.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@150983.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@150987.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@150981.4]
  assign regs_377_clock = clock; // @[:@150990.4]
  assign regs_377_reset = io_reset; // @[:@150991.4 RegFile.scala 76:16:@150998.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@150997.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@151001.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@150995.4]
  assign regs_378_clock = clock; // @[:@151004.4]
  assign regs_378_reset = io_reset; // @[:@151005.4 RegFile.scala 76:16:@151012.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@151011.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@151015.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@151009.4]
  assign regs_379_clock = clock; // @[:@151018.4]
  assign regs_379_reset = io_reset; // @[:@151019.4 RegFile.scala 76:16:@151026.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@151025.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@151029.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@151023.4]
  assign regs_380_clock = clock; // @[:@151032.4]
  assign regs_380_reset = io_reset; // @[:@151033.4 RegFile.scala 76:16:@151040.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@151039.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@151043.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@151037.4]
  assign regs_381_clock = clock; // @[:@151046.4]
  assign regs_381_reset = io_reset; // @[:@151047.4 RegFile.scala 76:16:@151054.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@151053.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@151057.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@151051.4]
  assign regs_382_clock = clock; // @[:@151060.4]
  assign regs_382_reset = io_reset; // @[:@151061.4 RegFile.scala 76:16:@151068.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@151067.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@151071.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@151065.4]
  assign regs_383_clock = clock; // @[:@151074.4]
  assign regs_383_reset = io_reset; // @[:@151075.4 RegFile.scala 76:16:@151082.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@151081.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@151085.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@151079.4]
  assign regs_384_clock = clock; // @[:@151088.4]
  assign regs_384_reset = io_reset; // @[:@151089.4 RegFile.scala 76:16:@151096.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@151095.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@151099.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@151093.4]
  assign regs_385_clock = clock; // @[:@151102.4]
  assign regs_385_reset = io_reset; // @[:@151103.4 RegFile.scala 76:16:@151110.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@151109.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@151113.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@151107.4]
  assign regs_386_clock = clock; // @[:@151116.4]
  assign regs_386_reset = io_reset; // @[:@151117.4 RegFile.scala 76:16:@151124.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@151123.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@151127.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@151121.4]
  assign regs_387_clock = clock; // @[:@151130.4]
  assign regs_387_reset = io_reset; // @[:@151131.4 RegFile.scala 76:16:@151138.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@151137.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@151141.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@151135.4]
  assign regs_388_clock = clock; // @[:@151144.4]
  assign regs_388_reset = io_reset; // @[:@151145.4 RegFile.scala 76:16:@151152.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@151151.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@151155.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@151149.4]
  assign regs_389_clock = clock; // @[:@151158.4]
  assign regs_389_reset = io_reset; // @[:@151159.4 RegFile.scala 76:16:@151166.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@151165.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@151169.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@151163.4]
  assign regs_390_clock = clock; // @[:@151172.4]
  assign regs_390_reset = io_reset; // @[:@151173.4 RegFile.scala 76:16:@151180.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@151179.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@151183.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@151177.4]
  assign regs_391_clock = clock; // @[:@151186.4]
  assign regs_391_reset = io_reset; // @[:@151187.4 RegFile.scala 76:16:@151194.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@151193.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@151197.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@151191.4]
  assign regs_392_clock = clock; // @[:@151200.4]
  assign regs_392_reset = io_reset; // @[:@151201.4 RegFile.scala 76:16:@151208.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@151207.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@151211.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@151205.4]
  assign regs_393_clock = clock; // @[:@151214.4]
  assign regs_393_reset = io_reset; // @[:@151215.4 RegFile.scala 76:16:@151222.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@151221.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@151225.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@151219.4]
  assign regs_394_clock = clock; // @[:@151228.4]
  assign regs_394_reset = io_reset; // @[:@151229.4 RegFile.scala 76:16:@151236.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@151235.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@151239.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@151233.4]
  assign regs_395_clock = clock; // @[:@151242.4]
  assign regs_395_reset = io_reset; // @[:@151243.4 RegFile.scala 76:16:@151250.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@151249.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@151253.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@151247.4]
  assign regs_396_clock = clock; // @[:@151256.4]
  assign regs_396_reset = io_reset; // @[:@151257.4 RegFile.scala 76:16:@151264.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@151263.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@151267.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@151261.4]
  assign regs_397_clock = clock; // @[:@151270.4]
  assign regs_397_reset = io_reset; // @[:@151271.4 RegFile.scala 76:16:@151278.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@151277.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@151281.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@151275.4]
  assign regs_398_clock = clock; // @[:@151284.4]
  assign regs_398_reset = io_reset; // @[:@151285.4 RegFile.scala 76:16:@151292.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@151291.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@151295.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@151289.4]
  assign regs_399_clock = clock; // @[:@151298.4]
  assign regs_399_reset = io_reset; // @[:@151299.4 RegFile.scala 76:16:@151306.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@151305.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@151309.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@151303.4]
  assign regs_400_clock = clock; // @[:@151312.4]
  assign regs_400_reset = io_reset; // @[:@151313.4 RegFile.scala 76:16:@151320.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@151319.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@151323.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@151317.4]
  assign regs_401_clock = clock; // @[:@151326.4]
  assign regs_401_reset = io_reset; // @[:@151327.4 RegFile.scala 76:16:@151334.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@151333.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@151337.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@151331.4]
  assign regs_402_clock = clock; // @[:@151340.4]
  assign regs_402_reset = io_reset; // @[:@151341.4 RegFile.scala 76:16:@151348.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@151347.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@151351.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@151345.4]
  assign regs_403_clock = clock; // @[:@151354.4]
  assign regs_403_reset = io_reset; // @[:@151355.4 RegFile.scala 76:16:@151362.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@151361.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@151365.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@151359.4]
  assign regs_404_clock = clock; // @[:@151368.4]
  assign regs_404_reset = io_reset; // @[:@151369.4 RegFile.scala 76:16:@151376.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@151375.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@151379.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@151373.4]
  assign regs_405_clock = clock; // @[:@151382.4]
  assign regs_405_reset = io_reset; // @[:@151383.4 RegFile.scala 76:16:@151390.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@151389.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@151393.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@151387.4]
  assign regs_406_clock = clock; // @[:@151396.4]
  assign regs_406_reset = io_reset; // @[:@151397.4 RegFile.scala 76:16:@151404.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@151403.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@151407.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@151401.4]
  assign regs_407_clock = clock; // @[:@151410.4]
  assign regs_407_reset = io_reset; // @[:@151411.4 RegFile.scala 76:16:@151418.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@151417.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@151421.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@151415.4]
  assign regs_408_clock = clock; // @[:@151424.4]
  assign regs_408_reset = io_reset; // @[:@151425.4 RegFile.scala 76:16:@151432.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@151431.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@151435.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@151429.4]
  assign regs_409_clock = clock; // @[:@151438.4]
  assign regs_409_reset = io_reset; // @[:@151439.4 RegFile.scala 76:16:@151446.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@151445.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@151449.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@151443.4]
  assign regs_410_clock = clock; // @[:@151452.4]
  assign regs_410_reset = io_reset; // @[:@151453.4 RegFile.scala 76:16:@151460.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@151459.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@151463.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@151457.4]
  assign regs_411_clock = clock; // @[:@151466.4]
  assign regs_411_reset = io_reset; // @[:@151467.4 RegFile.scala 76:16:@151474.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@151473.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@151477.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@151471.4]
  assign regs_412_clock = clock; // @[:@151480.4]
  assign regs_412_reset = io_reset; // @[:@151481.4 RegFile.scala 76:16:@151488.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@151487.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@151491.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@151485.4]
  assign regs_413_clock = clock; // @[:@151494.4]
  assign regs_413_reset = io_reset; // @[:@151495.4 RegFile.scala 76:16:@151502.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@151501.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@151505.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@151499.4]
  assign regs_414_clock = clock; // @[:@151508.4]
  assign regs_414_reset = io_reset; // @[:@151509.4 RegFile.scala 76:16:@151516.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@151515.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@151519.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@151513.4]
  assign regs_415_clock = clock; // @[:@151522.4]
  assign regs_415_reset = io_reset; // @[:@151523.4 RegFile.scala 76:16:@151530.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@151529.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@151533.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@151527.4]
  assign regs_416_clock = clock; // @[:@151536.4]
  assign regs_416_reset = io_reset; // @[:@151537.4 RegFile.scala 76:16:@151544.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@151543.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@151547.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@151541.4]
  assign regs_417_clock = clock; // @[:@151550.4]
  assign regs_417_reset = io_reset; // @[:@151551.4 RegFile.scala 76:16:@151558.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@151557.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@151561.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@151555.4]
  assign regs_418_clock = clock; // @[:@151564.4]
  assign regs_418_reset = io_reset; // @[:@151565.4 RegFile.scala 76:16:@151572.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@151571.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@151575.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@151569.4]
  assign regs_419_clock = clock; // @[:@151578.4]
  assign regs_419_reset = io_reset; // @[:@151579.4 RegFile.scala 76:16:@151586.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@151585.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@151589.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@151583.4]
  assign regs_420_clock = clock; // @[:@151592.4]
  assign regs_420_reset = io_reset; // @[:@151593.4 RegFile.scala 76:16:@151600.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@151599.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@151603.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@151597.4]
  assign regs_421_clock = clock; // @[:@151606.4]
  assign regs_421_reset = io_reset; // @[:@151607.4 RegFile.scala 76:16:@151614.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@151613.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@151617.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@151611.4]
  assign regs_422_clock = clock; // @[:@151620.4]
  assign regs_422_reset = io_reset; // @[:@151621.4 RegFile.scala 76:16:@151628.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@151627.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@151631.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@151625.4]
  assign regs_423_clock = clock; // @[:@151634.4]
  assign regs_423_reset = io_reset; // @[:@151635.4 RegFile.scala 76:16:@151642.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@151641.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@151645.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@151639.4]
  assign regs_424_clock = clock; // @[:@151648.4]
  assign regs_424_reset = io_reset; // @[:@151649.4 RegFile.scala 76:16:@151656.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@151655.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@151659.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@151653.4]
  assign regs_425_clock = clock; // @[:@151662.4]
  assign regs_425_reset = io_reset; // @[:@151663.4 RegFile.scala 76:16:@151670.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@151669.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@151673.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@151667.4]
  assign regs_426_clock = clock; // @[:@151676.4]
  assign regs_426_reset = io_reset; // @[:@151677.4 RegFile.scala 76:16:@151684.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@151683.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@151687.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@151681.4]
  assign regs_427_clock = clock; // @[:@151690.4]
  assign regs_427_reset = io_reset; // @[:@151691.4 RegFile.scala 76:16:@151698.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@151697.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@151701.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@151695.4]
  assign regs_428_clock = clock; // @[:@151704.4]
  assign regs_428_reset = io_reset; // @[:@151705.4 RegFile.scala 76:16:@151712.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@151711.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@151715.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@151709.4]
  assign regs_429_clock = clock; // @[:@151718.4]
  assign regs_429_reset = io_reset; // @[:@151719.4 RegFile.scala 76:16:@151726.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@151725.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@151729.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@151723.4]
  assign regs_430_clock = clock; // @[:@151732.4]
  assign regs_430_reset = io_reset; // @[:@151733.4 RegFile.scala 76:16:@151740.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@151739.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@151743.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@151737.4]
  assign regs_431_clock = clock; // @[:@151746.4]
  assign regs_431_reset = io_reset; // @[:@151747.4 RegFile.scala 76:16:@151754.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@151753.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@151757.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@151751.4]
  assign regs_432_clock = clock; // @[:@151760.4]
  assign regs_432_reset = io_reset; // @[:@151761.4 RegFile.scala 76:16:@151768.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@151767.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@151771.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@151765.4]
  assign regs_433_clock = clock; // @[:@151774.4]
  assign regs_433_reset = io_reset; // @[:@151775.4 RegFile.scala 76:16:@151782.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@151781.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@151785.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@151779.4]
  assign regs_434_clock = clock; // @[:@151788.4]
  assign regs_434_reset = io_reset; // @[:@151789.4 RegFile.scala 76:16:@151796.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@151795.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@151799.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@151793.4]
  assign regs_435_clock = clock; // @[:@151802.4]
  assign regs_435_reset = io_reset; // @[:@151803.4 RegFile.scala 76:16:@151810.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@151809.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@151813.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@151807.4]
  assign regs_436_clock = clock; // @[:@151816.4]
  assign regs_436_reset = io_reset; // @[:@151817.4 RegFile.scala 76:16:@151824.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@151823.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@151827.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@151821.4]
  assign regs_437_clock = clock; // @[:@151830.4]
  assign regs_437_reset = io_reset; // @[:@151831.4 RegFile.scala 76:16:@151838.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@151837.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@151841.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@151835.4]
  assign regs_438_clock = clock; // @[:@151844.4]
  assign regs_438_reset = io_reset; // @[:@151845.4 RegFile.scala 76:16:@151852.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@151851.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@151855.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@151849.4]
  assign regs_439_clock = clock; // @[:@151858.4]
  assign regs_439_reset = io_reset; // @[:@151859.4 RegFile.scala 76:16:@151866.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@151865.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@151869.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@151863.4]
  assign regs_440_clock = clock; // @[:@151872.4]
  assign regs_440_reset = io_reset; // @[:@151873.4 RegFile.scala 76:16:@151880.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@151879.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@151883.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@151877.4]
  assign regs_441_clock = clock; // @[:@151886.4]
  assign regs_441_reset = io_reset; // @[:@151887.4 RegFile.scala 76:16:@151894.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@151893.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@151897.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@151891.4]
  assign regs_442_clock = clock; // @[:@151900.4]
  assign regs_442_reset = io_reset; // @[:@151901.4 RegFile.scala 76:16:@151908.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@151907.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@151911.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@151905.4]
  assign regs_443_clock = clock; // @[:@151914.4]
  assign regs_443_reset = io_reset; // @[:@151915.4 RegFile.scala 76:16:@151922.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@151921.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@151925.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@151919.4]
  assign regs_444_clock = clock; // @[:@151928.4]
  assign regs_444_reset = io_reset; // @[:@151929.4 RegFile.scala 76:16:@151936.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@151935.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@151939.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@151933.4]
  assign regs_445_clock = clock; // @[:@151942.4]
  assign regs_445_reset = io_reset; // @[:@151943.4 RegFile.scala 76:16:@151950.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@151949.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@151953.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@151947.4]
  assign regs_446_clock = clock; // @[:@151956.4]
  assign regs_446_reset = io_reset; // @[:@151957.4 RegFile.scala 76:16:@151964.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@151963.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@151967.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@151961.4]
  assign regs_447_clock = clock; // @[:@151970.4]
  assign regs_447_reset = io_reset; // @[:@151971.4 RegFile.scala 76:16:@151978.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@151977.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@151981.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@151975.4]
  assign regs_448_clock = clock; // @[:@151984.4]
  assign regs_448_reset = io_reset; // @[:@151985.4 RegFile.scala 76:16:@151992.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@151991.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@151995.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@151989.4]
  assign regs_449_clock = clock; // @[:@151998.4]
  assign regs_449_reset = io_reset; // @[:@151999.4 RegFile.scala 76:16:@152006.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@152005.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@152009.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@152003.4]
  assign regs_450_clock = clock; // @[:@152012.4]
  assign regs_450_reset = io_reset; // @[:@152013.4 RegFile.scala 76:16:@152020.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@152019.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@152023.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@152017.4]
  assign regs_451_clock = clock; // @[:@152026.4]
  assign regs_451_reset = io_reset; // @[:@152027.4 RegFile.scala 76:16:@152034.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@152033.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@152037.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@152031.4]
  assign regs_452_clock = clock; // @[:@152040.4]
  assign regs_452_reset = io_reset; // @[:@152041.4 RegFile.scala 76:16:@152048.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@152047.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@152051.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@152045.4]
  assign regs_453_clock = clock; // @[:@152054.4]
  assign regs_453_reset = io_reset; // @[:@152055.4 RegFile.scala 76:16:@152062.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@152061.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@152065.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@152059.4]
  assign regs_454_clock = clock; // @[:@152068.4]
  assign regs_454_reset = io_reset; // @[:@152069.4 RegFile.scala 76:16:@152076.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@152075.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@152079.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@152073.4]
  assign regs_455_clock = clock; // @[:@152082.4]
  assign regs_455_reset = io_reset; // @[:@152083.4 RegFile.scala 76:16:@152090.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@152089.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@152093.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@152087.4]
  assign regs_456_clock = clock; // @[:@152096.4]
  assign regs_456_reset = io_reset; // @[:@152097.4 RegFile.scala 76:16:@152104.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@152103.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@152107.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@152101.4]
  assign regs_457_clock = clock; // @[:@152110.4]
  assign regs_457_reset = io_reset; // @[:@152111.4 RegFile.scala 76:16:@152118.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@152117.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@152121.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@152115.4]
  assign regs_458_clock = clock; // @[:@152124.4]
  assign regs_458_reset = io_reset; // @[:@152125.4 RegFile.scala 76:16:@152132.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@152131.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@152135.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@152129.4]
  assign regs_459_clock = clock; // @[:@152138.4]
  assign regs_459_reset = io_reset; // @[:@152139.4 RegFile.scala 76:16:@152146.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@152145.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@152149.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@152143.4]
  assign regs_460_clock = clock; // @[:@152152.4]
  assign regs_460_reset = io_reset; // @[:@152153.4 RegFile.scala 76:16:@152160.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@152159.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@152163.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@152157.4]
  assign regs_461_clock = clock; // @[:@152166.4]
  assign regs_461_reset = io_reset; // @[:@152167.4 RegFile.scala 76:16:@152174.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@152173.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@152177.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@152171.4]
  assign regs_462_clock = clock; // @[:@152180.4]
  assign regs_462_reset = io_reset; // @[:@152181.4 RegFile.scala 76:16:@152188.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@152187.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@152191.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@152185.4]
  assign regs_463_clock = clock; // @[:@152194.4]
  assign regs_463_reset = io_reset; // @[:@152195.4 RegFile.scala 76:16:@152202.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@152201.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@152205.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@152199.4]
  assign regs_464_clock = clock; // @[:@152208.4]
  assign regs_464_reset = io_reset; // @[:@152209.4 RegFile.scala 76:16:@152216.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@152215.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@152219.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@152213.4]
  assign regs_465_clock = clock; // @[:@152222.4]
  assign regs_465_reset = io_reset; // @[:@152223.4 RegFile.scala 76:16:@152230.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@152229.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@152233.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@152227.4]
  assign regs_466_clock = clock; // @[:@152236.4]
  assign regs_466_reset = io_reset; // @[:@152237.4 RegFile.scala 76:16:@152244.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@152243.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@152247.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@152241.4]
  assign regs_467_clock = clock; // @[:@152250.4]
  assign regs_467_reset = io_reset; // @[:@152251.4 RegFile.scala 76:16:@152258.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@152257.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@152261.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@152255.4]
  assign regs_468_clock = clock; // @[:@152264.4]
  assign regs_468_reset = io_reset; // @[:@152265.4 RegFile.scala 76:16:@152272.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@152271.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@152275.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@152269.4]
  assign regs_469_clock = clock; // @[:@152278.4]
  assign regs_469_reset = io_reset; // @[:@152279.4 RegFile.scala 76:16:@152286.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@152285.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@152289.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@152283.4]
  assign regs_470_clock = clock; // @[:@152292.4]
  assign regs_470_reset = io_reset; // @[:@152293.4 RegFile.scala 76:16:@152300.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@152299.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@152303.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@152297.4]
  assign regs_471_clock = clock; // @[:@152306.4]
  assign regs_471_reset = io_reset; // @[:@152307.4 RegFile.scala 76:16:@152314.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@152313.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@152317.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@152311.4]
  assign regs_472_clock = clock; // @[:@152320.4]
  assign regs_472_reset = io_reset; // @[:@152321.4 RegFile.scala 76:16:@152328.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@152327.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@152331.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@152325.4]
  assign regs_473_clock = clock; // @[:@152334.4]
  assign regs_473_reset = io_reset; // @[:@152335.4 RegFile.scala 76:16:@152342.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@152341.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@152345.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@152339.4]
  assign regs_474_clock = clock; // @[:@152348.4]
  assign regs_474_reset = io_reset; // @[:@152349.4 RegFile.scala 76:16:@152356.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@152355.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@152359.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@152353.4]
  assign regs_475_clock = clock; // @[:@152362.4]
  assign regs_475_reset = io_reset; // @[:@152363.4 RegFile.scala 76:16:@152370.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@152369.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@152373.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@152367.4]
  assign regs_476_clock = clock; // @[:@152376.4]
  assign regs_476_reset = io_reset; // @[:@152377.4 RegFile.scala 76:16:@152384.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@152383.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@152387.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@152381.4]
  assign regs_477_clock = clock; // @[:@152390.4]
  assign regs_477_reset = io_reset; // @[:@152391.4 RegFile.scala 76:16:@152398.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@152397.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@152401.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@152395.4]
  assign regs_478_clock = clock; // @[:@152404.4]
  assign regs_478_reset = io_reset; // @[:@152405.4 RegFile.scala 76:16:@152412.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@152411.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@152415.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@152409.4]
  assign regs_479_clock = clock; // @[:@152418.4]
  assign regs_479_reset = io_reset; // @[:@152419.4 RegFile.scala 76:16:@152426.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@152425.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@152429.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@152423.4]
  assign regs_480_clock = clock; // @[:@152432.4]
  assign regs_480_reset = io_reset; // @[:@152433.4 RegFile.scala 76:16:@152440.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@152439.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@152443.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@152437.4]
  assign regs_481_clock = clock; // @[:@152446.4]
  assign regs_481_reset = io_reset; // @[:@152447.4 RegFile.scala 76:16:@152454.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@152453.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@152457.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@152451.4]
  assign regs_482_clock = clock; // @[:@152460.4]
  assign regs_482_reset = io_reset; // @[:@152461.4 RegFile.scala 76:16:@152468.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@152467.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@152471.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@152465.4]
  assign regs_483_clock = clock; // @[:@152474.4]
  assign regs_483_reset = io_reset; // @[:@152475.4 RegFile.scala 76:16:@152482.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@152481.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@152485.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@152479.4]
  assign regs_484_clock = clock; // @[:@152488.4]
  assign regs_484_reset = io_reset; // @[:@152489.4 RegFile.scala 76:16:@152496.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@152495.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@152499.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@152493.4]
  assign regs_485_clock = clock; // @[:@152502.4]
  assign regs_485_reset = io_reset; // @[:@152503.4 RegFile.scala 76:16:@152510.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@152509.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@152513.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@152507.4]
  assign regs_486_clock = clock; // @[:@152516.4]
  assign regs_486_reset = io_reset; // @[:@152517.4 RegFile.scala 76:16:@152524.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@152523.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@152527.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@152521.4]
  assign regs_487_clock = clock; // @[:@152530.4]
  assign regs_487_reset = io_reset; // @[:@152531.4 RegFile.scala 76:16:@152538.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@152537.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@152541.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@152535.4]
  assign regs_488_clock = clock; // @[:@152544.4]
  assign regs_488_reset = io_reset; // @[:@152545.4 RegFile.scala 76:16:@152552.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@152551.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@152555.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@152549.4]
  assign regs_489_clock = clock; // @[:@152558.4]
  assign regs_489_reset = io_reset; // @[:@152559.4 RegFile.scala 76:16:@152566.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@152565.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@152569.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@152563.4]
  assign regs_490_clock = clock; // @[:@152572.4]
  assign regs_490_reset = io_reset; // @[:@152573.4 RegFile.scala 76:16:@152580.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@152579.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@152583.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@152577.4]
  assign regs_491_clock = clock; // @[:@152586.4]
  assign regs_491_reset = io_reset; // @[:@152587.4 RegFile.scala 76:16:@152594.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@152593.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@152597.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@152591.4]
  assign regs_492_clock = clock; // @[:@152600.4]
  assign regs_492_reset = io_reset; // @[:@152601.4 RegFile.scala 76:16:@152608.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@152607.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@152611.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@152605.4]
  assign regs_493_clock = clock; // @[:@152614.4]
  assign regs_493_reset = io_reset; // @[:@152615.4 RegFile.scala 76:16:@152622.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@152621.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@152625.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@152619.4]
  assign regs_494_clock = clock; // @[:@152628.4]
  assign regs_494_reset = io_reset; // @[:@152629.4 RegFile.scala 76:16:@152636.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@152635.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@152639.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@152633.4]
  assign regs_495_clock = clock; // @[:@152642.4]
  assign regs_495_reset = io_reset; // @[:@152643.4 RegFile.scala 76:16:@152650.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@152649.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@152653.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@152647.4]
  assign regs_496_clock = clock; // @[:@152656.4]
  assign regs_496_reset = io_reset; // @[:@152657.4 RegFile.scala 76:16:@152664.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@152663.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@152667.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@152661.4]
  assign regs_497_clock = clock; // @[:@152670.4]
  assign regs_497_reset = io_reset; // @[:@152671.4 RegFile.scala 76:16:@152678.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@152677.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@152681.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@152675.4]
  assign regs_498_clock = clock; // @[:@152684.4]
  assign regs_498_reset = io_reset; // @[:@152685.4 RegFile.scala 76:16:@152692.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@152691.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@152695.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@152689.4]
  assign regs_499_clock = clock; // @[:@152698.4]
  assign regs_499_reset = io_reset; // @[:@152699.4 RegFile.scala 76:16:@152706.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@152705.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@152709.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@152703.4]
  assign regs_500_clock = clock; // @[:@152712.4]
  assign regs_500_reset = io_reset; // @[:@152713.4 RegFile.scala 76:16:@152720.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@152719.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@152723.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@152717.4]
  assign regs_501_clock = clock; // @[:@152726.4]
  assign regs_501_reset = io_reset; // @[:@152727.4 RegFile.scala 76:16:@152734.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@152733.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@152737.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@152731.4]
  assign regs_502_clock = clock; // @[:@152740.4]
  assign regs_502_reset = io_reset; // @[:@152741.4 RegFile.scala 76:16:@152748.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@152747.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@152751.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@152745.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@153260.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@153261.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@153262.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@153263.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@153264.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@153265.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@153266.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@153267.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@153268.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@153269.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@153270.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@153271.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@153272.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@153273.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@153274.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@153275.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@153276.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@153277.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@153278.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@153279.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@153280.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@153281.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@153282.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@153283.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@153284.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@153285.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@153286.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@153287.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@153288.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@153289.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@153290.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@153291.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@153292.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@153293.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@153294.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@153295.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@153296.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@153297.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@153298.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@153299.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@153300.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@153301.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@153302.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@153303.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@153304.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@153305.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@153306.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@153307.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@153308.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@153309.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@153310.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@153311.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@153312.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@153313.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@153314.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@153315.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@153316.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@153317.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@153318.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@153319.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@153320.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@153321.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@153322.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@153323.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@153324.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@153325.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@153326.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@153327.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@153328.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@153329.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@153330.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@153331.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@153332.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@153333.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@153334.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@153335.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@153336.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@153337.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@153338.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@153339.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@153340.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@153341.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@153342.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@153343.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@153344.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@153345.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@153346.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@153347.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@153348.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@153349.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@153350.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@153351.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@153352.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@153353.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@153354.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@153355.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@153356.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@153357.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@153358.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@153359.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@153360.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@153361.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@153362.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@153363.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@153364.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@153365.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@153366.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@153367.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@153368.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@153369.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@153370.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@153371.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@153372.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@153373.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@153374.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@153375.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@153376.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@153377.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@153378.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@153379.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@153380.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@153381.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@153382.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@153383.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@153384.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@153385.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@153386.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@153387.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@153388.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@153389.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@153390.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@153391.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@153392.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@153393.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@153394.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@153395.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@153396.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@153397.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@153398.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@153399.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@153400.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@153401.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@153402.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@153403.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@153404.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@153405.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@153406.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@153407.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@153408.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@153409.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@153410.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@153411.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@153412.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@153413.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@153414.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@153415.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@153416.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@153417.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@153418.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@153419.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@153420.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@153421.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@153422.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@153423.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@153424.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@153425.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@153426.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@153427.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@153428.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@153429.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@153430.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@153431.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@153432.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@153433.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@153434.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@153435.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@153436.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@153437.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@153438.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@153439.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@153440.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@153441.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@153442.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@153443.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@153444.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@153445.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@153446.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@153447.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@153448.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@153449.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@153450.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@153451.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@153452.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@153453.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@153454.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@153455.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@153456.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@153457.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@153458.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@153459.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@153460.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@153461.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@153462.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@153463.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@153464.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@153465.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@153466.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@153467.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@153468.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@153469.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@153470.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@153471.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@153472.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@153473.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@153474.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@153475.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@153476.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@153477.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@153478.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@153479.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@153480.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@153481.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@153482.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@153483.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@153484.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@153485.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@153486.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@153487.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@153488.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@153489.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@153490.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@153491.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@153492.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@153493.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@153494.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@153495.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@153496.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@153497.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@153498.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@153499.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@153500.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@153501.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@153502.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@153503.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@153504.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@153505.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@153506.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@153507.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@153508.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@153509.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@153510.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@153511.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@153512.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@153513.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@153514.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@153515.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@153516.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@153517.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@153518.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@153519.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@153520.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@153521.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@153522.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@153523.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@153524.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@153525.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@153526.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@153527.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@153528.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@153529.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@153530.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@153531.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@153532.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@153533.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@153534.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@153535.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@153536.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@153537.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@153538.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@153539.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@153540.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@153541.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@153542.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@153543.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@153544.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@153545.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@153546.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@153547.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@153548.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@153549.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@153550.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@153551.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@153552.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@153553.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@153554.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@153555.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@153556.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@153557.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@153558.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@153559.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@153560.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@153561.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@153562.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@153563.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@153564.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@153565.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@153566.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@153567.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@153568.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@153569.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@153570.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@153571.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@153572.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@153573.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@153574.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@153575.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@153576.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@153577.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@153578.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@153579.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@153580.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@153581.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@153582.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@153583.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@153584.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@153585.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@153586.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@153587.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@153588.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@153589.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@153590.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@153591.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@153592.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@153593.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@153594.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@153595.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@153596.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@153597.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@153598.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@153599.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@153600.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@153601.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@153602.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@153603.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@153604.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@153605.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@153606.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@153607.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@153608.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@153609.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@153610.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@153611.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@153612.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@153613.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@153614.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@153615.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@153616.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@153617.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@153618.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@153619.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@153620.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@153621.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@153622.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@153623.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@153624.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@153625.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@153626.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@153627.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@153628.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@153629.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@153630.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@153631.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@153632.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@153633.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@153634.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@153635.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@153636.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@153637.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@153638.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@153639.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@153640.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@153641.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@153642.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@153643.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@153644.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@153645.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@153646.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@153647.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@153648.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@153649.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@153650.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@153651.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@153652.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@153653.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@153654.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@153655.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@153656.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@153657.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@153658.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@153659.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@153660.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@153661.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@153662.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@153663.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@153664.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@153665.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@153666.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@153667.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@153668.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@153669.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@153670.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@153671.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@153672.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@153673.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@153674.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@153675.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@153676.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@153677.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@153678.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@153679.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@153680.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@153681.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@153682.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@153683.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@153684.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@153685.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@153686.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@153687.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@153688.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@153689.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@153690.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@153691.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@153692.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@153693.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@153694.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@153695.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@153696.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@153697.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@153698.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@153699.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@153700.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@153701.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@153702.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@153703.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@153704.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@153705.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@153706.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@153707.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@153708.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@153709.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@153710.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@153711.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@153712.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@153713.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@153714.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@153715.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@153716.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@153717.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@153718.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@153719.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@153720.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@153721.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@153722.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@153723.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@153724.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@153725.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@153726.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@153727.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@153728.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@153729.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@153730.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@153731.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@153732.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@153733.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@153734.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@153735.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@153736.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@153737.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@153738.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@153739.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@153740.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@153741.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@153742.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@153743.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@153744.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@153745.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@153746.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@153747.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@153748.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@153749.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@153750.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@153751.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@153752.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@153753.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@153754.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@153755.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@153756.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@153757.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@153758.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@153759.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@153760.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@153761.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@153762.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@153763.4]
endmodule
module RetimeWrapper_1044( // @[:@153787.2]
  input         clock, // @[:@153788.4]
  input         reset, // @[:@153789.4]
  input  [39:0] io_in, // @[:@153790.4]
  output [39:0] io_out // @[:@153790.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@153792.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@153792.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@153792.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@153792.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@153792.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@153792.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@153792.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@153805.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@153804.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@153803.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@153802.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@153801.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@153799.4]
endmodule
module FringeFF_503( // @[:@153807.2]
  input         clock, // @[:@153808.4]
  input         reset, // @[:@153809.4]
  input  [39:0] io_in, // @[:@153810.4]
  output [39:0] io_out, // @[:@153810.4]
  input         io_enable // @[:@153810.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@153813.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@153813.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@153813.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@153813.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@153818.4 package.scala 96:25:@153819.4]
  RetimeWrapper_1044 RetimeWrapper ( // @[package.scala 93:22:@153813.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@153818.4 package.scala 96:25:@153819.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@153830.4]
  assign RetimeWrapper_clock = clock; // @[:@153814.4]
  assign RetimeWrapper_reset = reset; // @[:@153815.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@153816.4]
endmodule
module FringeCounter( // @[:@153832.2]
  input   clock, // @[:@153833.4]
  input   reset, // @[:@153834.4]
  input   io_enable, // @[:@153835.4]
  output  io_done // @[:@153835.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@153837.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@153837.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@153837.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@153837.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@153837.4]
  wire [40:0] count; // @[Cat.scala 30:58:@153844.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@153845.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@153846.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@153847.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@153849.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@153837.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@153844.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@153845.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@153846.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@153847.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@153849.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@153860.4]
  assign reg$_clock = clock; // @[:@153838.4]
  assign reg$_reset = reset; // @[:@153839.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@153851.6 FringeCounter.scala 37:15:@153854.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@153842.4]
endmodule
module FringeFF_504( // @[:@153894.2]
  input   clock, // @[:@153895.4]
  input   reset, // @[:@153896.4]
  input   io_in, // @[:@153897.4]
  input   io_reset, // @[:@153897.4]
  output  io_out, // @[:@153897.4]
  input   io_enable // @[:@153897.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@153900.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@153900.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@153900.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@153900.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@153900.4]
  wire  _T_18; // @[package.scala 96:25:@153905.4 package.scala 96:25:@153906.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@153911.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@153900.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@153905.4 package.scala 96:25:@153906.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@153911.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@153917.4]
  assign RetimeWrapper_clock = clock; // @[:@153901.4]
  assign RetimeWrapper_reset = reset; // @[:@153902.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@153904.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@153903.4]
endmodule
module Depulser( // @[:@153919.2]
  input   clock, // @[:@153920.4]
  input   reset, // @[:@153921.4]
  input   io_in, // @[:@153922.4]
  input   io_rst, // @[:@153922.4]
  output  io_out // @[:@153922.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@153924.4]
  wire  r_reset; // @[Depulser.scala 14:17:@153924.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@153924.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@153924.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@153924.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@153924.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@153924.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@153933.4]
  assign r_clock = clock; // @[:@153925.4]
  assign r_reset = reset; // @[:@153926.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@153928.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@153932.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@153931.4]
endmodule
module Fringe( // @[:@153935.2]
  input         clock, // @[:@153936.4]
  input         reset, // @[:@153937.4]
  input  [31:0] io_raddr, // @[:@153938.4]
  input         io_wen, // @[:@153938.4]
  input  [31:0] io_waddr, // @[:@153938.4]
  input  [63:0] io_wdata, // @[:@153938.4]
  output [63:0] io_rdata, // @[:@153938.4]
  output        io_enable, // @[:@153938.4]
  input         io_done, // @[:@153938.4]
  output        io_reset, // @[:@153938.4]
  output [63:0] io_argIns_0, // @[:@153938.4]
  output [63:0] io_argIns_1, // @[:@153938.4]
  input         io_argOuts_0_valid, // @[:@153938.4]
  input  [63:0] io_argOuts_0_bits, // @[:@153938.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@153938.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@153938.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@153938.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@153938.4]
  output        io_memStreams_stores_0_data_ready, // @[:@153938.4]
  input         io_memStreams_stores_0_data_valid, // @[:@153938.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@153938.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@153938.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@153938.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@153938.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@153938.4]
  input         io_dram_0_cmd_ready, // @[:@153938.4]
  output        io_dram_0_cmd_valid, // @[:@153938.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@153938.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@153938.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@153938.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@153938.4]
  input         io_dram_0_wdata_ready, // @[:@153938.4]
  output        io_dram_0_wdata_valid, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@153938.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@153938.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@153938.4]
  output        io_dram_0_rresp_ready, // @[:@153938.4]
  output        io_dram_0_wresp_ready, // @[:@153938.4]
  input         io_dram_0_wresp_valid, // @[:@153938.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@153938.4]
  input         io_dram_1_cmd_ready, // @[:@153938.4]
  output        io_dram_1_cmd_valid, // @[:@153938.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@153938.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@153938.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@153938.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@153938.4]
  input         io_dram_1_wdata_ready, // @[:@153938.4]
  output        io_dram_1_wdata_valid, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@153938.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@153938.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@153938.4]
  output        io_dram_1_rresp_ready, // @[:@153938.4]
  output        io_dram_1_wresp_ready, // @[:@153938.4]
  input         io_dram_1_wresp_valid, // @[:@153938.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@153938.4]
  input         io_dram_2_cmd_ready, // @[:@153938.4]
  output        io_dram_2_cmd_valid, // @[:@153938.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@153938.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@153938.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@153938.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@153938.4]
  input         io_dram_2_wdata_ready, // @[:@153938.4]
  output        io_dram_2_wdata_valid, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@153938.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@153938.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@153938.4]
  output        io_dram_2_rresp_ready, // @[:@153938.4]
  output        io_dram_2_wresp_ready, // @[:@153938.4]
  input         io_dram_2_wresp_valid, // @[:@153938.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@153938.4]
  input         io_dram_3_cmd_ready, // @[:@153938.4]
  output        io_dram_3_cmd_valid, // @[:@153938.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@153938.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@153938.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@153938.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@153938.4]
  input         io_dram_3_wdata_ready, // @[:@153938.4]
  output        io_dram_3_wdata_valid, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@153938.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@153938.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@153938.4]
  output        io_dram_3_rresp_ready, // @[:@153938.4]
  output        io_dram_3_wresp_ready, // @[:@153938.4]
  input         io_dram_3_wresp_valid, // @[:@153938.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@153938.4]
  input         io_heap_0_req_valid, // @[:@153938.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@153938.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@153938.4]
  output        io_heap_0_resp_valid, // @[:@153938.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@153938.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@153938.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@153944.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@153944.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@153944.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@153944.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@154937.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@154937.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@154937.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@155897.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@155897.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@155897.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@156857.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@156857.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@156857.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@156857.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@157817.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@157817.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@157817.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@157817.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@157817.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@157817.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@157817.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@157817.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@157817.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@157817.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@157817.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@157817.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@157826.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@157826.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@157826.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@157826.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@157826.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@157826.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@157826.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@157826.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@157826.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@159876.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@159876.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@159876.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@159876.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@159895.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@159895.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@159895.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@159895.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@159895.4]
  wire [63:0] _T_1020; // @[:@159853.4 :@159854.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@159855.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@159857.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@159859.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@159861.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@159863.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@159865.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@159867.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@159903.4]
  reg  _T_1047; // @[package.scala 152:20:@159906.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@159908.4]
  wire  _T_1049; // @[package.scala 153:8:@159909.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@159913.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@159914.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@159917.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@159918.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@159920.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@159921.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@159923.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@159926.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@159905.4 Fringe.scala 163:24:@159924.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@159905.4 Fringe.scala 162:28:@159922.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@159927.4]
  wire  alloc; // @[Fringe.scala 202:38:@161557.4]
  wire  dealloc; // @[Fringe.scala 203:40:@161558.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@161559.4]
  reg  _T_1572; // @[package.scala 152:20:@161560.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@161562.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@153944.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@154937.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@155897.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@156857.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@157817.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@157826.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@159876.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@159895.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@159853.4 :@159854.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@159855.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@159857.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@159859.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@159861.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@159863.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@159865.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@159867.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@159903.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@159908.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@159909.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@159913.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@159914.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@159917.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@159918.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@159920.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@159921.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@159923.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@159926.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@159905.4 Fringe.scala 163:24:@159924.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@159905.4 Fringe.scala 162:28:@159922.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@159927.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@161557.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@161558.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@161559.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@161562.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@159851.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@159871.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@159872.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@159893.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@159894.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@154863.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@154859.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@154854.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@154853.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@161055.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@161054.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@161053.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@161051.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@161050.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@161048.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@161032.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@161033.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@161034.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@161035.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@161036.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@161037.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@161038.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@161039.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@161040.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@161041.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@161042.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@161043.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@161044.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@161045.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@161046.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@161047.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@160968.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@160969.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@160970.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@160971.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@160972.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@160973.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@160974.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@160975.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@160976.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@160977.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@160978.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@160979.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@160980.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@160981.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@160982.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@160983.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@160984.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@160985.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@160986.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@160987.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@160988.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@160989.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@160990.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@160991.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@160992.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@160993.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@160994.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@160995.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@160996.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@160997.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@160998.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@160999.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@161000.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@161001.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@161002.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@161003.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@161004.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@161005.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@161006.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@161007.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@161008.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@161009.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@161010.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@161011.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@161012.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@161013.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@161014.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@161015.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@161016.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@161017.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@161018.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@161019.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@161020.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@161021.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@161022.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@161023.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@161024.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@161025.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@161026.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@161027.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@161028.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@161029.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@161030.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@161031.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@160967.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@160966.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@160947.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@161167.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@161166.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@161165.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@161163.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@161162.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@161160.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@161144.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@161145.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@161146.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@161147.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@161148.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@161149.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@161150.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@161151.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@161152.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@161153.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@161154.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@161155.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@161156.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@161157.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@161158.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@161159.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@161080.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@161081.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@161082.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@161083.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@161084.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@161085.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@161086.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@161087.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@161088.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@161089.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@161090.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@161091.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@161092.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@161093.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@161094.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@161095.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@161096.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@161097.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@161098.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@161099.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@161100.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@161101.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@161102.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@161103.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@161104.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@161105.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@161106.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@161107.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@161108.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@161109.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@161110.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@161111.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@161112.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@161113.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@161114.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@161115.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@161116.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@161117.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@161118.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@161119.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@161120.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@161121.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@161122.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@161123.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@161124.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@161125.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@161126.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@161127.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@161128.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@161129.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@161130.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@161131.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@161132.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@161133.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@161134.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@161135.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@161136.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@161137.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@161138.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@161139.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@161140.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@161141.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@161142.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@161143.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@161079.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@161078.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@161059.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@161279.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@161278.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@161277.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@161275.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@161274.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@161272.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@161256.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@161257.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@161258.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@161259.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@161260.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@161261.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@161262.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@161263.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@161264.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@161265.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@161266.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@161267.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@161268.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@161269.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@161270.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@161271.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@161192.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@161193.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@161194.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@161195.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@161196.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@161197.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@161198.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@161199.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@161200.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@161201.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@161202.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@161203.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@161204.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@161205.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@161206.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@161207.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@161208.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@161209.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@161210.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@161211.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@161212.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@161213.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@161214.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@161215.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@161216.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@161217.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@161218.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@161219.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@161220.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@161221.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@161222.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@161223.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@161224.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@161225.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@161226.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@161227.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@161228.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@161229.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@161230.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@161231.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@161232.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@161233.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@161234.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@161235.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@161236.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@161237.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@161238.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@161239.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@161240.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@161241.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@161242.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@161243.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@161244.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@161245.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@161246.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@161247.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@161248.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@161249.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@161250.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@161251.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@161252.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@161253.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@161254.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@161255.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@161191.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@161190.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@161171.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@161391.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@161390.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@161389.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@161387.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@161386.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@161384.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@161368.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@161369.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@161370.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@161371.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@161372.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@161373.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@161374.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@161375.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@161376.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@161377.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@161378.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@161379.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@161380.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@161381.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@161382.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@161383.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@161304.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@161305.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@161306.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@161307.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@161308.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@161309.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@161310.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@161311.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@161312.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@161313.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@161314.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@161315.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@161316.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@161317.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@161318.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@161319.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@161320.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@161321.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@161322.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@161323.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@161324.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@161325.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@161326.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@161327.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@161328.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@161329.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@161330.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@161331.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@161332.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@161333.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@161334.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@161335.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@161336.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@161337.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@161338.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@161339.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@161340.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@161341.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@161342.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@161343.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@161344.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@161345.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@161346.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@161347.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@161348.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@161349.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@161350.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@161351.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@161352.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@161353.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@161354.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@161355.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@161356.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@161357.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@161358.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@161359.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@161360.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@161361.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@161362.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@161363.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@161364.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@161365.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@161366.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@161367.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@161303.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@161302.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@161283.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@157822.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@157821.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@157820.4]
  assign dramArbs_0_clock = clock; // @[:@153945.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@153946.4 Fringe.scala 187:30:@160937.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@160941.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@154862.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@154861.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@154860.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@154858.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@154857.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@154856.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@154855.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@161056.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@161049.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@160946.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@160945.4]
  assign dramArbs_1_clock = clock; // @[:@154938.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@154939.4 Fringe.scala 187:30:@160938.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@160942.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@161168.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@161161.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@161058.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@161057.4]
  assign dramArbs_2_clock = clock; // @[:@155898.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@155899.4 Fringe.scala 187:30:@160939.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@160943.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@161280.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@161273.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@161170.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@161169.4]
  assign dramArbs_3_clock = clock; // @[:@156858.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@156859.4 Fringe.scala 187:30:@160940.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@160944.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@161392.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@161385.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@161282.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@161281.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@157825.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@157824.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@157823.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@161564.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@161565.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@161566.4]
  assign regs_clock = clock; // @[:@157827.4]
  assign regs_reset = reset; // @[:@157828.4 Fringe.scala 139:14:@159875.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@159847.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@159849.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@159848.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@159850.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@159873.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@159925.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@159929.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@159932.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@159931.4]
  assign timeoutCtr_clock = clock; // @[:@159877.4]
  assign timeoutCtr_reset = reset; // @[:@159878.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@159892.4]
  assign depulser_clock = clock; // @[:@159896.4]
  assign depulser_reset = reset; // @[:@159897.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@159902.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@159904.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@161581.2]
  input         clock, // @[:@161582.4]
  input         reset, // @[:@161583.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@161584.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@161584.4]
  input         io_S_AXI_AWVALID, // @[:@161584.4]
  output        io_S_AXI_AWREADY, // @[:@161584.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@161584.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@161584.4]
  input         io_S_AXI_ARVALID, // @[:@161584.4]
  output        io_S_AXI_ARREADY, // @[:@161584.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@161584.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@161584.4]
  input         io_S_AXI_WVALID, // @[:@161584.4]
  output        io_S_AXI_WREADY, // @[:@161584.4]
  output [31:0] io_S_AXI_RDATA, // @[:@161584.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@161584.4]
  output        io_S_AXI_RVALID, // @[:@161584.4]
  input         io_S_AXI_RREADY, // @[:@161584.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@161584.4]
  output        io_S_AXI_BVALID, // @[:@161584.4]
  input         io_S_AXI_BREADY, // @[:@161584.4]
  output [31:0] io_raddr, // @[:@161584.4]
  output        io_wen, // @[:@161584.4]
  output [31:0] io_waddr, // @[:@161584.4]
  output [31:0] io_wdata, // @[:@161584.4]
  input  [31:0] io_rdata // @[:@161584.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@161586.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@161610.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@161606.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@161602.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@161601.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@161600.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@161599.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@161597.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@161596.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@161618.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@161621.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@161619.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@161620.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@161622.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@161617.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@161614.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@161613.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@161612.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@161611.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@161609.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@161608.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@161607.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@161605.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@161604.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@161603.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@161598.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@161595.4]
endmodule
module MAGToAXI4Bridge( // @[:@161624.2]
  output         io_in_cmd_ready, // @[:@161627.4]
  input          io_in_cmd_valid, // @[:@161627.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@161627.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@161627.4]
  input          io_in_cmd_bits_isWr, // @[:@161627.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@161627.4]
  output         io_in_wdata_ready, // @[:@161627.4]
  input          io_in_wdata_valid, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@161627.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@161627.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@161627.4]
  input          io_in_wdata_bits_wlast, // @[:@161627.4]
  input          io_in_rresp_ready, // @[:@161627.4]
  input          io_in_wresp_ready, // @[:@161627.4]
  output         io_in_wresp_valid, // @[:@161627.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@161627.4]
  output [31:0]  io_M_AXI_AWID, // @[:@161627.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@161627.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@161627.4]
  output         io_M_AXI_AWVALID, // @[:@161627.4]
  input          io_M_AXI_AWREADY, // @[:@161627.4]
  output [31:0]  io_M_AXI_ARID, // @[:@161627.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@161627.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@161627.4]
  output         io_M_AXI_ARVALID, // @[:@161627.4]
  input          io_M_AXI_ARREADY, // @[:@161627.4]
  output [511:0] io_M_AXI_WDATA, // @[:@161627.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@161627.4]
  output         io_M_AXI_WLAST, // @[:@161627.4]
  output         io_M_AXI_WVALID, // @[:@161627.4]
  input          io_M_AXI_WREADY, // @[:@161627.4]
  output         io_M_AXI_RREADY, // @[:@161627.4]
  input  [31:0]  io_M_AXI_BID, // @[:@161627.4]
  input          io_M_AXI_BVALID, // @[:@161627.4]
  output         io_M_AXI_BREADY // @[:@161627.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@161784.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@161785.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@161786.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@161794.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@161821.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@161826.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@161837.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@161846.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@161855.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@161864.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@161873.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@161882.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@161890.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@161784.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@161785.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@161786.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@161794.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@161821.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@161826.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@161837.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@161846.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@161855.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@161864.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@161873.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@161882.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@161890.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@161798.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@161895.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@161948.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@161950.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@161799.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@161800.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@161804.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@161812.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@161782.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@161783.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@161787.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@161796.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@161828.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@161892.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@161893.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@161894.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@161945.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@161946.4]
endmodule
module FringeZynq( // @[:@162936.2]
  input          clock, // @[:@162937.4]
  input          reset, // @[:@162938.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@162939.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@162939.4]
  input          io_S_AXI_AWVALID, // @[:@162939.4]
  output         io_S_AXI_AWREADY, // @[:@162939.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@162939.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@162939.4]
  input          io_S_AXI_ARVALID, // @[:@162939.4]
  output         io_S_AXI_ARREADY, // @[:@162939.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@162939.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@162939.4]
  input          io_S_AXI_WVALID, // @[:@162939.4]
  output         io_S_AXI_WREADY, // @[:@162939.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@162939.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@162939.4]
  output         io_S_AXI_RVALID, // @[:@162939.4]
  input          io_S_AXI_RREADY, // @[:@162939.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@162939.4]
  output         io_S_AXI_BVALID, // @[:@162939.4]
  input          io_S_AXI_BREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@162939.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@162939.4]
  output         io_M_AXI_0_AWVALID, // @[:@162939.4]
  input          io_M_AXI_0_AWREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@162939.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@162939.4]
  output         io_M_AXI_0_ARVALID, // @[:@162939.4]
  input          io_M_AXI_0_ARREADY, // @[:@162939.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@162939.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@162939.4]
  output         io_M_AXI_0_WLAST, // @[:@162939.4]
  output         io_M_AXI_0_WVALID, // @[:@162939.4]
  input          io_M_AXI_0_WREADY, // @[:@162939.4]
  output         io_M_AXI_0_RREADY, // @[:@162939.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@162939.4]
  input          io_M_AXI_0_BVALID, // @[:@162939.4]
  output         io_M_AXI_0_BREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@162939.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@162939.4]
  output         io_M_AXI_1_AWVALID, // @[:@162939.4]
  input          io_M_AXI_1_AWREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@162939.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@162939.4]
  output         io_M_AXI_1_ARVALID, // @[:@162939.4]
  input          io_M_AXI_1_ARREADY, // @[:@162939.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@162939.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@162939.4]
  output         io_M_AXI_1_WLAST, // @[:@162939.4]
  output         io_M_AXI_1_WVALID, // @[:@162939.4]
  input          io_M_AXI_1_WREADY, // @[:@162939.4]
  output         io_M_AXI_1_RREADY, // @[:@162939.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@162939.4]
  input          io_M_AXI_1_BVALID, // @[:@162939.4]
  output         io_M_AXI_1_BREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@162939.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@162939.4]
  output         io_M_AXI_2_AWVALID, // @[:@162939.4]
  input          io_M_AXI_2_AWREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@162939.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@162939.4]
  output         io_M_AXI_2_ARVALID, // @[:@162939.4]
  input          io_M_AXI_2_ARREADY, // @[:@162939.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@162939.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@162939.4]
  output         io_M_AXI_2_WLAST, // @[:@162939.4]
  output         io_M_AXI_2_WVALID, // @[:@162939.4]
  input          io_M_AXI_2_WREADY, // @[:@162939.4]
  output         io_M_AXI_2_RREADY, // @[:@162939.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@162939.4]
  input          io_M_AXI_2_BVALID, // @[:@162939.4]
  output         io_M_AXI_2_BREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@162939.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@162939.4]
  output         io_M_AXI_3_AWVALID, // @[:@162939.4]
  input          io_M_AXI_3_AWREADY, // @[:@162939.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@162939.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@162939.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@162939.4]
  output         io_M_AXI_3_ARVALID, // @[:@162939.4]
  input          io_M_AXI_3_ARREADY, // @[:@162939.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@162939.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@162939.4]
  output         io_M_AXI_3_WLAST, // @[:@162939.4]
  output         io_M_AXI_3_WVALID, // @[:@162939.4]
  input          io_M_AXI_3_WREADY, // @[:@162939.4]
  output         io_M_AXI_3_RREADY, // @[:@162939.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@162939.4]
  input          io_M_AXI_3_BVALID, // @[:@162939.4]
  output         io_M_AXI_3_BREADY, // @[:@162939.4]
  output         io_enable, // @[:@162939.4]
  input          io_done, // @[:@162939.4]
  output         io_reset, // @[:@162939.4]
  output [63:0]  io_argIns_0, // @[:@162939.4]
  output [63:0]  io_argIns_1, // @[:@162939.4]
  input          io_argOuts_0_valid, // @[:@162939.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@162939.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@162939.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@162939.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@162939.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@162939.4]
  output         io_memStreams_stores_0_data_ready, // @[:@162939.4]
  input          io_memStreams_stores_0_data_valid, // @[:@162939.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@162939.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@162939.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@162939.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@162939.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@162939.4]
  input          io_heap_0_req_valid, // @[:@162939.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@162939.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@162939.4]
  output         io_heap_0_resp_valid, // @[:@162939.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@162939.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@162939.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@163410.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@163410.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@163410.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@164316.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@164316.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@164316.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@164316.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@164316.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@164316.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@164316.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@164316.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@164466.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@164466.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@164466.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@164466.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@164466.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@164466.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@164466.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@164622.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@164622.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@164622.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@164622.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@164622.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@164622.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@164622.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@164778.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@164778.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@164778.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@164778.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@164778.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@164778.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@164778.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@164934.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@164934.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@164934.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@164934.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@164934.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@164934.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@164934.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@164934.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@163410.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@164316.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@164466.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@164622.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@164778.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@164934.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@164334.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@164330.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@164326.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@164325.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@164324.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@164323.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@164321.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@164320.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@164621.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@164619.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@164618.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@164611.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@164609.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@164607.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@164606.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@164599.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@164597.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@164596.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@164595.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@164594.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@164586.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@164581.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@164777.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@164775.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@164774.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@164767.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@164765.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@164763.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@164762.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@164755.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@164753.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@164752.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@164751.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@164750.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@164742.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@164737.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@164933.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@164931.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@164930.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@164923.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@164921.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@164919.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@164918.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@164911.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@164909.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@164908.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@164907.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@164906.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@164898.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@164893.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@165089.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@165087.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@165086.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@165079.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@165077.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@165075.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@165074.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@165067.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@165065.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@165064.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@165063.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@165062.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@165054.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@165049.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@164344.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@164348.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@164349.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@164350.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@164437.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@164433.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@164428.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@164427.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@164462.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@164461.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@164460.4]
  assign fringeCommon_clock = clock; // @[:@163411.4]
  assign fringeCommon_reset = reset; // @[:@163412.4 FringeZynq.scala 117:22:@164347.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@164338.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@164339.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@164340.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@164341.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@164345.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@164352.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@164351.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@164436.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@164435.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@164434.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@164432.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@164431.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@164430.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@164429.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@164580.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@164573.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@164470.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@164469.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@164736.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@164729.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@164626.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@164625.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@164892.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@164885.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@164782.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@164781.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@165048.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@165041.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@164938.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@164937.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@164465.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@164464.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@164463.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@164317.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@164318.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@164337.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@164336.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@164335.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@164333.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@164332.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@164331.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@164329.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@164328.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@164327.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@164322.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@164319.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@164342.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@164579.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@164578.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@164577.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@164575.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@164574.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@164572.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@164556.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@164557.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@164558.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@164559.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@164560.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@164561.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@164562.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@164563.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@164564.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@164565.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@164566.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@164567.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@164568.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@164569.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@164570.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@164571.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@164492.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@164493.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@164494.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@164495.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@164496.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@164497.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@164498.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@164499.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@164500.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@164501.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@164502.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@164503.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@164504.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@164505.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@164506.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@164507.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@164508.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@164509.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@164510.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@164511.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@164512.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@164513.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@164514.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@164515.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@164516.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@164517.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@164518.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@164519.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@164520.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@164521.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@164522.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@164523.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@164524.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@164525.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@164526.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@164527.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@164528.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@164529.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@164530.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@164531.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@164532.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@164533.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@164534.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@164535.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@164536.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@164537.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@164538.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@164539.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@164540.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@164541.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@164542.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@164543.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@164544.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@164545.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@164546.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@164547.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@164548.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@164549.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@164550.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@164551.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@164552.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@164553.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@164554.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@164555.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@164491.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@164490.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@164471.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@164610.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@164598.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@164593.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@164585.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@164582.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@164735.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@164734.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@164733.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@164731.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@164730.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@164728.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@164712.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@164713.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@164714.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@164715.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@164716.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@164717.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@164718.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@164719.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@164720.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@164721.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@164722.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@164723.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@164724.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@164725.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@164726.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@164727.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@164648.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@164649.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@164650.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@164651.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@164652.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@164653.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@164654.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@164655.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@164656.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@164657.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@164658.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@164659.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@164660.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@164661.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@164662.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@164663.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@164664.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@164665.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@164666.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@164667.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@164668.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@164669.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@164670.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@164671.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@164672.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@164673.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@164674.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@164675.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@164676.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@164677.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@164678.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@164679.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@164680.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@164681.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@164682.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@164683.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@164684.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@164685.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@164686.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@164687.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@164688.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@164689.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@164690.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@164691.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@164692.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@164693.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@164694.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@164695.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@164696.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@164697.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@164698.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@164699.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@164700.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@164701.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@164702.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@164703.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@164704.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@164705.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@164706.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@164707.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@164708.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@164709.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@164710.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@164711.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@164647.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@164646.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@164627.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@164766.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@164754.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@164749.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@164741.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@164738.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@164891.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@164890.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@164889.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@164887.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@164886.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@164884.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@164868.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@164869.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@164870.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@164871.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@164872.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@164873.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@164874.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@164875.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@164876.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@164877.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@164878.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@164879.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@164880.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@164881.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@164882.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@164883.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@164804.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@164805.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@164806.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@164807.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@164808.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@164809.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@164810.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@164811.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@164812.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@164813.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@164814.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@164815.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@164816.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@164817.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@164818.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@164819.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@164820.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@164821.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@164822.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@164823.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@164824.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@164825.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@164826.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@164827.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@164828.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@164829.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@164830.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@164831.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@164832.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@164833.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@164834.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@164835.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@164836.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@164837.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@164838.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@164839.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@164840.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@164841.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@164842.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@164843.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@164844.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@164845.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@164846.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@164847.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@164848.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@164849.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@164850.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@164851.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@164852.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@164853.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@164854.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@164855.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@164856.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@164857.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@164858.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@164859.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@164860.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@164861.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@164862.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@164863.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@164864.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@164865.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@164866.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@164867.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@164803.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@164802.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@164783.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@164922.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@164910.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@164905.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@164897.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@164894.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@165047.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@165046.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@165045.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@165043.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@165042.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@165040.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@165024.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@165025.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@165026.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@165027.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@165028.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@165029.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@165030.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@165031.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@165032.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@165033.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@165034.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@165035.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@165036.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@165037.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@165038.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@165039.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@164960.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@164961.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@164962.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@164963.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@164964.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@164965.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@164966.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@164967.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@164968.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@164969.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@164970.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@164971.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@164972.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@164973.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@164974.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@164975.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@164976.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@164977.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@164978.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@164979.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@164980.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@164981.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@164982.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@164983.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@164984.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@164985.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@164986.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@164987.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@164988.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@164989.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@164990.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@164991.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@164992.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@164993.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@164994.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@164995.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@164996.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@164997.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@164998.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@164999.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@165000.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@165001.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@165002.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@165003.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@165004.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@165005.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@165006.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@165007.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@165008.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@165009.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@165010.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@165011.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@165012.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@165013.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@165014.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@165015.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@165016.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@165017.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@165018.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@165019.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@165020.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@165021.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@165022.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@165023.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@164959.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@164958.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@164939.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@165078.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@165066.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@165061.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@165053.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@165050.4]
endmodule
module SpatialIP( // @[:@165091.2]
  input          clock, // @[:@165092.4]
  input          reset, // @[:@165093.4]
  input          io_raddr, // @[:@165094.4]
  input          io_wen, // @[:@165094.4]
  input          io_waddr, // @[:@165094.4]
  input          io_wdata, // @[:@165094.4]
  output         io_rdata, // @[:@165094.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@165094.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@165094.4]
  input          io_S_AXI_AWVALID, // @[:@165094.4]
  output         io_S_AXI_AWREADY, // @[:@165094.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@165094.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@165094.4]
  input          io_S_AXI_ARVALID, // @[:@165094.4]
  output         io_S_AXI_ARREADY, // @[:@165094.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@165094.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@165094.4]
  input          io_S_AXI_WVALID, // @[:@165094.4]
  output         io_S_AXI_WREADY, // @[:@165094.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@165094.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@165094.4]
  output         io_S_AXI_RVALID, // @[:@165094.4]
  input          io_S_AXI_RREADY, // @[:@165094.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@165094.4]
  output         io_S_AXI_BVALID, // @[:@165094.4]
  input          io_S_AXI_BREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@165094.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@165094.4]
  output         io_M_AXI_0_AWLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@165094.4]
  output         io_M_AXI_0_AWVALID, // @[:@165094.4]
  input          io_M_AXI_0_AWREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@165094.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@165094.4]
  output         io_M_AXI_0_ARLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@165094.4]
  output         io_M_AXI_0_ARVALID, // @[:@165094.4]
  input          io_M_AXI_0_ARREADY, // @[:@165094.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@165094.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@165094.4]
  output         io_M_AXI_0_WLAST, // @[:@165094.4]
  output         io_M_AXI_0_WVALID, // @[:@165094.4]
  input          io_M_AXI_0_WREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@165094.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@165094.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@165094.4]
  input          io_M_AXI_0_RLAST, // @[:@165094.4]
  input          io_M_AXI_0_RVALID, // @[:@165094.4]
  output         io_M_AXI_0_RREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@165094.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@165094.4]
  input          io_M_AXI_0_BVALID, // @[:@165094.4]
  output         io_M_AXI_0_BREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@165094.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@165094.4]
  output         io_M_AXI_1_AWLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@165094.4]
  output         io_M_AXI_1_AWVALID, // @[:@165094.4]
  input          io_M_AXI_1_AWREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@165094.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@165094.4]
  output         io_M_AXI_1_ARLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@165094.4]
  output         io_M_AXI_1_ARVALID, // @[:@165094.4]
  input          io_M_AXI_1_ARREADY, // @[:@165094.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@165094.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@165094.4]
  output         io_M_AXI_1_WLAST, // @[:@165094.4]
  output         io_M_AXI_1_WVALID, // @[:@165094.4]
  input          io_M_AXI_1_WREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@165094.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@165094.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@165094.4]
  input          io_M_AXI_1_RLAST, // @[:@165094.4]
  input          io_M_AXI_1_RVALID, // @[:@165094.4]
  output         io_M_AXI_1_RREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@165094.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@165094.4]
  input          io_M_AXI_1_BVALID, // @[:@165094.4]
  output         io_M_AXI_1_BREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@165094.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@165094.4]
  output         io_M_AXI_2_AWLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@165094.4]
  output         io_M_AXI_2_AWVALID, // @[:@165094.4]
  input          io_M_AXI_2_AWREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@165094.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@165094.4]
  output         io_M_AXI_2_ARLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@165094.4]
  output         io_M_AXI_2_ARVALID, // @[:@165094.4]
  input          io_M_AXI_2_ARREADY, // @[:@165094.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@165094.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@165094.4]
  output         io_M_AXI_2_WLAST, // @[:@165094.4]
  output         io_M_AXI_2_WVALID, // @[:@165094.4]
  input          io_M_AXI_2_WREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@165094.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@165094.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@165094.4]
  input          io_M_AXI_2_RLAST, // @[:@165094.4]
  input          io_M_AXI_2_RVALID, // @[:@165094.4]
  output         io_M_AXI_2_RREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@165094.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@165094.4]
  input          io_M_AXI_2_BVALID, // @[:@165094.4]
  output         io_M_AXI_2_BREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@165094.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@165094.4]
  output         io_M_AXI_3_AWLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@165094.4]
  output         io_M_AXI_3_AWVALID, // @[:@165094.4]
  input          io_M_AXI_3_AWREADY, // @[:@165094.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@165094.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@165094.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@165094.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@165094.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@165094.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@165094.4]
  output         io_M_AXI_3_ARLOCK, // @[:@165094.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@165094.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@165094.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@165094.4]
  output         io_M_AXI_3_ARVALID, // @[:@165094.4]
  input          io_M_AXI_3_ARREADY, // @[:@165094.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@165094.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@165094.4]
  output         io_M_AXI_3_WLAST, // @[:@165094.4]
  output         io_M_AXI_3_WVALID, // @[:@165094.4]
  input          io_M_AXI_3_WREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@165094.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@165094.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@165094.4]
  input          io_M_AXI_3_RLAST, // @[:@165094.4]
  input          io_M_AXI_3_RVALID, // @[:@165094.4]
  output         io_M_AXI_3_RREADY, // @[:@165094.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@165094.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@165094.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@165094.4]
  input          io_M_AXI_3_BVALID, // @[:@165094.4]
  output         io_M_AXI_3_BREADY, // @[:@165094.4]
  input          io_TOP_AXI_AWID, // @[:@165094.4]
  input          io_TOP_AXI_AWUSER, // @[:@165094.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@165094.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@165094.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@165094.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@165094.4]
  input          io_TOP_AXI_AWLOCK, // @[:@165094.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@165094.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@165094.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@165094.4]
  input          io_TOP_AXI_AWVALID, // @[:@165094.4]
  input          io_TOP_AXI_AWREADY, // @[:@165094.4]
  input          io_TOP_AXI_ARID, // @[:@165094.4]
  input          io_TOP_AXI_ARUSER, // @[:@165094.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@165094.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@165094.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@165094.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@165094.4]
  input          io_TOP_AXI_ARLOCK, // @[:@165094.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@165094.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@165094.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@165094.4]
  input          io_TOP_AXI_ARVALID, // @[:@165094.4]
  input          io_TOP_AXI_ARREADY, // @[:@165094.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@165094.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@165094.4]
  input          io_TOP_AXI_WLAST, // @[:@165094.4]
  input          io_TOP_AXI_WVALID, // @[:@165094.4]
  input          io_TOP_AXI_WREADY, // @[:@165094.4]
  input          io_TOP_AXI_RID, // @[:@165094.4]
  input          io_TOP_AXI_RUSER, // @[:@165094.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@165094.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@165094.4]
  input          io_TOP_AXI_RLAST, // @[:@165094.4]
  input          io_TOP_AXI_RVALID, // @[:@165094.4]
  input          io_TOP_AXI_RREADY, // @[:@165094.4]
  input          io_TOP_AXI_BID, // @[:@165094.4]
  input          io_TOP_AXI_BUSER, // @[:@165094.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@165094.4]
  input          io_TOP_AXI_BVALID, // @[:@165094.4]
  input          io_TOP_AXI_BREADY, // @[:@165094.4]
  input          io_DWIDTH_AXI_AWID, // @[:@165094.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@165094.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@165094.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@165094.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@165094.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@165094.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@165094.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@165094.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@165094.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@165094.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@165094.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@165094.4]
  input          io_DWIDTH_AXI_ARID, // @[:@165094.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@165094.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@165094.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@165094.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@165094.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@165094.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@165094.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@165094.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@165094.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@165094.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@165094.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@165094.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@165094.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@165094.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@165094.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@165094.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@165094.4]
  input          io_DWIDTH_AXI_RID, // @[:@165094.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@165094.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@165094.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@165094.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@165094.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@165094.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@165094.4]
  input          io_DWIDTH_AXI_BID, // @[:@165094.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@165094.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@165094.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@165094.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@165094.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@165094.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@165094.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@165094.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@165094.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@165094.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@165094.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@165094.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@165094.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@165094.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@165094.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@165094.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@165094.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@165094.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@165094.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@165094.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@165094.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@165094.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@165094.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@165094.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@165094.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@165094.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@165094.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@165094.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@165094.4]
  input          io_PROTOCOL_AXI_RID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@165094.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@165094.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@165094.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@165094.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@165094.4]
  input          io_PROTOCOL_AXI_BID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@165094.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@165094.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@165094.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@165094.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@165094.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@165094.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@165094.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@165094.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@165094.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@165094.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@165094.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@165094.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@165094.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@165094.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@165094.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@165094.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@165094.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@165094.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@165094.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@165094.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@165094.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@165094.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@165094.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@165094.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@165096.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@165096.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@165096.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@165096.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@165096.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@165096.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@165096.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@165096.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@165096.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@165096.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@165238.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@165238.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@165238.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@165238.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@165238.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@165238.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@165238.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@165096.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@165238.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@165256.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@165252.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@165248.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@165247.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@165246.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@165245.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@165243.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@165242.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@165300.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@165299.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@165298.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@165297.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@165296.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@165295.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@165294.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@165293.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@165292.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@165291.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@165290.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@165288.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@165287.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@165286.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@165285.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@165284.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@165283.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@165282.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@165281.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@165280.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@165279.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@165278.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@165276.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@165275.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@165274.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@165273.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@165265.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@165260.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@165341.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@165340.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@165339.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@165338.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@165337.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@165336.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@165335.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@165334.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@165333.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@165332.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@165331.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@165329.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@165328.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@165327.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@165326.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@165325.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@165324.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@165323.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@165322.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@165321.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@165320.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@165319.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@165317.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@165316.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@165315.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@165314.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@165306.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@165301.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@165382.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@165381.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@165380.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@165379.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@165378.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@165377.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@165376.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@165375.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@165374.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@165373.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@165372.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@165370.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@165369.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@165368.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@165367.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@165366.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@165365.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@165364.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@165363.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@165362.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@165361.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@165360.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@165358.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@165357.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@165356.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@165355.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@165347.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@165342.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@165423.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@165422.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@165421.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@165420.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@165419.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@165418.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@165417.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@165416.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@165415.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@165414.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@165413.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@165411.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@165410.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@165409.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@165408.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@165407.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@165406.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@165405.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@165404.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@165403.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@165402.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@165401.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@165399.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@165398.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@165397.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@165396.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@165388.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@165383.4]
  assign accel_clock = clock; // @[:@165097.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@165098.4 Zynq.scala 54:17:@165712.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@165707.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@165700.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@165695.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@165679.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@165680.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@165681.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@165682.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@165683.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@165684.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@165685.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@165686.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@165687.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@165688.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@165689.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@165690.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@165691.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@165692.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@165693.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@165694.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@165678.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@165674.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@165669.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@165668.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@165667.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@165648.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@165632.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@165633.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@165634.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@165635.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@165636.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@165637.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@165638.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@165639.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@165640.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@165641.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@165642.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@165643.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@165644.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@165645.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@165646.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@165647.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@165631.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@165596.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@165595.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@165703.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@165702.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@165701.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@165589.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@165590.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@165593.4]
  assign FringeZynq_clock = clock; // @[:@165239.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@165240.4 Zynq.scala 53:18:@165711.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@165259.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@165258.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@165257.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@165255.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@165254.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@165253.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@165251.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@165250.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@165249.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@165244.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@165241.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@165289.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@165277.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@165272.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@165264.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@165261.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@165330.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@165318.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@165313.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@165305.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@165302.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@165371.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@165359.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@165354.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@165346.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@165343.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@165412.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@165400.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@165395.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@165387.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@165384.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@165708.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@165592.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@165591.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@165677.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@165676.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@165675.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@165673.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@165672.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@165671.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@165670.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@165706.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@165705.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@165704.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




