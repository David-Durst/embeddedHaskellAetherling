module FIFO(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7
);
  reg [15:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [15:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [15:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [15:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [15:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [15:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [15:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [15:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_8;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCounters_1(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters_1 NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input         clock,
  input         RE,
  input  [7:0]  RADDR,
  output [15:0] RDATA_0,
  output [15:0] RDATA_1,
  output [15:0] RDATA_2,
  output [15:0] RDATA_3,
  output [15:0] RDATA_4,
  output [15:0] RDATA_5,
  output [15:0] RDATA_6,
  output [15:0] RDATA_7,
  input         WE,
  input  [7:0]  WADDR,
  input  [15:0] WDATA_0,
  input  [15:0] WDATA_1,
  input  [15:0] WDATA_2,
  input  [15:0] WDATA_3,
  input  [15:0] WDATA_4,
  input  [15:0] WDATA_5,
  input  [15:0] WDATA_6,
  input  [15:0] WDATA_7
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [127:0] ram [0:239]; // @[RAM_ST.scala 29:24]
  reg [127:0] _RAND_0;
  wire [127:0] ram__T_15_data; // @[RAM_ST.scala 29:24]
  wire [7:0] ram__T_15_addr; // @[RAM_ST.scala 29:24]
  reg [127:0] _RAND_1;
  wire [127:0] ram__T_9_data; // @[RAM_ST.scala 29:24]
  wire [7:0] ram__T_9_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_9_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_9_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [7:0] ram__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [7:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_120; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_121; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_122; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_123; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_124; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_125; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_126; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_127; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_128; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_129; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_130; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_131; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_132; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_133; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_134; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_135; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_136; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_137; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_138; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_139; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_140; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_141; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_142; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_143; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_144; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_145; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_146; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_147; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_148; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_149; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_150; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_151; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_152; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_153; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_154; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_155; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_156; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_157; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_158; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_159; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_160; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_161; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_162; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_163; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_164; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_165; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_166; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_167; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_168; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_169; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_170; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_171; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_172; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_173; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_174; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_175; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_176; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_177; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_178; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_179; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_180; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_181; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_182; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_183; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_184; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_185; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_186; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_187; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_188; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_189; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_190; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_191; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_192; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_193; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_194; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_195; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_196; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_197; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_198; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_199; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_200; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_201; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_202; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_203; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_204; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_205; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_206; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_207; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_208; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_209; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_210; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_211; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_212; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_213; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_214; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_215; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_216; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_217; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_218; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_219; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_220; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_221; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_222; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_223; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_224; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_225; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_226; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_227; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_228; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_229; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_230; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_231; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_232; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_233; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_234; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_235; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_236; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_237; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_238; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_239; // @[RAM_ST.scala 31:71]
  wire [8:0] _T; // @[RAM_ST.scala 31:71]
  wire [63:0] _T_4; // @[RAM_ST.scala 31:115]
  wire [63:0] _T_7; // @[RAM_ST.scala 31:115]
  wire [7:0] _GEN_246; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_247; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_248; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_249; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_250; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_251; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_252; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_253; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_254; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_255; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_256; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_257; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_258; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_259; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_260; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_261; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_262; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_263; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_264; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_265; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_266; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_267; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_268; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_269; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_270; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_271; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_272; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_273; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_274; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_275; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_276; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_277; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_278; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_279; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_280; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_281; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_282; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_283; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_284; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_285; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_286; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_287; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_288; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_289; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_290; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_291; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_292; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_293; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_294; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_295; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_296; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_297; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_298; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_299; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_300; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_301; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_302; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_303; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_304; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_305; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_306; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_307; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_308; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_309; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_310; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_311; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_312; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_313; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_314; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_315; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_316; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_317; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_318; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_319; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_320; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_321; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_322; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_323; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_324; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_325; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_326; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_327; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_328; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_329; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_330; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_331; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_332; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_333; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_334; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_335; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_336; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_337; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_338; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_339; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_340; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_341; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_342; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_343; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_344; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_345; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_346; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_347; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_348; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_349; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_350; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_351; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_352; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_353; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_354; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_355; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_356; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_357; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_358; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_359; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_360; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_361; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_362; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_363; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_364; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_365; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_366; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_367; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_368; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_369; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_370; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_371; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_372; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_373; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_374; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_375; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_376; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_377; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_378; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_379; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_380; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_381; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_382; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_383; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_384; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_385; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_386; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_387; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_388; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_389; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_390; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_391; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_392; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_393; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_394; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_395; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_396; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_397; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_398; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_399; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_400; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_401; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_402; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_403; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_404; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_405; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_406; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_407; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_408; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_409; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_410; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_411; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_412; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_413; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_414; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_415; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_416; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_417; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_418; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_419; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_420; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_421; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_422; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_423; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_424; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_425; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_426; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_427; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_428; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_429; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_430; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_431; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_432; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_433; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_434; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_435; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_436; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_437; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_438; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_439; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_440; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_441; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_442; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_443; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_444; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_445; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_446; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_447; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_448; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_449; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_450; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_451; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_452; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_453; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_454; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_455; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_456; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_457; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_458; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_459; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_460; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_461; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_462; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_463; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_464; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_465; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_466; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_467; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_468; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_469; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_470; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_471; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_472; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_473; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_474; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_475; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_476; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_477; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_478; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_479; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_480; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_481; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_482; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_483; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_484; // @[RAM_ST.scala 32:46]
  wire [8:0] _T_10; // @[RAM_ST.scala 32:46]
  wire [127:0] _T_17;
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_15_addr = ram__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_15_data = ram[ram__T_15_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_15_data = ram__T_15_addr >= 8'hf0 ? _RAND_1[127:0] : ram[ram__T_15_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_9_data = {_T_7,_T_4};
  assign ram__T_9_addr = _T[7:0];
  assign ram__T_9_mask = 1'h1;
  assign ram__T_9_en = write_elem_counter_valid;
  assign _GEN_1 = 8'h1 == WADDR ? 8'h1 : 8'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 8'h2 == WADDR ? 8'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 8'h3 == WADDR ? 8'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 8'h4 == WADDR ? 8'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 8'h5 == WADDR ? 8'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 8'h6 == WADDR ? 8'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 8'h7 == WADDR ? 8'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 8'h8 == WADDR ? 8'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 8'h9 == WADDR ? 8'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 8'ha == WADDR ? 8'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 8'hb == WADDR ? 8'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 8'hc == WADDR ? 8'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 8'hd == WADDR ? 8'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 8'he == WADDR ? 8'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 8'hf == WADDR ? 8'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 8'h10 == WADDR ? 8'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 8'h11 == WADDR ? 8'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 8'h12 == WADDR ? 8'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 8'h13 == WADDR ? 8'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 8'h14 == WADDR ? 8'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 8'h15 == WADDR ? 8'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 8'h16 == WADDR ? 8'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 8'h17 == WADDR ? 8'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 8'h18 == WADDR ? 8'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 8'h19 == WADDR ? 8'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 8'h1a == WADDR ? 8'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 8'h1b == WADDR ? 8'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 8'h1c == WADDR ? 8'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 8'h1d == WADDR ? 8'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 8'h1e == WADDR ? 8'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 8'h1f == WADDR ? 8'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 8'h20 == WADDR ? 8'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 8'h21 == WADDR ? 8'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 8'h22 == WADDR ? 8'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 8'h23 == WADDR ? 8'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 8'h24 == WADDR ? 8'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 8'h25 == WADDR ? 8'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 8'h26 == WADDR ? 8'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 8'h27 == WADDR ? 8'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 8'h28 == WADDR ? 8'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 8'h29 == WADDR ? 8'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 8'h2a == WADDR ? 8'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 8'h2b == WADDR ? 8'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 8'h2c == WADDR ? 8'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 8'h2d == WADDR ? 8'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 8'h2e == WADDR ? 8'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 8'h2f == WADDR ? 8'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 8'h30 == WADDR ? 8'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 8'h31 == WADDR ? 8'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 8'h32 == WADDR ? 8'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 8'h33 == WADDR ? 8'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 8'h34 == WADDR ? 8'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 8'h35 == WADDR ? 8'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 8'h36 == WADDR ? 8'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 8'h37 == WADDR ? 8'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 8'h38 == WADDR ? 8'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 8'h39 == WADDR ? 8'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 8'h3a == WADDR ? 8'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 8'h3b == WADDR ? 8'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 8'h3c == WADDR ? 8'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 8'h3d == WADDR ? 8'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 8'h3e == WADDR ? 8'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 8'h3f == WADDR ? 8'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 8'h40 == WADDR ? 8'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 8'h41 == WADDR ? 8'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 8'h42 == WADDR ? 8'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 8'h43 == WADDR ? 8'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 8'h44 == WADDR ? 8'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 8'h45 == WADDR ? 8'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 8'h46 == WADDR ? 8'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 8'h47 == WADDR ? 8'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 8'h48 == WADDR ? 8'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 8'h49 == WADDR ? 8'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 8'h4a == WADDR ? 8'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 8'h4b == WADDR ? 8'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 8'h4c == WADDR ? 8'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 8'h4d == WADDR ? 8'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 8'h4e == WADDR ? 8'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 8'h4f == WADDR ? 8'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 8'h50 == WADDR ? 8'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 8'h51 == WADDR ? 8'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 8'h52 == WADDR ? 8'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 8'h53 == WADDR ? 8'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 8'h54 == WADDR ? 8'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 8'h55 == WADDR ? 8'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 8'h56 == WADDR ? 8'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 8'h57 == WADDR ? 8'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 8'h58 == WADDR ? 8'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 8'h59 == WADDR ? 8'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 8'h5a == WADDR ? 8'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 8'h5b == WADDR ? 8'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 8'h5c == WADDR ? 8'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 8'h5d == WADDR ? 8'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 8'h5e == WADDR ? 8'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 8'h5f == WADDR ? 8'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 8'h60 == WADDR ? 8'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 8'h61 == WADDR ? 8'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 8'h62 == WADDR ? 8'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 8'h63 == WADDR ? 8'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 8'h64 == WADDR ? 8'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 8'h65 == WADDR ? 8'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 8'h66 == WADDR ? 8'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 8'h67 == WADDR ? 8'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 8'h68 == WADDR ? 8'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 8'h69 == WADDR ? 8'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 8'h6a == WADDR ? 8'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 8'h6b == WADDR ? 8'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 8'h6c == WADDR ? 8'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 8'h6d == WADDR ? 8'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 8'h6e == WADDR ? 8'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 8'h6f == WADDR ? 8'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 8'h70 == WADDR ? 8'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 8'h71 == WADDR ? 8'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 8'h72 == WADDR ? 8'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 8'h73 == WADDR ? 8'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 8'h74 == WADDR ? 8'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 8'h75 == WADDR ? 8'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 8'h76 == WADDR ? 8'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 8'h77 == WADDR ? 8'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _GEN_120 = 8'h78 == WADDR ? 8'h78 : _GEN_119; // @[RAM_ST.scala 31:71]
  assign _GEN_121 = 8'h79 == WADDR ? 8'h79 : _GEN_120; // @[RAM_ST.scala 31:71]
  assign _GEN_122 = 8'h7a == WADDR ? 8'h7a : _GEN_121; // @[RAM_ST.scala 31:71]
  assign _GEN_123 = 8'h7b == WADDR ? 8'h7b : _GEN_122; // @[RAM_ST.scala 31:71]
  assign _GEN_124 = 8'h7c == WADDR ? 8'h7c : _GEN_123; // @[RAM_ST.scala 31:71]
  assign _GEN_125 = 8'h7d == WADDR ? 8'h7d : _GEN_124; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 8'h7e == WADDR ? 8'h7e : _GEN_125; // @[RAM_ST.scala 31:71]
  assign _GEN_127 = 8'h7f == WADDR ? 8'h7f : _GEN_126; // @[RAM_ST.scala 31:71]
  assign _GEN_128 = 8'h80 == WADDR ? 8'h80 : _GEN_127; // @[RAM_ST.scala 31:71]
  assign _GEN_129 = 8'h81 == WADDR ? 8'h81 : _GEN_128; // @[RAM_ST.scala 31:71]
  assign _GEN_130 = 8'h82 == WADDR ? 8'h82 : _GEN_129; // @[RAM_ST.scala 31:71]
  assign _GEN_131 = 8'h83 == WADDR ? 8'h83 : _GEN_130; // @[RAM_ST.scala 31:71]
  assign _GEN_132 = 8'h84 == WADDR ? 8'h84 : _GEN_131; // @[RAM_ST.scala 31:71]
  assign _GEN_133 = 8'h85 == WADDR ? 8'h85 : _GEN_132; // @[RAM_ST.scala 31:71]
  assign _GEN_134 = 8'h86 == WADDR ? 8'h86 : _GEN_133; // @[RAM_ST.scala 31:71]
  assign _GEN_135 = 8'h87 == WADDR ? 8'h87 : _GEN_134; // @[RAM_ST.scala 31:71]
  assign _GEN_136 = 8'h88 == WADDR ? 8'h88 : _GEN_135; // @[RAM_ST.scala 31:71]
  assign _GEN_137 = 8'h89 == WADDR ? 8'h89 : _GEN_136; // @[RAM_ST.scala 31:71]
  assign _GEN_138 = 8'h8a == WADDR ? 8'h8a : _GEN_137; // @[RAM_ST.scala 31:71]
  assign _GEN_139 = 8'h8b == WADDR ? 8'h8b : _GEN_138; // @[RAM_ST.scala 31:71]
  assign _GEN_140 = 8'h8c == WADDR ? 8'h8c : _GEN_139; // @[RAM_ST.scala 31:71]
  assign _GEN_141 = 8'h8d == WADDR ? 8'h8d : _GEN_140; // @[RAM_ST.scala 31:71]
  assign _GEN_142 = 8'h8e == WADDR ? 8'h8e : _GEN_141; // @[RAM_ST.scala 31:71]
  assign _GEN_143 = 8'h8f == WADDR ? 8'h8f : _GEN_142; // @[RAM_ST.scala 31:71]
  assign _GEN_144 = 8'h90 == WADDR ? 8'h90 : _GEN_143; // @[RAM_ST.scala 31:71]
  assign _GEN_145 = 8'h91 == WADDR ? 8'h91 : _GEN_144; // @[RAM_ST.scala 31:71]
  assign _GEN_146 = 8'h92 == WADDR ? 8'h92 : _GEN_145; // @[RAM_ST.scala 31:71]
  assign _GEN_147 = 8'h93 == WADDR ? 8'h93 : _GEN_146; // @[RAM_ST.scala 31:71]
  assign _GEN_148 = 8'h94 == WADDR ? 8'h94 : _GEN_147; // @[RAM_ST.scala 31:71]
  assign _GEN_149 = 8'h95 == WADDR ? 8'h95 : _GEN_148; // @[RAM_ST.scala 31:71]
  assign _GEN_150 = 8'h96 == WADDR ? 8'h96 : _GEN_149; // @[RAM_ST.scala 31:71]
  assign _GEN_151 = 8'h97 == WADDR ? 8'h97 : _GEN_150; // @[RAM_ST.scala 31:71]
  assign _GEN_152 = 8'h98 == WADDR ? 8'h98 : _GEN_151; // @[RAM_ST.scala 31:71]
  assign _GEN_153 = 8'h99 == WADDR ? 8'h99 : _GEN_152; // @[RAM_ST.scala 31:71]
  assign _GEN_154 = 8'h9a == WADDR ? 8'h9a : _GEN_153; // @[RAM_ST.scala 31:71]
  assign _GEN_155 = 8'h9b == WADDR ? 8'h9b : _GEN_154; // @[RAM_ST.scala 31:71]
  assign _GEN_156 = 8'h9c == WADDR ? 8'h9c : _GEN_155; // @[RAM_ST.scala 31:71]
  assign _GEN_157 = 8'h9d == WADDR ? 8'h9d : _GEN_156; // @[RAM_ST.scala 31:71]
  assign _GEN_158 = 8'h9e == WADDR ? 8'h9e : _GEN_157; // @[RAM_ST.scala 31:71]
  assign _GEN_159 = 8'h9f == WADDR ? 8'h9f : _GEN_158; // @[RAM_ST.scala 31:71]
  assign _GEN_160 = 8'ha0 == WADDR ? 8'ha0 : _GEN_159; // @[RAM_ST.scala 31:71]
  assign _GEN_161 = 8'ha1 == WADDR ? 8'ha1 : _GEN_160; // @[RAM_ST.scala 31:71]
  assign _GEN_162 = 8'ha2 == WADDR ? 8'ha2 : _GEN_161; // @[RAM_ST.scala 31:71]
  assign _GEN_163 = 8'ha3 == WADDR ? 8'ha3 : _GEN_162; // @[RAM_ST.scala 31:71]
  assign _GEN_164 = 8'ha4 == WADDR ? 8'ha4 : _GEN_163; // @[RAM_ST.scala 31:71]
  assign _GEN_165 = 8'ha5 == WADDR ? 8'ha5 : _GEN_164; // @[RAM_ST.scala 31:71]
  assign _GEN_166 = 8'ha6 == WADDR ? 8'ha6 : _GEN_165; // @[RAM_ST.scala 31:71]
  assign _GEN_167 = 8'ha7 == WADDR ? 8'ha7 : _GEN_166; // @[RAM_ST.scala 31:71]
  assign _GEN_168 = 8'ha8 == WADDR ? 8'ha8 : _GEN_167; // @[RAM_ST.scala 31:71]
  assign _GEN_169 = 8'ha9 == WADDR ? 8'ha9 : _GEN_168; // @[RAM_ST.scala 31:71]
  assign _GEN_170 = 8'haa == WADDR ? 8'haa : _GEN_169; // @[RAM_ST.scala 31:71]
  assign _GEN_171 = 8'hab == WADDR ? 8'hab : _GEN_170; // @[RAM_ST.scala 31:71]
  assign _GEN_172 = 8'hac == WADDR ? 8'hac : _GEN_171; // @[RAM_ST.scala 31:71]
  assign _GEN_173 = 8'had == WADDR ? 8'had : _GEN_172; // @[RAM_ST.scala 31:71]
  assign _GEN_174 = 8'hae == WADDR ? 8'hae : _GEN_173; // @[RAM_ST.scala 31:71]
  assign _GEN_175 = 8'haf == WADDR ? 8'haf : _GEN_174; // @[RAM_ST.scala 31:71]
  assign _GEN_176 = 8'hb0 == WADDR ? 8'hb0 : _GEN_175; // @[RAM_ST.scala 31:71]
  assign _GEN_177 = 8'hb1 == WADDR ? 8'hb1 : _GEN_176; // @[RAM_ST.scala 31:71]
  assign _GEN_178 = 8'hb2 == WADDR ? 8'hb2 : _GEN_177; // @[RAM_ST.scala 31:71]
  assign _GEN_179 = 8'hb3 == WADDR ? 8'hb3 : _GEN_178; // @[RAM_ST.scala 31:71]
  assign _GEN_180 = 8'hb4 == WADDR ? 8'hb4 : _GEN_179; // @[RAM_ST.scala 31:71]
  assign _GEN_181 = 8'hb5 == WADDR ? 8'hb5 : _GEN_180; // @[RAM_ST.scala 31:71]
  assign _GEN_182 = 8'hb6 == WADDR ? 8'hb6 : _GEN_181; // @[RAM_ST.scala 31:71]
  assign _GEN_183 = 8'hb7 == WADDR ? 8'hb7 : _GEN_182; // @[RAM_ST.scala 31:71]
  assign _GEN_184 = 8'hb8 == WADDR ? 8'hb8 : _GEN_183; // @[RAM_ST.scala 31:71]
  assign _GEN_185 = 8'hb9 == WADDR ? 8'hb9 : _GEN_184; // @[RAM_ST.scala 31:71]
  assign _GEN_186 = 8'hba == WADDR ? 8'hba : _GEN_185; // @[RAM_ST.scala 31:71]
  assign _GEN_187 = 8'hbb == WADDR ? 8'hbb : _GEN_186; // @[RAM_ST.scala 31:71]
  assign _GEN_188 = 8'hbc == WADDR ? 8'hbc : _GEN_187; // @[RAM_ST.scala 31:71]
  assign _GEN_189 = 8'hbd == WADDR ? 8'hbd : _GEN_188; // @[RAM_ST.scala 31:71]
  assign _GEN_190 = 8'hbe == WADDR ? 8'hbe : _GEN_189; // @[RAM_ST.scala 31:71]
  assign _GEN_191 = 8'hbf == WADDR ? 8'hbf : _GEN_190; // @[RAM_ST.scala 31:71]
  assign _GEN_192 = 8'hc0 == WADDR ? 8'hc0 : _GEN_191; // @[RAM_ST.scala 31:71]
  assign _GEN_193 = 8'hc1 == WADDR ? 8'hc1 : _GEN_192; // @[RAM_ST.scala 31:71]
  assign _GEN_194 = 8'hc2 == WADDR ? 8'hc2 : _GEN_193; // @[RAM_ST.scala 31:71]
  assign _GEN_195 = 8'hc3 == WADDR ? 8'hc3 : _GEN_194; // @[RAM_ST.scala 31:71]
  assign _GEN_196 = 8'hc4 == WADDR ? 8'hc4 : _GEN_195; // @[RAM_ST.scala 31:71]
  assign _GEN_197 = 8'hc5 == WADDR ? 8'hc5 : _GEN_196; // @[RAM_ST.scala 31:71]
  assign _GEN_198 = 8'hc6 == WADDR ? 8'hc6 : _GEN_197; // @[RAM_ST.scala 31:71]
  assign _GEN_199 = 8'hc7 == WADDR ? 8'hc7 : _GEN_198; // @[RAM_ST.scala 31:71]
  assign _GEN_200 = 8'hc8 == WADDR ? 8'hc8 : _GEN_199; // @[RAM_ST.scala 31:71]
  assign _GEN_201 = 8'hc9 == WADDR ? 8'hc9 : _GEN_200; // @[RAM_ST.scala 31:71]
  assign _GEN_202 = 8'hca == WADDR ? 8'hca : _GEN_201; // @[RAM_ST.scala 31:71]
  assign _GEN_203 = 8'hcb == WADDR ? 8'hcb : _GEN_202; // @[RAM_ST.scala 31:71]
  assign _GEN_204 = 8'hcc == WADDR ? 8'hcc : _GEN_203; // @[RAM_ST.scala 31:71]
  assign _GEN_205 = 8'hcd == WADDR ? 8'hcd : _GEN_204; // @[RAM_ST.scala 31:71]
  assign _GEN_206 = 8'hce == WADDR ? 8'hce : _GEN_205; // @[RAM_ST.scala 31:71]
  assign _GEN_207 = 8'hcf == WADDR ? 8'hcf : _GEN_206; // @[RAM_ST.scala 31:71]
  assign _GEN_208 = 8'hd0 == WADDR ? 8'hd0 : _GEN_207; // @[RAM_ST.scala 31:71]
  assign _GEN_209 = 8'hd1 == WADDR ? 8'hd1 : _GEN_208; // @[RAM_ST.scala 31:71]
  assign _GEN_210 = 8'hd2 == WADDR ? 8'hd2 : _GEN_209; // @[RAM_ST.scala 31:71]
  assign _GEN_211 = 8'hd3 == WADDR ? 8'hd3 : _GEN_210; // @[RAM_ST.scala 31:71]
  assign _GEN_212 = 8'hd4 == WADDR ? 8'hd4 : _GEN_211; // @[RAM_ST.scala 31:71]
  assign _GEN_213 = 8'hd5 == WADDR ? 8'hd5 : _GEN_212; // @[RAM_ST.scala 31:71]
  assign _GEN_214 = 8'hd6 == WADDR ? 8'hd6 : _GEN_213; // @[RAM_ST.scala 31:71]
  assign _GEN_215 = 8'hd7 == WADDR ? 8'hd7 : _GEN_214; // @[RAM_ST.scala 31:71]
  assign _GEN_216 = 8'hd8 == WADDR ? 8'hd8 : _GEN_215; // @[RAM_ST.scala 31:71]
  assign _GEN_217 = 8'hd9 == WADDR ? 8'hd9 : _GEN_216; // @[RAM_ST.scala 31:71]
  assign _GEN_218 = 8'hda == WADDR ? 8'hda : _GEN_217; // @[RAM_ST.scala 31:71]
  assign _GEN_219 = 8'hdb == WADDR ? 8'hdb : _GEN_218; // @[RAM_ST.scala 31:71]
  assign _GEN_220 = 8'hdc == WADDR ? 8'hdc : _GEN_219; // @[RAM_ST.scala 31:71]
  assign _GEN_221 = 8'hdd == WADDR ? 8'hdd : _GEN_220; // @[RAM_ST.scala 31:71]
  assign _GEN_222 = 8'hde == WADDR ? 8'hde : _GEN_221; // @[RAM_ST.scala 31:71]
  assign _GEN_223 = 8'hdf == WADDR ? 8'hdf : _GEN_222; // @[RAM_ST.scala 31:71]
  assign _GEN_224 = 8'he0 == WADDR ? 8'he0 : _GEN_223; // @[RAM_ST.scala 31:71]
  assign _GEN_225 = 8'he1 == WADDR ? 8'he1 : _GEN_224; // @[RAM_ST.scala 31:71]
  assign _GEN_226 = 8'he2 == WADDR ? 8'he2 : _GEN_225; // @[RAM_ST.scala 31:71]
  assign _GEN_227 = 8'he3 == WADDR ? 8'he3 : _GEN_226; // @[RAM_ST.scala 31:71]
  assign _GEN_228 = 8'he4 == WADDR ? 8'he4 : _GEN_227; // @[RAM_ST.scala 31:71]
  assign _GEN_229 = 8'he5 == WADDR ? 8'he5 : _GEN_228; // @[RAM_ST.scala 31:71]
  assign _GEN_230 = 8'he6 == WADDR ? 8'he6 : _GEN_229; // @[RAM_ST.scala 31:71]
  assign _GEN_231 = 8'he7 == WADDR ? 8'he7 : _GEN_230; // @[RAM_ST.scala 31:71]
  assign _GEN_232 = 8'he8 == WADDR ? 8'he8 : _GEN_231; // @[RAM_ST.scala 31:71]
  assign _GEN_233 = 8'he9 == WADDR ? 8'he9 : _GEN_232; // @[RAM_ST.scala 31:71]
  assign _GEN_234 = 8'hea == WADDR ? 8'hea : _GEN_233; // @[RAM_ST.scala 31:71]
  assign _GEN_235 = 8'heb == WADDR ? 8'heb : _GEN_234; // @[RAM_ST.scala 31:71]
  assign _GEN_236 = 8'hec == WADDR ? 8'hec : _GEN_235; // @[RAM_ST.scala 31:71]
  assign _GEN_237 = 8'hed == WADDR ? 8'hed : _GEN_236; // @[RAM_ST.scala 31:71]
  assign _GEN_238 = 8'hee == WADDR ? 8'hee : _GEN_237; // @[RAM_ST.scala 31:71]
  assign _GEN_239 = 8'hef == WADDR ? 8'hef : _GEN_238; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_239}; // @[RAM_ST.scala 31:71]
  assign _T_4 = {WDATA_3,WDATA_2,WDATA_1,WDATA_0}; // @[RAM_ST.scala 31:115]
  assign _T_7 = {WDATA_7,WDATA_6,WDATA_5,WDATA_4}; // @[RAM_ST.scala 31:115]
  assign _GEN_246 = 8'h1 == RADDR ? 8'h1 : 8'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_247 = 8'h2 == RADDR ? 8'h2 : _GEN_246; // @[RAM_ST.scala 32:46]
  assign _GEN_248 = 8'h3 == RADDR ? 8'h3 : _GEN_247; // @[RAM_ST.scala 32:46]
  assign _GEN_249 = 8'h4 == RADDR ? 8'h4 : _GEN_248; // @[RAM_ST.scala 32:46]
  assign _GEN_250 = 8'h5 == RADDR ? 8'h5 : _GEN_249; // @[RAM_ST.scala 32:46]
  assign _GEN_251 = 8'h6 == RADDR ? 8'h6 : _GEN_250; // @[RAM_ST.scala 32:46]
  assign _GEN_252 = 8'h7 == RADDR ? 8'h7 : _GEN_251; // @[RAM_ST.scala 32:46]
  assign _GEN_253 = 8'h8 == RADDR ? 8'h8 : _GEN_252; // @[RAM_ST.scala 32:46]
  assign _GEN_254 = 8'h9 == RADDR ? 8'h9 : _GEN_253; // @[RAM_ST.scala 32:46]
  assign _GEN_255 = 8'ha == RADDR ? 8'ha : _GEN_254; // @[RAM_ST.scala 32:46]
  assign _GEN_256 = 8'hb == RADDR ? 8'hb : _GEN_255; // @[RAM_ST.scala 32:46]
  assign _GEN_257 = 8'hc == RADDR ? 8'hc : _GEN_256; // @[RAM_ST.scala 32:46]
  assign _GEN_258 = 8'hd == RADDR ? 8'hd : _GEN_257; // @[RAM_ST.scala 32:46]
  assign _GEN_259 = 8'he == RADDR ? 8'he : _GEN_258; // @[RAM_ST.scala 32:46]
  assign _GEN_260 = 8'hf == RADDR ? 8'hf : _GEN_259; // @[RAM_ST.scala 32:46]
  assign _GEN_261 = 8'h10 == RADDR ? 8'h10 : _GEN_260; // @[RAM_ST.scala 32:46]
  assign _GEN_262 = 8'h11 == RADDR ? 8'h11 : _GEN_261; // @[RAM_ST.scala 32:46]
  assign _GEN_263 = 8'h12 == RADDR ? 8'h12 : _GEN_262; // @[RAM_ST.scala 32:46]
  assign _GEN_264 = 8'h13 == RADDR ? 8'h13 : _GEN_263; // @[RAM_ST.scala 32:46]
  assign _GEN_265 = 8'h14 == RADDR ? 8'h14 : _GEN_264; // @[RAM_ST.scala 32:46]
  assign _GEN_266 = 8'h15 == RADDR ? 8'h15 : _GEN_265; // @[RAM_ST.scala 32:46]
  assign _GEN_267 = 8'h16 == RADDR ? 8'h16 : _GEN_266; // @[RAM_ST.scala 32:46]
  assign _GEN_268 = 8'h17 == RADDR ? 8'h17 : _GEN_267; // @[RAM_ST.scala 32:46]
  assign _GEN_269 = 8'h18 == RADDR ? 8'h18 : _GEN_268; // @[RAM_ST.scala 32:46]
  assign _GEN_270 = 8'h19 == RADDR ? 8'h19 : _GEN_269; // @[RAM_ST.scala 32:46]
  assign _GEN_271 = 8'h1a == RADDR ? 8'h1a : _GEN_270; // @[RAM_ST.scala 32:46]
  assign _GEN_272 = 8'h1b == RADDR ? 8'h1b : _GEN_271; // @[RAM_ST.scala 32:46]
  assign _GEN_273 = 8'h1c == RADDR ? 8'h1c : _GEN_272; // @[RAM_ST.scala 32:46]
  assign _GEN_274 = 8'h1d == RADDR ? 8'h1d : _GEN_273; // @[RAM_ST.scala 32:46]
  assign _GEN_275 = 8'h1e == RADDR ? 8'h1e : _GEN_274; // @[RAM_ST.scala 32:46]
  assign _GEN_276 = 8'h1f == RADDR ? 8'h1f : _GEN_275; // @[RAM_ST.scala 32:46]
  assign _GEN_277 = 8'h20 == RADDR ? 8'h20 : _GEN_276; // @[RAM_ST.scala 32:46]
  assign _GEN_278 = 8'h21 == RADDR ? 8'h21 : _GEN_277; // @[RAM_ST.scala 32:46]
  assign _GEN_279 = 8'h22 == RADDR ? 8'h22 : _GEN_278; // @[RAM_ST.scala 32:46]
  assign _GEN_280 = 8'h23 == RADDR ? 8'h23 : _GEN_279; // @[RAM_ST.scala 32:46]
  assign _GEN_281 = 8'h24 == RADDR ? 8'h24 : _GEN_280; // @[RAM_ST.scala 32:46]
  assign _GEN_282 = 8'h25 == RADDR ? 8'h25 : _GEN_281; // @[RAM_ST.scala 32:46]
  assign _GEN_283 = 8'h26 == RADDR ? 8'h26 : _GEN_282; // @[RAM_ST.scala 32:46]
  assign _GEN_284 = 8'h27 == RADDR ? 8'h27 : _GEN_283; // @[RAM_ST.scala 32:46]
  assign _GEN_285 = 8'h28 == RADDR ? 8'h28 : _GEN_284; // @[RAM_ST.scala 32:46]
  assign _GEN_286 = 8'h29 == RADDR ? 8'h29 : _GEN_285; // @[RAM_ST.scala 32:46]
  assign _GEN_287 = 8'h2a == RADDR ? 8'h2a : _GEN_286; // @[RAM_ST.scala 32:46]
  assign _GEN_288 = 8'h2b == RADDR ? 8'h2b : _GEN_287; // @[RAM_ST.scala 32:46]
  assign _GEN_289 = 8'h2c == RADDR ? 8'h2c : _GEN_288; // @[RAM_ST.scala 32:46]
  assign _GEN_290 = 8'h2d == RADDR ? 8'h2d : _GEN_289; // @[RAM_ST.scala 32:46]
  assign _GEN_291 = 8'h2e == RADDR ? 8'h2e : _GEN_290; // @[RAM_ST.scala 32:46]
  assign _GEN_292 = 8'h2f == RADDR ? 8'h2f : _GEN_291; // @[RAM_ST.scala 32:46]
  assign _GEN_293 = 8'h30 == RADDR ? 8'h30 : _GEN_292; // @[RAM_ST.scala 32:46]
  assign _GEN_294 = 8'h31 == RADDR ? 8'h31 : _GEN_293; // @[RAM_ST.scala 32:46]
  assign _GEN_295 = 8'h32 == RADDR ? 8'h32 : _GEN_294; // @[RAM_ST.scala 32:46]
  assign _GEN_296 = 8'h33 == RADDR ? 8'h33 : _GEN_295; // @[RAM_ST.scala 32:46]
  assign _GEN_297 = 8'h34 == RADDR ? 8'h34 : _GEN_296; // @[RAM_ST.scala 32:46]
  assign _GEN_298 = 8'h35 == RADDR ? 8'h35 : _GEN_297; // @[RAM_ST.scala 32:46]
  assign _GEN_299 = 8'h36 == RADDR ? 8'h36 : _GEN_298; // @[RAM_ST.scala 32:46]
  assign _GEN_300 = 8'h37 == RADDR ? 8'h37 : _GEN_299; // @[RAM_ST.scala 32:46]
  assign _GEN_301 = 8'h38 == RADDR ? 8'h38 : _GEN_300; // @[RAM_ST.scala 32:46]
  assign _GEN_302 = 8'h39 == RADDR ? 8'h39 : _GEN_301; // @[RAM_ST.scala 32:46]
  assign _GEN_303 = 8'h3a == RADDR ? 8'h3a : _GEN_302; // @[RAM_ST.scala 32:46]
  assign _GEN_304 = 8'h3b == RADDR ? 8'h3b : _GEN_303; // @[RAM_ST.scala 32:46]
  assign _GEN_305 = 8'h3c == RADDR ? 8'h3c : _GEN_304; // @[RAM_ST.scala 32:46]
  assign _GEN_306 = 8'h3d == RADDR ? 8'h3d : _GEN_305; // @[RAM_ST.scala 32:46]
  assign _GEN_307 = 8'h3e == RADDR ? 8'h3e : _GEN_306; // @[RAM_ST.scala 32:46]
  assign _GEN_308 = 8'h3f == RADDR ? 8'h3f : _GEN_307; // @[RAM_ST.scala 32:46]
  assign _GEN_309 = 8'h40 == RADDR ? 8'h40 : _GEN_308; // @[RAM_ST.scala 32:46]
  assign _GEN_310 = 8'h41 == RADDR ? 8'h41 : _GEN_309; // @[RAM_ST.scala 32:46]
  assign _GEN_311 = 8'h42 == RADDR ? 8'h42 : _GEN_310; // @[RAM_ST.scala 32:46]
  assign _GEN_312 = 8'h43 == RADDR ? 8'h43 : _GEN_311; // @[RAM_ST.scala 32:46]
  assign _GEN_313 = 8'h44 == RADDR ? 8'h44 : _GEN_312; // @[RAM_ST.scala 32:46]
  assign _GEN_314 = 8'h45 == RADDR ? 8'h45 : _GEN_313; // @[RAM_ST.scala 32:46]
  assign _GEN_315 = 8'h46 == RADDR ? 8'h46 : _GEN_314; // @[RAM_ST.scala 32:46]
  assign _GEN_316 = 8'h47 == RADDR ? 8'h47 : _GEN_315; // @[RAM_ST.scala 32:46]
  assign _GEN_317 = 8'h48 == RADDR ? 8'h48 : _GEN_316; // @[RAM_ST.scala 32:46]
  assign _GEN_318 = 8'h49 == RADDR ? 8'h49 : _GEN_317; // @[RAM_ST.scala 32:46]
  assign _GEN_319 = 8'h4a == RADDR ? 8'h4a : _GEN_318; // @[RAM_ST.scala 32:46]
  assign _GEN_320 = 8'h4b == RADDR ? 8'h4b : _GEN_319; // @[RAM_ST.scala 32:46]
  assign _GEN_321 = 8'h4c == RADDR ? 8'h4c : _GEN_320; // @[RAM_ST.scala 32:46]
  assign _GEN_322 = 8'h4d == RADDR ? 8'h4d : _GEN_321; // @[RAM_ST.scala 32:46]
  assign _GEN_323 = 8'h4e == RADDR ? 8'h4e : _GEN_322; // @[RAM_ST.scala 32:46]
  assign _GEN_324 = 8'h4f == RADDR ? 8'h4f : _GEN_323; // @[RAM_ST.scala 32:46]
  assign _GEN_325 = 8'h50 == RADDR ? 8'h50 : _GEN_324; // @[RAM_ST.scala 32:46]
  assign _GEN_326 = 8'h51 == RADDR ? 8'h51 : _GEN_325; // @[RAM_ST.scala 32:46]
  assign _GEN_327 = 8'h52 == RADDR ? 8'h52 : _GEN_326; // @[RAM_ST.scala 32:46]
  assign _GEN_328 = 8'h53 == RADDR ? 8'h53 : _GEN_327; // @[RAM_ST.scala 32:46]
  assign _GEN_329 = 8'h54 == RADDR ? 8'h54 : _GEN_328; // @[RAM_ST.scala 32:46]
  assign _GEN_330 = 8'h55 == RADDR ? 8'h55 : _GEN_329; // @[RAM_ST.scala 32:46]
  assign _GEN_331 = 8'h56 == RADDR ? 8'h56 : _GEN_330; // @[RAM_ST.scala 32:46]
  assign _GEN_332 = 8'h57 == RADDR ? 8'h57 : _GEN_331; // @[RAM_ST.scala 32:46]
  assign _GEN_333 = 8'h58 == RADDR ? 8'h58 : _GEN_332; // @[RAM_ST.scala 32:46]
  assign _GEN_334 = 8'h59 == RADDR ? 8'h59 : _GEN_333; // @[RAM_ST.scala 32:46]
  assign _GEN_335 = 8'h5a == RADDR ? 8'h5a : _GEN_334; // @[RAM_ST.scala 32:46]
  assign _GEN_336 = 8'h5b == RADDR ? 8'h5b : _GEN_335; // @[RAM_ST.scala 32:46]
  assign _GEN_337 = 8'h5c == RADDR ? 8'h5c : _GEN_336; // @[RAM_ST.scala 32:46]
  assign _GEN_338 = 8'h5d == RADDR ? 8'h5d : _GEN_337; // @[RAM_ST.scala 32:46]
  assign _GEN_339 = 8'h5e == RADDR ? 8'h5e : _GEN_338; // @[RAM_ST.scala 32:46]
  assign _GEN_340 = 8'h5f == RADDR ? 8'h5f : _GEN_339; // @[RAM_ST.scala 32:46]
  assign _GEN_341 = 8'h60 == RADDR ? 8'h60 : _GEN_340; // @[RAM_ST.scala 32:46]
  assign _GEN_342 = 8'h61 == RADDR ? 8'h61 : _GEN_341; // @[RAM_ST.scala 32:46]
  assign _GEN_343 = 8'h62 == RADDR ? 8'h62 : _GEN_342; // @[RAM_ST.scala 32:46]
  assign _GEN_344 = 8'h63 == RADDR ? 8'h63 : _GEN_343; // @[RAM_ST.scala 32:46]
  assign _GEN_345 = 8'h64 == RADDR ? 8'h64 : _GEN_344; // @[RAM_ST.scala 32:46]
  assign _GEN_346 = 8'h65 == RADDR ? 8'h65 : _GEN_345; // @[RAM_ST.scala 32:46]
  assign _GEN_347 = 8'h66 == RADDR ? 8'h66 : _GEN_346; // @[RAM_ST.scala 32:46]
  assign _GEN_348 = 8'h67 == RADDR ? 8'h67 : _GEN_347; // @[RAM_ST.scala 32:46]
  assign _GEN_349 = 8'h68 == RADDR ? 8'h68 : _GEN_348; // @[RAM_ST.scala 32:46]
  assign _GEN_350 = 8'h69 == RADDR ? 8'h69 : _GEN_349; // @[RAM_ST.scala 32:46]
  assign _GEN_351 = 8'h6a == RADDR ? 8'h6a : _GEN_350; // @[RAM_ST.scala 32:46]
  assign _GEN_352 = 8'h6b == RADDR ? 8'h6b : _GEN_351; // @[RAM_ST.scala 32:46]
  assign _GEN_353 = 8'h6c == RADDR ? 8'h6c : _GEN_352; // @[RAM_ST.scala 32:46]
  assign _GEN_354 = 8'h6d == RADDR ? 8'h6d : _GEN_353; // @[RAM_ST.scala 32:46]
  assign _GEN_355 = 8'h6e == RADDR ? 8'h6e : _GEN_354; // @[RAM_ST.scala 32:46]
  assign _GEN_356 = 8'h6f == RADDR ? 8'h6f : _GEN_355; // @[RAM_ST.scala 32:46]
  assign _GEN_357 = 8'h70 == RADDR ? 8'h70 : _GEN_356; // @[RAM_ST.scala 32:46]
  assign _GEN_358 = 8'h71 == RADDR ? 8'h71 : _GEN_357; // @[RAM_ST.scala 32:46]
  assign _GEN_359 = 8'h72 == RADDR ? 8'h72 : _GEN_358; // @[RAM_ST.scala 32:46]
  assign _GEN_360 = 8'h73 == RADDR ? 8'h73 : _GEN_359; // @[RAM_ST.scala 32:46]
  assign _GEN_361 = 8'h74 == RADDR ? 8'h74 : _GEN_360; // @[RAM_ST.scala 32:46]
  assign _GEN_362 = 8'h75 == RADDR ? 8'h75 : _GEN_361; // @[RAM_ST.scala 32:46]
  assign _GEN_363 = 8'h76 == RADDR ? 8'h76 : _GEN_362; // @[RAM_ST.scala 32:46]
  assign _GEN_364 = 8'h77 == RADDR ? 8'h77 : _GEN_363; // @[RAM_ST.scala 32:46]
  assign _GEN_365 = 8'h78 == RADDR ? 8'h78 : _GEN_364; // @[RAM_ST.scala 32:46]
  assign _GEN_366 = 8'h79 == RADDR ? 8'h79 : _GEN_365; // @[RAM_ST.scala 32:46]
  assign _GEN_367 = 8'h7a == RADDR ? 8'h7a : _GEN_366; // @[RAM_ST.scala 32:46]
  assign _GEN_368 = 8'h7b == RADDR ? 8'h7b : _GEN_367; // @[RAM_ST.scala 32:46]
  assign _GEN_369 = 8'h7c == RADDR ? 8'h7c : _GEN_368; // @[RAM_ST.scala 32:46]
  assign _GEN_370 = 8'h7d == RADDR ? 8'h7d : _GEN_369; // @[RAM_ST.scala 32:46]
  assign _GEN_371 = 8'h7e == RADDR ? 8'h7e : _GEN_370; // @[RAM_ST.scala 32:46]
  assign _GEN_372 = 8'h7f == RADDR ? 8'h7f : _GEN_371; // @[RAM_ST.scala 32:46]
  assign _GEN_373 = 8'h80 == RADDR ? 8'h80 : _GEN_372; // @[RAM_ST.scala 32:46]
  assign _GEN_374 = 8'h81 == RADDR ? 8'h81 : _GEN_373; // @[RAM_ST.scala 32:46]
  assign _GEN_375 = 8'h82 == RADDR ? 8'h82 : _GEN_374; // @[RAM_ST.scala 32:46]
  assign _GEN_376 = 8'h83 == RADDR ? 8'h83 : _GEN_375; // @[RAM_ST.scala 32:46]
  assign _GEN_377 = 8'h84 == RADDR ? 8'h84 : _GEN_376; // @[RAM_ST.scala 32:46]
  assign _GEN_378 = 8'h85 == RADDR ? 8'h85 : _GEN_377; // @[RAM_ST.scala 32:46]
  assign _GEN_379 = 8'h86 == RADDR ? 8'h86 : _GEN_378; // @[RAM_ST.scala 32:46]
  assign _GEN_380 = 8'h87 == RADDR ? 8'h87 : _GEN_379; // @[RAM_ST.scala 32:46]
  assign _GEN_381 = 8'h88 == RADDR ? 8'h88 : _GEN_380; // @[RAM_ST.scala 32:46]
  assign _GEN_382 = 8'h89 == RADDR ? 8'h89 : _GEN_381; // @[RAM_ST.scala 32:46]
  assign _GEN_383 = 8'h8a == RADDR ? 8'h8a : _GEN_382; // @[RAM_ST.scala 32:46]
  assign _GEN_384 = 8'h8b == RADDR ? 8'h8b : _GEN_383; // @[RAM_ST.scala 32:46]
  assign _GEN_385 = 8'h8c == RADDR ? 8'h8c : _GEN_384; // @[RAM_ST.scala 32:46]
  assign _GEN_386 = 8'h8d == RADDR ? 8'h8d : _GEN_385; // @[RAM_ST.scala 32:46]
  assign _GEN_387 = 8'h8e == RADDR ? 8'h8e : _GEN_386; // @[RAM_ST.scala 32:46]
  assign _GEN_388 = 8'h8f == RADDR ? 8'h8f : _GEN_387; // @[RAM_ST.scala 32:46]
  assign _GEN_389 = 8'h90 == RADDR ? 8'h90 : _GEN_388; // @[RAM_ST.scala 32:46]
  assign _GEN_390 = 8'h91 == RADDR ? 8'h91 : _GEN_389; // @[RAM_ST.scala 32:46]
  assign _GEN_391 = 8'h92 == RADDR ? 8'h92 : _GEN_390; // @[RAM_ST.scala 32:46]
  assign _GEN_392 = 8'h93 == RADDR ? 8'h93 : _GEN_391; // @[RAM_ST.scala 32:46]
  assign _GEN_393 = 8'h94 == RADDR ? 8'h94 : _GEN_392; // @[RAM_ST.scala 32:46]
  assign _GEN_394 = 8'h95 == RADDR ? 8'h95 : _GEN_393; // @[RAM_ST.scala 32:46]
  assign _GEN_395 = 8'h96 == RADDR ? 8'h96 : _GEN_394; // @[RAM_ST.scala 32:46]
  assign _GEN_396 = 8'h97 == RADDR ? 8'h97 : _GEN_395; // @[RAM_ST.scala 32:46]
  assign _GEN_397 = 8'h98 == RADDR ? 8'h98 : _GEN_396; // @[RAM_ST.scala 32:46]
  assign _GEN_398 = 8'h99 == RADDR ? 8'h99 : _GEN_397; // @[RAM_ST.scala 32:46]
  assign _GEN_399 = 8'h9a == RADDR ? 8'h9a : _GEN_398; // @[RAM_ST.scala 32:46]
  assign _GEN_400 = 8'h9b == RADDR ? 8'h9b : _GEN_399; // @[RAM_ST.scala 32:46]
  assign _GEN_401 = 8'h9c == RADDR ? 8'h9c : _GEN_400; // @[RAM_ST.scala 32:46]
  assign _GEN_402 = 8'h9d == RADDR ? 8'h9d : _GEN_401; // @[RAM_ST.scala 32:46]
  assign _GEN_403 = 8'h9e == RADDR ? 8'h9e : _GEN_402; // @[RAM_ST.scala 32:46]
  assign _GEN_404 = 8'h9f == RADDR ? 8'h9f : _GEN_403; // @[RAM_ST.scala 32:46]
  assign _GEN_405 = 8'ha0 == RADDR ? 8'ha0 : _GEN_404; // @[RAM_ST.scala 32:46]
  assign _GEN_406 = 8'ha1 == RADDR ? 8'ha1 : _GEN_405; // @[RAM_ST.scala 32:46]
  assign _GEN_407 = 8'ha2 == RADDR ? 8'ha2 : _GEN_406; // @[RAM_ST.scala 32:46]
  assign _GEN_408 = 8'ha3 == RADDR ? 8'ha3 : _GEN_407; // @[RAM_ST.scala 32:46]
  assign _GEN_409 = 8'ha4 == RADDR ? 8'ha4 : _GEN_408; // @[RAM_ST.scala 32:46]
  assign _GEN_410 = 8'ha5 == RADDR ? 8'ha5 : _GEN_409; // @[RAM_ST.scala 32:46]
  assign _GEN_411 = 8'ha6 == RADDR ? 8'ha6 : _GEN_410; // @[RAM_ST.scala 32:46]
  assign _GEN_412 = 8'ha7 == RADDR ? 8'ha7 : _GEN_411; // @[RAM_ST.scala 32:46]
  assign _GEN_413 = 8'ha8 == RADDR ? 8'ha8 : _GEN_412; // @[RAM_ST.scala 32:46]
  assign _GEN_414 = 8'ha9 == RADDR ? 8'ha9 : _GEN_413; // @[RAM_ST.scala 32:46]
  assign _GEN_415 = 8'haa == RADDR ? 8'haa : _GEN_414; // @[RAM_ST.scala 32:46]
  assign _GEN_416 = 8'hab == RADDR ? 8'hab : _GEN_415; // @[RAM_ST.scala 32:46]
  assign _GEN_417 = 8'hac == RADDR ? 8'hac : _GEN_416; // @[RAM_ST.scala 32:46]
  assign _GEN_418 = 8'had == RADDR ? 8'had : _GEN_417; // @[RAM_ST.scala 32:46]
  assign _GEN_419 = 8'hae == RADDR ? 8'hae : _GEN_418; // @[RAM_ST.scala 32:46]
  assign _GEN_420 = 8'haf == RADDR ? 8'haf : _GEN_419; // @[RAM_ST.scala 32:46]
  assign _GEN_421 = 8'hb0 == RADDR ? 8'hb0 : _GEN_420; // @[RAM_ST.scala 32:46]
  assign _GEN_422 = 8'hb1 == RADDR ? 8'hb1 : _GEN_421; // @[RAM_ST.scala 32:46]
  assign _GEN_423 = 8'hb2 == RADDR ? 8'hb2 : _GEN_422; // @[RAM_ST.scala 32:46]
  assign _GEN_424 = 8'hb3 == RADDR ? 8'hb3 : _GEN_423; // @[RAM_ST.scala 32:46]
  assign _GEN_425 = 8'hb4 == RADDR ? 8'hb4 : _GEN_424; // @[RAM_ST.scala 32:46]
  assign _GEN_426 = 8'hb5 == RADDR ? 8'hb5 : _GEN_425; // @[RAM_ST.scala 32:46]
  assign _GEN_427 = 8'hb6 == RADDR ? 8'hb6 : _GEN_426; // @[RAM_ST.scala 32:46]
  assign _GEN_428 = 8'hb7 == RADDR ? 8'hb7 : _GEN_427; // @[RAM_ST.scala 32:46]
  assign _GEN_429 = 8'hb8 == RADDR ? 8'hb8 : _GEN_428; // @[RAM_ST.scala 32:46]
  assign _GEN_430 = 8'hb9 == RADDR ? 8'hb9 : _GEN_429; // @[RAM_ST.scala 32:46]
  assign _GEN_431 = 8'hba == RADDR ? 8'hba : _GEN_430; // @[RAM_ST.scala 32:46]
  assign _GEN_432 = 8'hbb == RADDR ? 8'hbb : _GEN_431; // @[RAM_ST.scala 32:46]
  assign _GEN_433 = 8'hbc == RADDR ? 8'hbc : _GEN_432; // @[RAM_ST.scala 32:46]
  assign _GEN_434 = 8'hbd == RADDR ? 8'hbd : _GEN_433; // @[RAM_ST.scala 32:46]
  assign _GEN_435 = 8'hbe == RADDR ? 8'hbe : _GEN_434; // @[RAM_ST.scala 32:46]
  assign _GEN_436 = 8'hbf == RADDR ? 8'hbf : _GEN_435; // @[RAM_ST.scala 32:46]
  assign _GEN_437 = 8'hc0 == RADDR ? 8'hc0 : _GEN_436; // @[RAM_ST.scala 32:46]
  assign _GEN_438 = 8'hc1 == RADDR ? 8'hc1 : _GEN_437; // @[RAM_ST.scala 32:46]
  assign _GEN_439 = 8'hc2 == RADDR ? 8'hc2 : _GEN_438; // @[RAM_ST.scala 32:46]
  assign _GEN_440 = 8'hc3 == RADDR ? 8'hc3 : _GEN_439; // @[RAM_ST.scala 32:46]
  assign _GEN_441 = 8'hc4 == RADDR ? 8'hc4 : _GEN_440; // @[RAM_ST.scala 32:46]
  assign _GEN_442 = 8'hc5 == RADDR ? 8'hc5 : _GEN_441; // @[RAM_ST.scala 32:46]
  assign _GEN_443 = 8'hc6 == RADDR ? 8'hc6 : _GEN_442; // @[RAM_ST.scala 32:46]
  assign _GEN_444 = 8'hc7 == RADDR ? 8'hc7 : _GEN_443; // @[RAM_ST.scala 32:46]
  assign _GEN_445 = 8'hc8 == RADDR ? 8'hc8 : _GEN_444; // @[RAM_ST.scala 32:46]
  assign _GEN_446 = 8'hc9 == RADDR ? 8'hc9 : _GEN_445; // @[RAM_ST.scala 32:46]
  assign _GEN_447 = 8'hca == RADDR ? 8'hca : _GEN_446; // @[RAM_ST.scala 32:46]
  assign _GEN_448 = 8'hcb == RADDR ? 8'hcb : _GEN_447; // @[RAM_ST.scala 32:46]
  assign _GEN_449 = 8'hcc == RADDR ? 8'hcc : _GEN_448; // @[RAM_ST.scala 32:46]
  assign _GEN_450 = 8'hcd == RADDR ? 8'hcd : _GEN_449; // @[RAM_ST.scala 32:46]
  assign _GEN_451 = 8'hce == RADDR ? 8'hce : _GEN_450; // @[RAM_ST.scala 32:46]
  assign _GEN_452 = 8'hcf == RADDR ? 8'hcf : _GEN_451; // @[RAM_ST.scala 32:46]
  assign _GEN_453 = 8'hd0 == RADDR ? 8'hd0 : _GEN_452; // @[RAM_ST.scala 32:46]
  assign _GEN_454 = 8'hd1 == RADDR ? 8'hd1 : _GEN_453; // @[RAM_ST.scala 32:46]
  assign _GEN_455 = 8'hd2 == RADDR ? 8'hd2 : _GEN_454; // @[RAM_ST.scala 32:46]
  assign _GEN_456 = 8'hd3 == RADDR ? 8'hd3 : _GEN_455; // @[RAM_ST.scala 32:46]
  assign _GEN_457 = 8'hd4 == RADDR ? 8'hd4 : _GEN_456; // @[RAM_ST.scala 32:46]
  assign _GEN_458 = 8'hd5 == RADDR ? 8'hd5 : _GEN_457; // @[RAM_ST.scala 32:46]
  assign _GEN_459 = 8'hd6 == RADDR ? 8'hd6 : _GEN_458; // @[RAM_ST.scala 32:46]
  assign _GEN_460 = 8'hd7 == RADDR ? 8'hd7 : _GEN_459; // @[RAM_ST.scala 32:46]
  assign _GEN_461 = 8'hd8 == RADDR ? 8'hd8 : _GEN_460; // @[RAM_ST.scala 32:46]
  assign _GEN_462 = 8'hd9 == RADDR ? 8'hd9 : _GEN_461; // @[RAM_ST.scala 32:46]
  assign _GEN_463 = 8'hda == RADDR ? 8'hda : _GEN_462; // @[RAM_ST.scala 32:46]
  assign _GEN_464 = 8'hdb == RADDR ? 8'hdb : _GEN_463; // @[RAM_ST.scala 32:46]
  assign _GEN_465 = 8'hdc == RADDR ? 8'hdc : _GEN_464; // @[RAM_ST.scala 32:46]
  assign _GEN_466 = 8'hdd == RADDR ? 8'hdd : _GEN_465; // @[RAM_ST.scala 32:46]
  assign _GEN_467 = 8'hde == RADDR ? 8'hde : _GEN_466; // @[RAM_ST.scala 32:46]
  assign _GEN_468 = 8'hdf == RADDR ? 8'hdf : _GEN_467; // @[RAM_ST.scala 32:46]
  assign _GEN_469 = 8'he0 == RADDR ? 8'he0 : _GEN_468; // @[RAM_ST.scala 32:46]
  assign _GEN_470 = 8'he1 == RADDR ? 8'he1 : _GEN_469; // @[RAM_ST.scala 32:46]
  assign _GEN_471 = 8'he2 == RADDR ? 8'he2 : _GEN_470; // @[RAM_ST.scala 32:46]
  assign _GEN_472 = 8'he3 == RADDR ? 8'he3 : _GEN_471; // @[RAM_ST.scala 32:46]
  assign _GEN_473 = 8'he4 == RADDR ? 8'he4 : _GEN_472; // @[RAM_ST.scala 32:46]
  assign _GEN_474 = 8'he5 == RADDR ? 8'he5 : _GEN_473; // @[RAM_ST.scala 32:46]
  assign _GEN_475 = 8'he6 == RADDR ? 8'he6 : _GEN_474; // @[RAM_ST.scala 32:46]
  assign _GEN_476 = 8'he7 == RADDR ? 8'he7 : _GEN_475; // @[RAM_ST.scala 32:46]
  assign _GEN_477 = 8'he8 == RADDR ? 8'he8 : _GEN_476; // @[RAM_ST.scala 32:46]
  assign _GEN_478 = 8'he9 == RADDR ? 8'he9 : _GEN_477; // @[RAM_ST.scala 32:46]
  assign _GEN_479 = 8'hea == RADDR ? 8'hea : _GEN_478; // @[RAM_ST.scala 32:46]
  assign _GEN_480 = 8'heb == RADDR ? 8'heb : _GEN_479; // @[RAM_ST.scala 32:46]
  assign _GEN_481 = 8'hec == RADDR ? 8'hec : _GEN_480; // @[RAM_ST.scala 32:46]
  assign _GEN_482 = 8'hed == RADDR ? 8'hed : _GEN_481; // @[RAM_ST.scala 32:46]
  assign _GEN_483 = 8'hee == RADDR ? 8'hee : _GEN_482; // @[RAM_ST.scala 32:46]
  assign _GEN_484 = 8'hef == RADDR ? 8'hef : _GEN_483; // @[RAM_ST.scala 32:46]
  assign _T_10 = {{1'd0}, _GEN_484}; // @[RAM_ST.scala 32:46]
  assign _T_17 = ram__T_15_data;
  assign RDATA_0 = _T_17[15:0]; // @[RAM_ST.scala 32:9]
  assign RDATA_1 = _T_17[31:16]; // @[RAM_ST.scala 32:9]
  assign RDATA_2 = _T_17[47:32]; // @[RAM_ST.scala 32:9]
  assign RDATA_3 = _T_17[63:48]; // @[RAM_ST.scala 32:9]
  assign RDATA_4 = _T_17[79:64]; // @[RAM_ST.scala 32:9]
  assign RDATA_5 = _T_17[95:80]; // @[RAM_ST.scala 32:9]
  assign RDATA_6 = _T_17[111:96]; // @[RAM_ST.scala 32:9]
  assign RDATA_7 = _T_17[127:112]; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 240; initvar = initvar+1)
    ram[initvar] = _RAND_0[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_15_addr_pipe_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_9_en & ram__T_9_mask) begin
      ram[ram__T_9_addr] <= ram__T_9_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_15_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_15_addr_pipe_0 <= _T_10[7:0];
    end
  end
endmodule
module ShiftT(
  input         clock,
  input         reset,
  input         valid_up,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_0; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_1; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_2; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_3; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_4; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_5; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_6; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_7; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_0; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_1; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_2; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_3; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_4; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_5; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_6; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_7; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [7:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [7:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA_0(RAM_ST_RDATA_0),
    .RDATA_1(RAM_ST_RDATA_1),
    .RDATA_2(RAM_ST_RDATA_2),
    .RDATA_3(RAM_ST_RDATA_3),
    .RDATA_4(RAM_ST_RDATA_4),
    .RDATA_5(RAM_ST_RDATA_5),
    .RDATA_6(RAM_ST_RDATA_6),
    .RDATA_7(RAM_ST_RDATA_7),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA_0(RAM_ST_WDATA_0),
    .WDATA_1(RAM_ST_WDATA_1),
    .WDATA_2(RAM_ST_WDATA_2),
    .WDATA_3(RAM_ST_WDATA_3),
    .WDATA_4(RAM_ST_WDATA_4),
    .WDATA_5(RAM_ST_WDATA_5),
    .WDATA_6(RAM_ST_WDATA_6),
    .WDATA_7(RAM_ST_WDATA_7)
  );
  NestedCounters_1 NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 8'hef; // @[Counter.scala 37:24]
  assign _T_3 = value + 8'h1; // @[Counter.scala 38:22]
  assign O_0 = RAM_ST_RDATA_0; // @[ShiftT.scala 51:7]
  assign O_1 = RAM_ST_RDATA_1; // @[ShiftT.scala 51:7]
  assign O_2 = RAM_ST_RDATA_2; // @[ShiftT.scala 51:7]
  assign O_3 = RAM_ST_RDATA_3; // @[ShiftT.scala 51:7]
  assign O_4 = RAM_ST_RDATA_4; // @[ShiftT.scala 51:7]
  assign O_5 = RAM_ST_RDATA_5; // @[ShiftT.scala 51:7]
  assign O_6 = RAM_ST_RDATA_6; // @[ShiftT.scala 51:7]
  assign O_7 = RAM_ST_RDATA_7; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 8'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA_0 = I_0; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_1 = I_1; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_2 = I_2; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_3 = I_3; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_4 = I_4; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_5 = I_5; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_6 = I_6; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_7 = I_7; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 8'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 8'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:26]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_1; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_2; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_3; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_4; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_5; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_6; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_7; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_1; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_2; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_3; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_4; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_5; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_6; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_7; // @[ShiftTS.scala 32:26]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I_0(ShiftT_I_0),
    .I_1(ShiftT_I_1),
    .I_2(ShiftT_I_2),
    .I_3(ShiftT_I_3),
    .I_4(ShiftT_I_4),
    .I_5(ShiftT_I_5),
    .I_6(ShiftT_I_6),
    .I_7(ShiftT_I_7),
    .O_0(ShiftT_O_0),
    .O_1(ShiftT_O_1),
    .O_2(ShiftT_O_2),
    .O_3(ShiftT_O_3),
    .O_4(ShiftT_O_4),
    .O_5(ShiftT_O_5),
    .O_6(ShiftT_O_6),
    .O_7(ShiftT_O_7)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = ShiftT_O_1; // @[ShiftTS.scala 51:36]
  assign O_2 = ShiftT_O_2; // @[ShiftTS.scala 51:36]
  assign O_3 = ShiftT_O_3; // @[ShiftTS.scala 51:36]
  assign O_4 = ShiftT_O_4; // @[ShiftTS.scala 51:36]
  assign O_5 = ShiftT_O_5; // @[ShiftTS.scala 51:36]
  assign O_6 = ShiftT_O_6; // @[ShiftTS.scala 51:36]
  assign O_7 = ShiftT_O_7; // @[ShiftTS.scala 51:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 53:29]
  assign ShiftT_I_0 = I_0; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_1 = I_1; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_2 = I_2; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_3 = I_3; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_4 = I_4; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_5 = I_5; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_6 = I_6; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_7 = I_7; // @[ShiftTS.scala 50:25]
endmodule
module ShiftT_2(
  input         clock,
  input  [15:0] I_0,
  output [15:0] O_0
);
  reg [15:0] _T_0; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O_0 = _T_0; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= I_0;
  end
endmodule
module ShiftTS_2(
  input         clock,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  ShiftT_2 ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .I_0(ShiftT_I_0),
    .O_0(ShiftT_O_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = I_0; // @[ShiftTS.scala 40:36]
  assign O_2 = I_1; // @[ShiftTS.scala 40:36]
  assign O_3 = I_2; // @[ShiftTS.scala 40:36]
  assign O_4 = I_3; // @[ShiftTS.scala 40:36]
  assign O_5 = I_4; // @[ShiftTS.scala 40:36]
  assign O_6 = I_5; // @[ShiftTS.scala 40:36]
  assign O_7 = I_6; // @[ShiftTS.scala 40:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I_0 = I_7; // @[ShiftTS.scala 50:25]
endmodule
module SSeqTupleCreator(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  input  [15:0] I1,
  output [15:0] O_0,
  output [15:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I0_3,
  input  [15:0] I0_4,
  input  [15:0] I0_5,
  input  [15:0] I0_6,
  input  [15:0] I0_7,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_7_0,
  output [15:0] O_7_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  SSeqTupleCreator other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  SSeqTupleCreator other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  SSeqTupleCreator other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1)
  );
  SSeqTupleCreator other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1)
  );
  SSeqTupleCreator other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1)
  );
  SSeqTupleCreator other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I0_3,
  input  [15:0] I0_4,
  input  [15:0] I0_5,
  input  [15:0] I0_6,
  input  [15:0] I0_7,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_7_0,
  output [15:0] O_7_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I1,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  SSeqTupleAppender other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  SSeqTupleAppender other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  SSeqTupleAppender other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  SSeqTupleAppender other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  SSeqTupleAppender other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  SSeqTupleAppender other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_2_2 = other_ops_1_O_2; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_3_2 = other_ops_2_O_2; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_4_2 = other_ops_3_O_2; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_5_2 = other_ops_4_O_2; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_6_2 = other_ops_5_O_2; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_7_2 = other_ops_6_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_1_2 = op_O_1_2; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_2_2 = op_O_2_2; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_3_2 = op_O_3_2; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_4_2 = op_O_4_2; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_5_2 = op_O_5_2; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_6_2 = op_O_6_2; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_7_2 = op_O_7_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
endmodule
module PartitionS(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  input  [15:0] I_4_0,
  input  [15:0] I_4_1,
  input  [15:0] I_4_2,
  input  [15:0] I_5_0,
  input  [15:0] I_5_1,
  input  [15:0] I_5_2,
  input  [15:0] I_6_0,
  input  [15:0] I_6_1,
  input  [15:0] I_6_2,
  input  [15:0] I_7_0,
  input  [15:0] I_7_1,
  input  [15:0] I_7_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2 = I_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_3_0_2 = I_3_2; // @[Partition.scala 15:39]
  assign O_4_0_0 = I_4_0; // @[Partition.scala 15:39]
  assign O_4_0_1 = I_4_1; // @[Partition.scala 15:39]
  assign O_4_0_2 = I_4_2; // @[Partition.scala 15:39]
  assign O_5_0_0 = I_5_0; // @[Partition.scala 15:39]
  assign O_5_0_1 = I_5_1; // @[Partition.scala 15:39]
  assign O_5_0_2 = I_5_2; // @[Partition.scala 15:39]
  assign O_6_0_0 = I_6_0; // @[Partition.scala 15:39]
  assign O_6_0_1 = I_6_1; // @[Partition.scala 15:39]
  assign O_6_0_2 = I_6_2; // @[Partition.scala 15:39]
  assign O_7_0_0 = I_7_0; // @[Partition.scala 15:39]
  assign O_7_0_1 = I_7_1; // @[Partition.scala 15:39]
  assign O_7_0_2 = I_7_2; // @[Partition.scala 15:39]
endmodule
module MapT(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  input  [15:0] I_4_0,
  input  [15:0] I_4_1,
  input  [15:0] I_4_2,
  input  [15:0] I_5_0,
  input  [15:0] I_5_1,
  input  [15:0] I_5_2,
  input  [15:0] I_6_0,
  input  [15:0] I_6_1,
  input  [15:0] I_6_2,
  input  [15:0] I_7_0,
  input  [15:0] I_7_1,
  input  [15:0] I_7_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[MapT.scala 8:20]
  PartitionS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_1_2(op_I_1_2),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_2_2(op_I_2_2),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .I_3_2(op_I_3_2),
    .I_4_0(op_I_4_0),
    .I_4_1(op_I_4_1),
    .I_4_2(op_I_4_2),
    .I_5_0(op_I_5_0),
    .I_5_1(op_I_5_1),
    .I_5_2(op_I_5_2),
    .I_6_0(op_I_6_0),
    .I_6_1(op_I_6_1),
    .I_6_2(op_I_6_2),
    .I_7_0(op_I_7_0),
    .I_7_1(op_I_7_1),
    .I_7_2(op_I_7_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_1_2 = I_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2 = I_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
  assign op_I_3_2 = I_3_2; // @[MapT.scala 14:10]
  assign op_I_4_0 = I_4_0; // @[MapT.scala 14:10]
  assign op_I_4_1 = I_4_1; // @[MapT.scala 14:10]
  assign op_I_4_2 = I_4_2; // @[MapT.scala 14:10]
  assign op_I_5_0 = I_5_0; // @[MapT.scala 14:10]
  assign op_I_5_1 = I_5_1; // @[MapT.scala 14:10]
  assign op_I_5_2 = I_5_2; // @[MapT.scala 14:10]
  assign op_I_6_0 = I_6_0; // @[MapT.scala 14:10]
  assign op_I_6_1 = I_6_1; // @[MapT.scala 14:10]
  assign op_I_6_2 = I_6_2; // @[MapT.scala 14:10]
  assign op_I_7_0 = I_7_0; // @[MapT.scala 14:10]
  assign op_I_7_1 = I_7_1; // @[MapT.scala 14:10]
  assign op_I_7_2 = I_7_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  Remove1S other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  Remove1S other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  Remove1S other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  Remove1S other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  Remove1S other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  Remove1S other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_3_2 = other_ops_2_O_2; // @[MapS.scala 21:12]
  assign O_4_0 = other_ops_3_O_0; // @[MapS.scala 21:12]
  assign O_4_1 = other_ops_3_O_1; // @[MapS.scala 21:12]
  assign O_4_2 = other_ops_3_O_2; // @[MapS.scala 21:12]
  assign O_5_0 = other_ops_4_O_0; // @[MapS.scala 21:12]
  assign O_5_1 = other_ops_4_O_1; // @[MapS.scala 21:12]
  assign O_5_2 = other_ops_4_O_2; // @[MapS.scala 21:12]
  assign O_6_0 = other_ops_5_O_0; // @[MapS.scala 21:12]
  assign O_6_1 = other_ops_5_O_1; // @[MapS.scala 21:12]
  assign O_6_2 = other_ops_5_O_2; // @[MapS.scala 21:12]
  assign O_7_0 = other_ops_6_O_0; // @[MapS.scala 21:12]
  assign O_7_1 = other_ops_6_O_1; // @[MapS.scala 21:12]
  assign O_7_2 = other_ops_6_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
endmodule
module MapT_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_0_2 = op_O_0_2; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_1_2 = op_O_1_2; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_2_2 = op_O_2_2; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign O_3_2 = op_O_3_2; // @[MapT.scala 15:7]
  assign O_4_0 = op_O_4_0; // @[MapT.scala 15:7]
  assign O_4_1 = op_O_4_1; // @[MapT.scala 15:7]
  assign O_4_2 = op_O_4_2; // @[MapT.scala 15:7]
  assign O_5_0 = op_O_5_0; // @[MapT.scala 15:7]
  assign O_5_1 = op_O_5_1; // @[MapT.scala 15:7]
  assign O_5_2 = op_O_5_2; // @[MapT.scala 15:7]
  assign O_6_0 = op_O_6_0; // @[MapT.scala 15:7]
  assign O_6_1 = op_O_6_1; // @[MapT.scala 15:7]
  assign O_6_2 = op_O_6_2; // @[MapT.scala 15:7]
  assign O_7_0 = op_O_7_0; // @[MapT.scala 15:7]
  assign O_7_1 = op_O_7_1; // @[MapT.scala 15:7]
  assign O_7_2 = op_O_7_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_3_2,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_4_2,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_5_2,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_6_2,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I0_7_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I0_2(other_ops_2_I0_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I0_2(other_ops_3_I0_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I0_2(other_ops_4_I0_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I0_2(other_ops_5_I0_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I0_2(other_ops_6_I0_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2 = I0_3_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2 = I0_4_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2 = I0_5_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2 = I0_6_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2 = I0_7_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_3_2,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_4_2,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_5_2,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_6_2,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I0_7_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_0_2(op_I0_0_2),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_1_2(op_I0_1_2),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_2_2(op_I0_2_2),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_3_2(op_I0_3_2),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_4_2(op_I0_4_2),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_5_2(op_I0_5_2),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_6_2(op_I0_6_2),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_7_2(op_I0_7_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2 = I0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2 = I0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2 = I0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2 = I0_3_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_4_2 = I0_4_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_5_2 = I0_5_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_6_2 = I0_6_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_7_2 = I0_7_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0_0,
  input  [15:0] I0_0_0_1,
  input  [15:0] I0_0_0_2,
  input  [15:0] I0_0_1_0,
  input  [15:0] I0_0_1_1,
  input  [15:0] I0_0_1_2,
  input  [15:0] I0_1_0_0,
  input  [15:0] I0_1_0_1,
  input  [15:0] I0_1_0_2,
  input  [15:0] I0_1_1_0,
  input  [15:0] I0_1_1_1,
  input  [15:0] I0_1_1_2,
  input  [15:0] I0_2_0_0,
  input  [15:0] I0_2_0_1,
  input  [15:0] I0_2_0_2,
  input  [15:0] I0_2_1_0,
  input  [15:0] I0_2_1_1,
  input  [15:0] I0_2_1_2,
  input  [15:0] I0_3_0_0,
  input  [15:0] I0_3_0_1,
  input  [15:0] I0_3_0_2,
  input  [15:0] I0_3_1_0,
  input  [15:0] I0_3_1_1,
  input  [15:0] I0_3_1_2,
  input  [15:0] I0_4_0_0,
  input  [15:0] I0_4_0_1,
  input  [15:0] I0_4_0_2,
  input  [15:0] I0_4_1_0,
  input  [15:0] I0_4_1_1,
  input  [15:0] I0_4_1_2,
  input  [15:0] I0_5_0_0,
  input  [15:0] I0_5_0_1,
  input  [15:0] I0_5_0_2,
  input  [15:0] I0_5_1_0,
  input  [15:0] I0_5_1_1,
  input  [15:0] I0_5_1_2,
  input  [15:0] I0_6_0_0,
  input  [15:0] I0_6_0_1,
  input  [15:0] I0_6_0_2,
  input  [15:0] I0_6_1_0,
  input  [15:0] I0_6_1_1,
  input  [15:0] I0_6_1_2,
  input  [15:0] I0_7_0_0,
  input  [15:0] I0_7_0_1,
  input  [15:0] I0_7_0_2,
  input  [15:0] I0_7_1_0,
  input  [15:0] I0_7_1_1,
  input  [15:0] I0_7_1_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[Map2S.scala 24:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[Map2S.scala 24:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[Map2S.scala 24:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[Map2S.scala 24:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[Map2S.scala 24:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[Map2S.scala 24:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[Map2S.scala 24:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[Map2S.scala 24:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[Map2S.scala 24:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[Map2S.scala 24:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[Map2S.scala 24:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[Map2S.scala 24:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0_0,
  input  [15:0] I0_0_0_1,
  input  [15:0] I0_0_0_2,
  input  [15:0] I0_0_1_0,
  input  [15:0] I0_0_1_1,
  input  [15:0] I0_0_1_2,
  input  [15:0] I0_1_0_0,
  input  [15:0] I0_1_0_1,
  input  [15:0] I0_1_0_2,
  input  [15:0] I0_1_1_0,
  input  [15:0] I0_1_1_1,
  input  [15:0] I0_1_1_2,
  input  [15:0] I0_2_0_0,
  input  [15:0] I0_2_0_1,
  input  [15:0] I0_2_0_2,
  input  [15:0] I0_2_1_0,
  input  [15:0] I0_2_1_1,
  input  [15:0] I0_2_1_2,
  input  [15:0] I0_3_0_0,
  input  [15:0] I0_3_0_1,
  input  [15:0] I0_3_0_2,
  input  [15:0] I0_3_1_0,
  input  [15:0] I0_3_1_1,
  input  [15:0] I0_3_1_2,
  input  [15:0] I0_4_0_0,
  input  [15:0] I0_4_0_1,
  input  [15:0] I0_4_0_2,
  input  [15:0] I0_4_1_0,
  input  [15:0] I0_4_1_1,
  input  [15:0] I0_4_1_2,
  input  [15:0] I0_5_0_0,
  input  [15:0] I0_5_0_1,
  input  [15:0] I0_5_0_2,
  input  [15:0] I0_5_1_0,
  input  [15:0] I0_5_1_1,
  input  [15:0] I0_5_1_2,
  input  [15:0] I0_6_0_0,
  input  [15:0] I0_6_0_1,
  input  [15:0] I0_6_0_2,
  input  [15:0] I0_6_1_0,
  input  [15:0] I0_6_1_1,
  input  [15:0] I0_6_1_2,
  input  [15:0] I0_7_0_0,
  input  [15:0] I0_7_0_1,
  input  [15:0] I0_7_0_2,
  input  [15:0] I0_7_1_0,
  input  [15:0] I0_7_1_1,
  input  [15:0] I0_7_1_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2_2; // @[Map2T.scala 8:20]
  Map2S_7 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_4_1_0(op_I0_4_1_0),
    .I0_4_1_1(op_I0_4_1_1),
    .I0_4_1_2(op_I0_4_1_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_5_1_0(op_I0_5_1_0),
    .I0_5_1_1(op_I0_5_1_1),
    .I0_5_1_2(op_I0_5_1_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_6_1_0(op_I0_6_1_0),
    .I0_6_1_1(op_I0_6_1_1),
    .I0_6_1_2(op_I0_6_1_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_7_1_0(op_I0_7_1_0),
    .I0_7_1_1(op_I0_7_1_1),
    .I0_7_1_2(op_I0_7_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_2_0 = op_O_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_2_1 = op_O_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_2_2 = op_O_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_1_2_0 = op_O_1_2_0; // @[Map2T.scala 17:7]
  assign O_1_2_1 = op_O_1_2_1; // @[Map2T.scala 17:7]
  assign O_1_2_2 = op_O_1_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_2_2_0 = op_O_2_2_0; // @[Map2T.scala 17:7]
  assign O_2_2_1 = op_O_2_2_1; // @[Map2T.scala 17:7]
  assign O_2_2_2 = op_O_2_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_3_2_0 = op_O_3_2_0; // @[Map2T.scala 17:7]
  assign O_3_2_1 = op_O_3_2_1; // @[Map2T.scala 17:7]
  assign O_3_2_2 = op_O_3_2_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_4_2_0 = op_O_4_2_0; // @[Map2T.scala 17:7]
  assign O_4_2_1 = op_O_4_2_1; // @[Map2T.scala 17:7]
  assign O_4_2_2 = op_O_4_2_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_5_2_0 = op_O_5_2_0; // @[Map2T.scala 17:7]
  assign O_5_2_1 = op_O_5_2_1; // @[Map2T.scala 17:7]
  assign O_5_2_2 = op_O_5_2_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_6_2_0 = op_O_6_2_0; // @[Map2T.scala 17:7]
  assign O_6_2_1 = op_O_6_2_1; // @[Map2T.scala 17:7]
  assign O_6_2_2 = op_O_6_2_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_7_2_0 = op_O_7_2_0; // @[Map2T.scala 17:7]
  assign O_7_2_1 = op_O_7_2_1; // @[Map2T.scala 17:7]
  assign O_7_2_2 = op_O_7_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_1_0 = I0_4_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1_1 = I0_4_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_1_2 = I0_4_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_1_0 = I0_5_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1_1 = I0_5_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_1_2 = I0_5_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_1_0 = I0_6_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1_1 = I0_6_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_1_2 = I0_6_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_1_0 = I0_7_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1_1 = I0_7_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_1_2 = I0_7_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
endmodule
module PartitionS_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_0_2,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_0_0_1_2,
  output [15:0] O_0_0_2_0,
  output [15:0] O_0_0_2_1,
  output [15:0] O_0_0_2_2,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_0_2,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_1_0_1_2,
  output [15:0] O_1_0_2_0,
  output [15:0] O_1_0_2_1,
  output [15:0] O_1_0_2_2,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_0_2,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_2_0_1_2,
  output [15:0] O_2_0_2_0,
  output [15:0] O_2_0_2_1,
  output [15:0] O_2_0_2_2,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_0_2,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1,
  output [15:0] O_3_0_1_2,
  output [15:0] O_3_0_2_0,
  output [15:0] O_3_0_2_1,
  output [15:0] O_3_0_2_2,
  output [15:0] O_4_0_0_0,
  output [15:0] O_4_0_0_1,
  output [15:0] O_4_0_0_2,
  output [15:0] O_4_0_1_0,
  output [15:0] O_4_0_1_1,
  output [15:0] O_4_0_1_2,
  output [15:0] O_4_0_2_0,
  output [15:0] O_4_0_2_1,
  output [15:0] O_4_0_2_2,
  output [15:0] O_5_0_0_0,
  output [15:0] O_5_0_0_1,
  output [15:0] O_5_0_0_2,
  output [15:0] O_5_0_1_0,
  output [15:0] O_5_0_1_1,
  output [15:0] O_5_0_1_2,
  output [15:0] O_5_0_2_0,
  output [15:0] O_5_0_2_1,
  output [15:0] O_5_0_2_2,
  output [15:0] O_6_0_0_0,
  output [15:0] O_6_0_0_1,
  output [15:0] O_6_0_0_2,
  output [15:0] O_6_0_1_0,
  output [15:0] O_6_0_1_1,
  output [15:0] O_6_0_1_2,
  output [15:0] O_6_0_2_0,
  output [15:0] O_6_0_2_1,
  output [15:0] O_6_0_2_2,
  output [15:0] O_7_0_0_0,
  output [15:0] O_7_0_0_1,
  output [15:0] O_7_0_0_2,
  output [15:0] O_7_0_1_0,
  output [15:0] O_7_0_1_1,
  output [15:0] O_7_0_1_2,
  output [15:0] O_7_0_2_0,
  output [15:0] O_7_0_2_1,
  output [15:0] O_7_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_0_2 = I_2_0_2; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_2_0_1_2 = I_2_1_2; // @[Partition.scala 15:39]
  assign O_2_0_2_0 = I_2_2_0; // @[Partition.scala 15:39]
  assign O_2_0_2_1 = I_2_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2_2 = I_2_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_0_2 = I_3_0_2; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_3_0_1_2 = I_3_1_2; // @[Partition.scala 15:39]
  assign O_3_0_2_0 = I_3_2_0; // @[Partition.scala 15:39]
  assign O_3_0_2_1 = I_3_2_1; // @[Partition.scala 15:39]
  assign O_3_0_2_2 = I_3_2_2; // @[Partition.scala 15:39]
  assign O_4_0_0_0 = I_4_0_0; // @[Partition.scala 15:39]
  assign O_4_0_0_1 = I_4_0_1; // @[Partition.scala 15:39]
  assign O_4_0_0_2 = I_4_0_2; // @[Partition.scala 15:39]
  assign O_4_0_1_0 = I_4_1_0; // @[Partition.scala 15:39]
  assign O_4_0_1_1 = I_4_1_1; // @[Partition.scala 15:39]
  assign O_4_0_1_2 = I_4_1_2; // @[Partition.scala 15:39]
  assign O_4_0_2_0 = I_4_2_0; // @[Partition.scala 15:39]
  assign O_4_0_2_1 = I_4_2_1; // @[Partition.scala 15:39]
  assign O_4_0_2_2 = I_4_2_2; // @[Partition.scala 15:39]
  assign O_5_0_0_0 = I_5_0_0; // @[Partition.scala 15:39]
  assign O_5_0_0_1 = I_5_0_1; // @[Partition.scala 15:39]
  assign O_5_0_0_2 = I_5_0_2; // @[Partition.scala 15:39]
  assign O_5_0_1_0 = I_5_1_0; // @[Partition.scala 15:39]
  assign O_5_0_1_1 = I_5_1_1; // @[Partition.scala 15:39]
  assign O_5_0_1_2 = I_5_1_2; // @[Partition.scala 15:39]
  assign O_5_0_2_0 = I_5_2_0; // @[Partition.scala 15:39]
  assign O_5_0_2_1 = I_5_2_1; // @[Partition.scala 15:39]
  assign O_5_0_2_2 = I_5_2_2; // @[Partition.scala 15:39]
  assign O_6_0_0_0 = I_6_0_0; // @[Partition.scala 15:39]
  assign O_6_0_0_1 = I_6_0_1; // @[Partition.scala 15:39]
  assign O_6_0_0_2 = I_6_0_2; // @[Partition.scala 15:39]
  assign O_6_0_1_0 = I_6_1_0; // @[Partition.scala 15:39]
  assign O_6_0_1_1 = I_6_1_1; // @[Partition.scala 15:39]
  assign O_6_0_1_2 = I_6_1_2; // @[Partition.scala 15:39]
  assign O_6_0_2_0 = I_6_2_0; // @[Partition.scala 15:39]
  assign O_6_0_2_1 = I_6_2_1; // @[Partition.scala 15:39]
  assign O_6_0_2_2 = I_6_2_2; // @[Partition.scala 15:39]
  assign O_7_0_0_0 = I_7_0_0; // @[Partition.scala 15:39]
  assign O_7_0_0_1 = I_7_0_1; // @[Partition.scala 15:39]
  assign O_7_0_0_2 = I_7_0_2; // @[Partition.scala 15:39]
  assign O_7_0_1_0 = I_7_1_0; // @[Partition.scala 15:39]
  assign O_7_0_1_1 = I_7_1_1; // @[Partition.scala 15:39]
  assign O_7_0_1_2 = I_7_1_2; // @[Partition.scala 15:39]
  assign O_7_0_2_0 = I_7_2_0; // @[Partition.scala 15:39]
  assign O_7_0_2_1 = I_7_2_1; // @[Partition.scala 15:39]
  assign O_7_0_2_2 = I_7_2_2; // @[Partition.scala 15:39]
endmodule
module MapT_6(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_0_2,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_0_0_1_2,
  output [15:0] O_0_0_2_0,
  output [15:0] O_0_0_2_1,
  output [15:0] O_0_0_2_2,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_0_2,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_1_0_1_2,
  output [15:0] O_1_0_2_0,
  output [15:0] O_1_0_2_1,
  output [15:0] O_1_0_2_2,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_0_2,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_2_0_1_2,
  output [15:0] O_2_0_2_0,
  output [15:0] O_2_0_2_1,
  output [15:0] O_2_0_2_2,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_0_2,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1,
  output [15:0] O_3_0_1_2,
  output [15:0] O_3_0_2_0,
  output [15:0] O_3_0_2_1,
  output [15:0] O_3_0_2_2,
  output [15:0] O_4_0_0_0,
  output [15:0] O_4_0_0_1,
  output [15:0] O_4_0_0_2,
  output [15:0] O_4_0_1_0,
  output [15:0] O_4_0_1_1,
  output [15:0] O_4_0_1_2,
  output [15:0] O_4_0_2_0,
  output [15:0] O_4_0_2_1,
  output [15:0] O_4_0_2_2,
  output [15:0] O_5_0_0_0,
  output [15:0] O_5_0_0_1,
  output [15:0] O_5_0_0_2,
  output [15:0] O_5_0_1_0,
  output [15:0] O_5_0_1_1,
  output [15:0] O_5_0_1_2,
  output [15:0] O_5_0_2_0,
  output [15:0] O_5_0_2_1,
  output [15:0] O_5_0_2_2,
  output [15:0] O_6_0_0_0,
  output [15:0] O_6_0_0_1,
  output [15:0] O_6_0_0_2,
  output [15:0] O_6_0_1_0,
  output [15:0] O_6_0_1_1,
  output [15:0] O_6_0_1_2,
  output [15:0] O_6_0_2_0,
  output [15:0] O_6_0_2_1,
  output [15:0] O_6_0_2_2,
  output [15:0] O_7_0_0_0,
  output [15:0] O_7_0_0_1,
  output [15:0] O_7_0_0_2,
  output [15:0] O_7_0_1_0,
  output [15:0] O_7_0_1_1,
  output [15:0] O_7_0_1_2,
  output [15:0] O_7_0_2_0,
  output [15:0] O_7_0_2_1,
  output [15:0] O_7_0_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2_2; // @[MapT.scala 8:20]
  PartitionS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_4_0_2_0(op_O_4_0_2_0),
    .O_4_0_2_1(op_O_4_0_2_1),
    .O_4_0_2_2(op_O_4_0_2_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_5_0_2_0(op_O_5_0_2_0),
    .O_5_0_2_1(op_O_5_0_2_1),
    .O_5_0_2_2(op_O_5_0_2_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_6_0_2_0(op_O_6_0_2_0),
    .O_6_0_2_1(op_O_6_0_2_1),
    .O_6_0_2_2(op_O_6_0_2_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_7_0_2_0(op_O_7_0_2_0),
    .O_7_0_2_1(op_O_7_0_2_1),
    .O_7_0_2_2(op_O_7_0_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[MapT.scala 15:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[MapT.scala 15:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[MapT.scala 15:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[MapT.scala 15:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[MapT.scala 15:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[MapT.scala 15:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[MapT.scala 15:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[MapT.scala 15:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[MapT.scala 15:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[MapT.scala 15:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[MapT.scala 15:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[MapT.scala 15:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[MapT.scala 15:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[MapT.scala 15:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[MapT.scala 15:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[MapT.scala 15:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[MapT.scala 15:7]
  assign O_4_0_2_0 = op_O_4_0_2_0; // @[MapT.scala 15:7]
  assign O_4_0_2_1 = op_O_4_0_2_1; // @[MapT.scala 15:7]
  assign O_4_0_2_2 = op_O_4_0_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[MapT.scala 15:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[MapT.scala 15:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[MapT.scala 15:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[MapT.scala 15:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[MapT.scala 15:7]
  assign O_5_0_2_0 = op_O_5_0_2_0; // @[MapT.scala 15:7]
  assign O_5_0_2_1 = op_O_5_0_2_1; // @[MapT.scala 15:7]
  assign O_5_0_2_2 = op_O_5_0_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[MapT.scala 15:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[MapT.scala 15:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[MapT.scala 15:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[MapT.scala 15:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[MapT.scala 15:7]
  assign O_6_0_2_0 = op_O_6_0_2_0; // @[MapT.scala 15:7]
  assign O_6_0_2_1 = op_O_6_0_2_1; // @[MapT.scala 15:7]
  assign O_6_0_2_2 = op_O_6_0_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[MapT.scala 15:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[MapT.scala 15:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[MapT.scala 15:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[MapT.scala 15:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[MapT.scala 15:7]
  assign O_7_0_2_0 = op_O_7_0_2_0; // @[MapT.scala 15:7]
  assign O_7_0_2_1 = op_O_7_0_2_1; // @[MapT.scala 15:7]
  assign O_7_0_2_2 = op_O_7_0_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_0_2,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_0_0_1_2,
  input  [15:0] I_0_0_2_0,
  input  [15:0] I_0_0_2_1,
  input  [15:0] I_0_0_2_2,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_0_2,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_1_0_1_2,
  input  [15:0] I_1_0_2_0,
  input  [15:0] I_1_0_2_1,
  input  [15:0] I_1_0_2_2,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_0_2,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_2_0_1_2,
  input  [15:0] I_2_0_2_0,
  input  [15:0] I_2_0_2_1,
  input  [15:0] I_2_0_2_2,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_0_2,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  input  [15:0] I_3_0_1_2,
  input  [15:0] I_3_0_2_0,
  input  [15:0] I_3_0_2_1,
  input  [15:0] I_3_0_2_2,
  input  [15:0] I_4_0_0_0,
  input  [15:0] I_4_0_0_1,
  input  [15:0] I_4_0_0_2,
  input  [15:0] I_4_0_1_0,
  input  [15:0] I_4_0_1_1,
  input  [15:0] I_4_0_1_2,
  input  [15:0] I_4_0_2_0,
  input  [15:0] I_4_0_2_1,
  input  [15:0] I_4_0_2_2,
  input  [15:0] I_5_0_0_0,
  input  [15:0] I_5_0_0_1,
  input  [15:0] I_5_0_0_2,
  input  [15:0] I_5_0_1_0,
  input  [15:0] I_5_0_1_1,
  input  [15:0] I_5_0_1_2,
  input  [15:0] I_5_0_2_0,
  input  [15:0] I_5_0_2_1,
  input  [15:0] I_5_0_2_2,
  input  [15:0] I_6_0_0_0,
  input  [15:0] I_6_0_0_1,
  input  [15:0] I_6_0_0_2,
  input  [15:0] I_6_0_1_0,
  input  [15:0] I_6_0_1_1,
  input  [15:0] I_6_0_1_2,
  input  [15:0] I_6_0_2_0,
  input  [15:0] I_6_0_2_1,
  input  [15:0] I_6_0_2_2,
  input  [15:0] I_7_0_0_0,
  input  [15:0] I_7_0_0_1,
  input  [15:0] I_7_0_0_2,
  input  [15:0] I_7_0_1_0,
  input  [15:0] I_7_0_1_1,
  input  [15:0] I_7_0_1_2,
  input  [15:0] I_7_0_2_0,
  input  [15:0] I_7_0_2_1,
  input  [15:0] I_7_0_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_0_2,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_0_0_1_2,
  input  [15:0] I_0_0_2_0,
  input  [15:0] I_0_0_2_1,
  input  [15:0] I_0_0_2_2,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_0_2,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_1_0_1_2,
  input  [15:0] I_1_0_2_0,
  input  [15:0] I_1_0_2_1,
  input  [15:0] I_1_0_2_2,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_0_2,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_2_0_1_2,
  input  [15:0] I_2_0_2_0,
  input  [15:0] I_2_0_2_1,
  input  [15:0] I_2_0_2_2,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_0_2,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  input  [15:0] I_3_0_1_2,
  input  [15:0] I_3_0_2_0,
  input  [15:0] I_3_0_2_1,
  input  [15:0] I_3_0_2_2,
  input  [15:0] I_4_0_0_0,
  input  [15:0] I_4_0_0_1,
  input  [15:0] I_4_0_0_2,
  input  [15:0] I_4_0_1_0,
  input  [15:0] I_4_0_1_1,
  input  [15:0] I_4_0_1_2,
  input  [15:0] I_4_0_2_0,
  input  [15:0] I_4_0_2_1,
  input  [15:0] I_4_0_2_2,
  input  [15:0] I_5_0_0_0,
  input  [15:0] I_5_0_0_1,
  input  [15:0] I_5_0_0_2,
  input  [15:0] I_5_0_1_0,
  input  [15:0] I_5_0_1_1,
  input  [15:0] I_5_0_1_2,
  input  [15:0] I_5_0_2_0,
  input  [15:0] I_5_0_2_1,
  input  [15:0] I_5_0_2_2,
  input  [15:0] I_6_0_0_0,
  input  [15:0] I_6_0_0_1,
  input  [15:0] I_6_0_0_2,
  input  [15:0] I_6_0_1_0,
  input  [15:0] I_6_0_1_1,
  input  [15:0] I_6_0_1_2,
  input  [15:0] I_6_0_2_0,
  input  [15:0] I_6_0_2_1,
  input  [15:0] I_6_0_2_2,
  input  [15:0] I_7_0_0_0,
  input  [15:0] I_7_0_0_1,
  input  [15:0] I_7_0_0_2,
  input  [15:0] I_7_0_1_0,
  input  [15:0] I_7_0_1_1,
  input  [15:0] I_7_0_1_2,
  input  [15:0] I_7_0_2_0,
  input  [15:0] I_7_0_2_1,
  input  [15:0] I_7_0_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_4_0_1_2(op_I_4_0_1_2),
    .I_4_0_2_0(op_I_4_0_2_0),
    .I_4_0_2_1(op_I_4_0_2_1),
    .I_4_0_2_2(op_I_4_0_2_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_5_0_1_2(op_I_5_0_1_2),
    .I_5_0_2_0(op_I_5_0_2_0),
    .I_5_0_2_1(op_I_5_0_2_1),
    .I_5_0_2_2(op_I_5_0_2_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_6_0_1_2(op_I_6_0_1_2),
    .I_6_0_2_0(op_I_6_0_2_0),
    .I_6_0_2_1(op_I_6_0_2_1),
    .I_6_0_2_2(op_I_6_0_2_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_7_0_1_2(op_I_7_0_1_2),
    .I_7_0_2_0(op_I_7_0_2_0),
    .I_7_0_2_1(op_I_7_0_2_1),
    .I_7_0_2_2(op_I_7_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_4_1_2 = op_O_4_1_2; // @[MapT.scala 15:7]
  assign O_4_2_0 = op_O_4_2_0; // @[MapT.scala 15:7]
  assign O_4_2_1 = op_O_4_2_1; // @[MapT.scala 15:7]
  assign O_4_2_2 = op_O_4_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_5_1_2 = op_O_5_1_2; // @[MapT.scala 15:7]
  assign O_5_2_0 = op_O_5_2_0; // @[MapT.scala 15:7]
  assign O_5_2_1 = op_O_5_2_1; // @[MapT.scala 15:7]
  assign O_5_2_2 = op_O_5_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_6_1_2 = op_O_6_1_2; // @[MapT.scala 15:7]
  assign O_6_2_0 = op_O_6_2_0; // @[MapT.scala 15:7]
  assign O_6_2_1 = op_O_6_2_1; // @[MapT.scala 15:7]
  assign O_6_2_2 = op_O_6_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_7_1_2 = op_O_7_1_2; // @[MapT.scala 15:7]
  assign O_7_2_0 = op_O_7_2_0; // @[MapT.scala 15:7]
  assign O_7_2_1 = op_O_7_2_1; // @[MapT.scala 15:7]
  assign O_7_2_2 = op_O_7_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_2 = I_4_0_1_2; // @[MapT.scala 14:10]
  assign op_I_4_0_2_0 = I_4_0_2_0; // @[MapT.scala 14:10]
  assign op_I_4_0_2_1 = I_4_0_2_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2_2 = I_4_0_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_2 = I_5_0_1_2; // @[MapT.scala 14:10]
  assign op_I_5_0_2_0 = I_5_0_2_0; // @[MapT.scala 14:10]
  assign op_I_5_0_2_1 = I_5_0_2_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2_2 = I_5_0_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_2 = I_6_0_1_2; // @[MapT.scala 14:10]
  assign op_I_6_0_2_0 = I_6_0_2_0; // @[MapT.scala 14:10]
  assign op_I_6_0_2_1 = I_6_0_2_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2_2 = I_6_0_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_2 = I_7_0_1_2; // @[MapT.scala 14:10]
  assign op_I_7_0_2_0 = I_7_0_2_0; // @[MapT.scala 14:10]
  assign op_I_7_0_2_1 = I_7_0_2_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2_2 = I_7_0_2_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  input  [15:0] I1,
  output [15:0] O_t0b,
  output [15:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_t0b,
  output [15:0] O_0_t1b,
  output [15:0] O_1_t0b,
  output [15:0] O_1_t1b,
  output [15:0] O_2_t0b,
  output [15:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_9(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  output [15:0] O_0_0_t0b,
  output [15:0] O_0_0_t1b,
  output [15:0] O_0_1_t0b,
  output [15:0] O_0_1_t1b,
  output [15:0] O_0_2_t0b,
  output [15:0] O_0_2_t1b,
  output [15:0] O_1_0_t0b,
  output [15:0] O_1_0_t1b,
  output [15:0] O_1_1_t0b,
  output [15:0] O_1_1_t1b,
  output [15:0] O_1_2_t0b,
  output [15:0] O_1_2_t1b,
  output [15:0] O_2_0_t0b,
  output [15:0] O_2_0_t1b,
  output [15:0] O_2_1_t0b,
  output [15:0] O_2_1_t1b,
  output [15:0] O_2_2_t0b,
  output [15:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_8 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_8 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_8 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 16'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 16'h2; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 16'h1; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 16'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 16'h4; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 16'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 16'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 16'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 16'h1; // @[Map2S.scala 23:43]
endmodule
module Mul(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_t0b,
  input  [15:0] I_t1b,
  output [15:0] O
);
  wire [15:0] BlackBoxMulUInt16_I0; // @[Arithmetic.scala 180:27]
  wire [15:0] BlackBoxMulUInt16_I1; // @[Arithmetic.scala 180:27]
  wire [31:0] BlackBoxMulUInt16_O; // @[Arithmetic.scala 180:27]
  wire  BlackBoxMulUInt16_clock; // @[Arithmetic.scala 180:27]
  reg  _T_1; // @[Arithmetic.scala 217:42]
  reg [31:0] _RAND_0;
  reg  _T_2; // @[Arithmetic.scala 217:34]
  reg [31:0] _RAND_1;
  reg  _T_3; // @[Arithmetic.scala 217:26]
  reg [31:0] _RAND_2;
  BlackBoxMulUInt16 BlackBoxMulUInt16 ( // @[Arithmetic.scala 180:27]
    .I0(BlackBoxMulUInt16_I0),
    .I1(BlackBoxMulUInt16_I1),
    .O(BlackBoxMulUInt16_O),
    .clock(BlackBoxMulUInt16_clock)
  );
  assign valid_down = _T_3; // @[Arithmetic.scala 217:16]
  assign O = BlackBoxMulUInt16_O[15:0]; // @[Arithmetic.scala 183:7]
  assign BlackBoxMulUInt16_I0 = I_t0b; // @[Arithmetic.scala 181:21]
  assign BlackBoxMulUInt16_I1 = I_t1b; // @[Arithmetic.scala 182:21]
  assign BlackBoxMulUInt16_clock = clock; // @[Arithmetic.scala 184:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _T_1;
    end
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= _T_2;
    end
  end
endmodule
module MapS_4(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_t0b,
  input  [15:0] I_0_t1b,
  input  [15:0] I_1_t0b,
  input  [15:0] I_1_t1b,
  input  [15:0] I_2_t0b,
  input  [15:0] I_2_t1b,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  Mul fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  Mul other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  Mul other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_5(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_t0b,
  input  [15:0] I_0_0_t1b,
  input  [15:0] I_0_1_t0b,
  input  [15:0] I_0_1_t1b,
  input  [15:0] I_0_2_t0b,
  input  [15:0] I_0_2_t1b,
  input  [15:0] I_1_0_t0b,
  input  [15:0] I_1_0_t1b,
  input  [15:0] I_1_1_t0b,
  input  [15:0] I_1_1_t1b,
  input  [15:0] I_1_2_t0b,
  input  [15:0] I_1_2_t1b,
  input  [15:0] I_2_0_t0b,
  input  [15:0] I_2_0_t1b,
  input  [15:0] I_2_1_t0b,
  input  [15:0] I_2_1_t1b,
  input  [15:0] I_2_2_t0b,
  input  [15:0] I_2_2_t1b,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_4 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_4 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_4 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [15:0] I_t0b,
  input  [15:0] I_t1b,
  output [15:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  output [15:0] O_0
);
  wire [15:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [15:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [15:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [15:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [15:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = _T_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module MapS_6(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0,
  output [15:0] O_1_0,
  output [15:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [15:0] I_0_t0b,
  input  [15:0] I_0_t1b,
  output [15:0] O_0
);
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [15:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [15:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_1_0,
  input  [15:0] I_2_0,
  output [15:0] O_0_0
);
  wire [15:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [15:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [15:0] _T_1_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [15:0] _T_2_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [15:0] _T_3_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = _T_2_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = _T_3_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = _T_1_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1_0 <= I_0_0;
    _T_2_0 <= I_1_0;
    _T_3_0 <= I_2_0;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [3:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [3:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 4'h8; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 4'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 4'h8; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 4'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  output [15:0] O_t0b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
endmodule
module Map2S_10(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  output [15:0] O_0_t0b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  AtomTuple_1 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .O_t0b(fst_op_O_t0b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
endmodule
module Map2S_11(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  output [15:0] O_0_0_t0b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  Map2S_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .O_0_t0b(fst_op_O_0_t0b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
endmodule
module Div(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_t0b,
  output [15:0] O
);
  wire [15:0] BlackBoxMulUInt16_I0; // @[Arithmetic.scala 349:27]
  wire [15:0] BlackBoxMulUInt16_I1; // @[Arithmetic.scala 349:27]
  wire [31:0] BlackBoxMulUInt16_O; // @[Arithmetic.scala 349:27]
  wire  BlackBoxMulUInt16_clock; // @[Arithmetic.scala 349:27]
  reg  _T_3; // @[Arithmetic.scala 370:42]
  reg [31:0] _RAND_0;
  reg  _T_4; // @[Arithmetic.scala 370:34]
  reg [31:0] _RAND_1;
  reg  _T_5; // @[Arithmetic.scala 370:26]
  reg [31:0] _RAND_2;
  BlackBoxMulUInt16 BlackBoxMulUInt16 ( // @[Arithmetic.scala 349:27]
    .I0(BlackBoxMulUInt16_I0),
    .I1(BlackBoxMulUInt16_I1),
    .O(BlackBoxMulUInt16_O),
    .clock(BlackBoxMulUInt16_clock)
  );
  assign valid_down = _T_5; // @[Arithmetic.scala 370:16]
  assign O = BlackBoxMulUInt16_O[22:7]; // @[Arithmetic.scala 352:7]
  assign BlackBoxMulUInt16_I0 = I_t0b; // @[Arithmetic.scala 350:21]
  assign BlackBoxMulUInt16_I1 = 16'h8; // @[Arithmetic.scala 351:21]
  assign BlackBoxMulUInt16_clock = clock; // @[Arithmetic.scala 353:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_5 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= valid_up;
    end
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= _T_3;
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= _T_4;
    end
  end
endmodule
module MapS_7(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_t0b,
  output [15:0] O_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O; // @[MapS.scala 9:22]
  Div fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
endmodule
module MapS_8(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_t0b,
  output [15:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n110_valid_up; // @[Top.scala 18:22]
  wire  n110_valid_down; // @[Top.scala 18:22]
  wire [15:0] n110_I0_0_0; // @[Top.scala 18:22]
  wire [15:0] n110_I0_0_1; // @[Top.scala 18:22]
  wire [15:0] n110_I0_0_2; // @[Top.scala 18:22]
  wire [15:0] n110_I0_1_0; // @[Top.scala 18:22]
  wire [15:0] n110_I0_1_1; // @[Top.scala 18:22]
  wire [15:0] n110_I0_1_2; // @[Top.scala 18:22]
  wire [15:0] n110_I0_2_0; // @[Top.scala 18:22]
  wire [15:0] n110_I0_2_1; // @[Top.scala 18:22]
  wire [15:0] n110_I0_2_2; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_0_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_1_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_2_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_2_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_0_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_1_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_2_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_2_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_0_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_1_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_2_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_2_t1b; // @[Top.scala 18:22]
  wire  n121_clock; // @[Top.scala 22:22]
  wire  n121_reset; // @[Top.scala 22:22]
  wire  n121_valid_up; // @[Top.scala 22:22]
  wire  n121_valid_down; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_0_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_1_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_2_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_0_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_1_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_2_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_0_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_1_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_2_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_O_0_0; // @[Top.scala 22:22]
  wire [15:0] n121_O_0_1; // @[Top.scala 22:22]
  wire [15:0] n121_O_0_2; // @[Top.scala 22:22]
  wire [15:0] n121_O_1_0; // @[Top.scala 22:22]
  wire [15:0] n121_O_1_1; // @[Top.scala 22:22]
  wire [15:0] n121_O_1_2; // @[Top.scala 22:22]
  wire [15:0] n121_O_2_0; // @[Top.scala 22:22]
  wire [15:0] n121_O_2_1; // @[Top.scala 22:22]
  wire [15:0] n121_O_2_2; // @[Top.scala 22:22]
  wire  n126_clock; // @[Top.scala 25:22]
  wire  n126_reset; // @[Top.scala 25:22]
  wire  n126_valid_up; // @[Top.scala 25:22]
  wire  n126_valid_down; // @[Top.scala 25:22]
  wire [15:0] n126_I_0_0; // @[Top.scala 25:22]
  wire [15:0] n126_I_0_1; // @[Top.scala 25:22]
  wire [15:0] n126_I_0_2; // @[Top.scala 25:22]
  wire [15:0] n126_I_1_0; // @[Top.scala 25:22]
  wire [15:0] n126_I_1_1; // @[Top.scala 25:22]
  wire [15:0] n126_I_1_2; // @[Top.scala 25:22]
  wire [15:0] n126_I_2_0; // @[Top.scala 25:22]
  wire [15:0] n126_I_2_1; // @[Top.scala 25:22]
  wire [15:0] n126_I_2_2; // @[Top.scala 25:22]
  wire [15:0] n126_O_0_0; // @[Top.scala 25:22]
  wire [15:0] n126_O_1_0; // @[Top.scala 25:22]
  wire [15:0] n126_O_2_0; // @[Top.scala 25:22]
  wire  n131_clock; // @[Top.scala 28:22]
  wire  n131_reset; // @[Top.scala 28:22]
  wire  n131_valid_up; // @[Top.scala 28:22]
  wire  n131_valid_down; // @[Top.scala 28:22]
  wire [15:0] n131_I_0_0; // @[Top.scala 28:22]
  wire [15:0] n131_I_1_0; // @[Top.scala 28:22]
  wire [15:0] n131_I_2_0; // @[Top.scala 28:22]
  wire [15:0] n131_O_0_0; // @[Top.scala 28:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n134_valid_up; // @[Top.scala 32:22]
  wire  n134_valid_down; // @[Top.scala 32:22]
  wire [15:0] n134_I0_0_0; // @[Top.scala 32:22]
  wire [15:0] n134_O_0_0_t0b; // @[Top.scala 32:22]
  wire  n145_clock; // @[Top.scala 36:22]
  wire  n145_reset; // @[Top.scala 36:22]
  wire  n145_valid_up; // @[Top.scala 36:22]
  wire  n145_valid_down; // @[Top.scala 36:22]
  wire [15:0] n145_I_0_0_t0b; // @[Top.scala 36:22]
  wire [15:0] n145_O_0_0; // @[Top.scala 36:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_9 n110 ( // @[Top.scala 18:22]
    .valid_up(n110_valid_up),
    .valid_down(n110_valid_down),
    .I0_0_0(n110_I0_0_0),
    .I0_0_1(n110_I0_0_1),
    .I0_0_2(n110_I0_0_2),
    .I0_1_0(n110_I0_1_0),
    .I0_1_1(n110_I0_1_1),
    .I0_1_2(n110_I0_1_2),
    .I0_2_0(n110_I0_2_0),
    .I0_2_1(n110_I0_2_1),
    .I0_2_2(n110_I0_2_2),
    .O_0_0_t0b(n110_O_0_0_t0b),
    .O_0_0_t1b(n110_O_0_0_t1b),
    .O_0_1_t0b(n110_O_0_1_t0b),
    .O_0_1_t1b(n110_O_0_1_t1b),
    .O_0_2_t0b(n110_O_0_2_t0b),
    .O_0_2_t1b(n110_O_0_2_t1b),
    .O_1_0_t0b(n110_O_1_0_t0b),
    .O_1_0_t1b(n110_O_1_0_t1b),
    .O_1_1_t0b(n110_O_1_1_t0b),
    .O_1_1_t1b(n110_O_1_1_t1b),
    .O_1_2_t0b(n110_O_1_2_t0b),
    .O_1_2_t1b(n110_O_1_2_t1b),
    .O_2_0_t0b(n110_O_2_0_t0b),
    .O_2_0_t1b(n110_O_2_0_t1b),
    .O_2_1_t0b(n110_O_2_1_t0b),
    .O_2_1_t1b(n110_O_2_1_t1b),
    .O_2_2_t0b(n110_O_2_2_t0b),
    .O_2_2_t1b(n110_O_2_2_t1b)
  );
  MapS_5 n121 ( // @[Top.scala 22:22]
    .clock(n121_clock),
    .reset(n121_reset),
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I_0_0_t0b(n121_I_0_0_t0b),
    .I_0_0_t1b(n121_I_0_0_t1b),
    .I_0_1_t0b(n121_I_0_1_t0b),
    .I_0_1_t1b(n121_I_0_1_t1b),
    .I_0_2_t0b(n121_I_0_2_t0b),
    .I_0_2_t1b(n121_I_0_2_t1b),
    .I_1_0_t0b(n121_I_1_0_t0b),
    .I_1_0_t1b(n121_I_1_0_t1b),
    .I_1_1_t0b(n121_I_1_1_t0b),
    .I_1_1_t1b(n121_I_1_1_t1b),
    .I_1_2_t0b(n121_I_1_2_t0b),
    .I_1_2_t1b(n121_I_1_2_t1b),
    .I_2_0_t0b(n121_I_2_0_t0b),
    .I_2_0_t1b(n121_I_2_0_t1b),
    .I_2_1_t0b(n121_I_2_1_t0b),
    .I_2_1_t1b(n121_I_2_1_t1b),
    .I_2_2_t0b(n121_I_2_2_t0b),
    .I_2_2_t1b(n121_I_2_2_t1b),
    .O_0_0(n121_O_0_0),
    .O_0_1(n121_O_0_1),
    .O_0_2(n121_O_0_2),
    .O_1_0(n121_O_1_0),
    .O_1_1(n121_O_1_1),
    .O_1_2(n121_O_1_2),
    .O_2_0(n121_O_2_0),
    .O_2_1(n121_O_2_1),
    .O_2_2(n121_O_2_2)
  );
  MapS_6 n126 ( // @[Top.scala 25:22]
    .clock(n126_clock),
    .reset(n126_reset),
    .valid_up(n126_valid_up),
    .valid_down(n126_valid_down),
    .I_0_0(n126_I_0_0),
    .I_0_1(n126_I_0_1),
    .I_0_2(n126_I_0_2),
    .I_1_0(n126_I_1_0),
    .I_1_1(n126_I_1_1),
    .I_1_2(n126_I_1_2),
    .I_2_0(n126_I_2_0),
    .I_2_1(n126_I_2_1),
    .I_2_2(n126_I_2_2),
    .O_0_0(n126_O_0_0),
    .O_1_0(n126_O_1_0),
    .O_2_0(n126_O_2_0)
  );
  ReduceS_1 n131 ( // @[Top.scala 28:22]
    .clock(n131_clock),
    .reset(n131_reset),
    .valid_up(n131_valid_up),
    .valid_down(n131_valid_down),
    .I_0_0(n131_I_0_0),
    .I_1_0(n131_I_1_0),
    .I_2_0(n131_I_2_0),
    .O_0_0(n131_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n134 ( // @[Top.scala 32:22]
    .valid_up(n134_valid_up),
    .valid_down(n134_valid_down),
    .I0_0_0(n134_I0_0_0),
    .O_0_0_t0b(n134_O_0_0_t0b)
  );
  MapS_8 n145 ( // @[Top.scala 36:22]
    .clock(n145_clock),
    .reset(n145_reset),
    .valid_up(n145_valid_up),
    .valid_down(n145_valid_down),
    .I_0_0_t0b(n145_I_0_0_t0b),
    .O_0_0(n145_O_0_0)
  );
  assign valid_down = n145_valid_down; // @[Top.scala 40:16]
  assign O_0_0 = n145_O_0_0; // @[Top.scala 39:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n110_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 21:19]
  assign n110_I0_0_0 = I_0_0; // @[Top.scala 19:13]
  assign n110_I0_0_1 = I_0_1; // @[Top.scala 19:13]
  assign n110_I0_0_2 = I_0_2; // @[Top.scala 19:13]
  assign n110_I0_1_0 = I_1_0; // @[Top.scala 19:13]
  assign n110_I0_1_1 = I_1_1; // @[Top.scala 19:13]
  assign n110_I0_1_2 = I_1_2; // @[Top.scala 19:13]
  assign n110_I0_2_0 = I_2_0; // @[Top.scala 19:13]
  assign n110_I0_2_1 = I_2_1; // @[Top.scala 19:13]
  assign n110_I0_2_2 = I_2_2; // @[Top.scala 19:13]
  assign n121_clock = clock;
  assign n121_reset = reset;
  assign n121_valid_up = n110_valid_down; // @[Top.scala 24:19]
  assign n121_I_0_0_t0b = n110_O_0_0_t0b; // @[Top.scala 23:12]
  assign n121_I_0_0_t1b = n110_O_0_0_t1b; // @[Top.scala 23:12]
  assign n121_I_0_1_t0b = n110_O_0_1_t0b; // @[Top.scala 23:12]
  assign n121_I_0_1_t1b = n110_O_0_1_t1b; // @[Top.scala 23:12]
  assign n121_I_0_2_t0b = n110_O_0_2_t0b; // @[Top.scala 23:12]
  assign n121_I_0_2_t1b = n110_O_0_2_t1b; // @[Top.scala 23:12]
  assign n121_I_1_0_t0b = n110_O_1_0_t0b; // @[Top.scala 23:12]
  assign n121_I_1_0_t1b = n110_O_1_0_t1b; // @[Top.scala 23:12]
  assign n121_I_1_1_t0b = n110_O_1_1_t0b; // @[Top.scala 23:12]
  assign n121_I_1_1_t1b = n110_O_1_1_t1b; // @[Top.scala 23:12]
  assign n121_I_1_2_t0b = n110_O_1_2_t0b; // @[Top.scala 23:12]
  assign n121_I_1_2_t1b = n110_O_1_2_t1b; // @[Top.scala 23:12]
  assign n121_I_2_0_t0b = n110_O_2_0_t0b; // @[Top.scala 23:12]
  assign n121_I_2_0_t1b = n110_O_2_0_t1b; // @[Top.scala 23:12]
  assign n121_I_2_1_t0b = n110_O_2_1_t0b; // @[Top.scala 23:12]
  assign n121_I_2_1_t1b = n110_O_2_1_t1b; // @[Top.scala 23:12]
  assign n121_I_2_2_t0b = n110_O_2_2_t0b; // @[Top.scala 23:12]
  assign n121_I_2_2_t1b = n110_O_2_2_t1b; // @[Top.scala 23:12]
  assign n126_clock = clock;
  assign n126_reset = reset;
  assign n126_valid_up = n121_valid_down; // @[Top.scala 27:19]
  assign n126_I_0_0 = n121_O_0_0; // @[Top.scala 26:12]
  assign n126_I_0_1 = n121_O_0_1; // @[Top.scala 26:12]
  assign n126_I_0_2 = n121_O_0_2; // @[Top.scala 26:12]
  assign n126_I_1_0 = n121_O_1_0; // @[Top.scala 26:12]
  assign n126_I_1_1 = n121_O_1_1; // @[Top.scala 26:12]
  assign n126_I_1_2 = n121_O_1_2; // @[Top.scala 26:12]
  assign n126_I_2_0 = n121_O_2_0; // @[Top.scala 26:12]
  assign n126_I_2_1 = n121_O_2_1; // @[Top.scala 26:12]
  assign n126_I_2_2 = n121_O_2_2; // @[Top.scala 26:12]
  assign n131_clock = clock;
  assign n131_reset = reset;
  assign n131_valid_up = n126_valid_down; // @[Top.scala 30:19]
  assign n131_I_0_0 = n126_O_0_0; // @[Top.scala 29:12]
  assign n131_I_1_0 = n126_O_1_0; // @[Top.scala 29:12]
  assign n131_I_2_0 = n126_O_2_0; // @[Top.scala 29:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n134_valid_up = n131_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 35:19]
  assign n134_I0_0_0 = n131_O_0_0; // @[Top.scala 33:13]
  assign n145_clock = clock;
  assign n145_reset = reset;
  assign n145_valid_up = n134_valid_down; // @[Top.scala 38:19]
  assign n145_I_0_0_t0b = n134_O_0_0_t0b; // @[Top.scala 37:12]
endmodule
module MapS_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0,
  output [15:0] O_4_0_0,
  output [15:0] O_5_0_0,
  output [15:0] O_6_0_0,
  output [15:0] O_7_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_8(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0,
  output [15:0] O_4_0_0,
  output [15:0] O_5_0_0,
  output [15:0] O_6_0_0,
  output [15:0] O_7_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[MapT.scala 8:20]
  MapS_9 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_1_0_0,
  input  [15:0] I_2_0_0,
  input  [15:0] I_3_0_0,
  input  [15:0] I_4_0_0,
  input  [15:0] I_5_0_0,
  input  [15:0] I_6_0_0,
  input  [15:0] I_7_0_0,
  output [15:0] O_0_0,
  output [15:0] O_1_0,
  output [15:0] O_2_0,
  output [15:0] O_3_0,
  output [15:0] O_4_0,
  output [15:0] O_5_0,
  output [15:0] O_6_0,
  output [15:0] O_7_0
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0 = I_1_0_0; // @[Passthrough.scala 17:68]
  assign O_2_0 = I_2_0_0; // @[Passthrough.scala 17:68]
  assign O_3_0 = I_3_0_0; // @[Passthrough.scala 17:68]
  assign O_4_0 = I_4_0_0; // @[Passthrough.scala 17:68]
  assign O_5_0 = I_5_0_0; // @[Passthrough.scala 17:68]
  assign O_6_0 = I_6_0_0; // @[Passthrough.scala 17:68]
  assign O_7_0 = I_7_0_0; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_1_0,
  input  [15:0] I_2_0,
  input  [15:0] I_3_0,
  input  [15:0] I_4_0,
  input  [15:0] I_5_0,
  input  [15:0] I_6_0,
  input  [15:0] I_7_0,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_1_0; // @[Passthrough.scala 17:68]
  assign O_2 = I_2_0; // @[Passthrough.scala 17:68]
  assign O_3 = I_3_0; // @[Passthrough.scala 17:68]
  assign O_4 = I_4_0; // @[Passthrough.scala 17:68]
  assign O_5 = I_5_0; // @[Passthrough.scala 17:68]
  assign O_6 = I_6_0; // @[Passthrough.scala 17:68]
  assign O_7 = I_7_0; // @[Passthrough.scala 17:68]
endmodule
module Top(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7
);
  wire  n1_clock; // @[Top.scala 46:20]
  wire  n1_reset; // @[Top.scala 46:20]
  wire  n1_valid_up; // @[Top.scala 46:20]
  wire  n1_valid_down; // @[Top.scala 46:20]
  wire [15:0] n1_I_0; // @[Top.scala 46:20]
  wire [15:0] n1_I_1; // @[Top.scala 46:20]
  wire [15:0] n1_I_2; // @[Top.scala 46:20]
  wire [15:0] n1_I_3; // @[Top.scala 46:20]
  wire [15:0] n1_I_4; // @[Top.scala 46:20]
  wire [15:0] n1_I_5; // @[Top.scala 46:20]
  wire [15:0] n1_I_6; // @[Top.scala 46:20]
  wire [15:0] n1_I_7; // @[Top.scala 46:20]
  wire [15:0] n1_O_0; // @[Top.scala 46:20]
  wire [15:0] n1_O_1; // @[Top.scala 46:20]
  wire [15:0] n1_O_2; // @[Top.scala 46:20]
  wire [15:0] n1_O_3; // @[Top.scala 46:20]
  wire [15:0] n1_O_4; // @[Top.scala 46:20]
  wire [15:0] n1_O_5; // @[Top.scala 46:20]
  wire [15:0] n1_O_6; // @[Top.scala 46:20]
  wire [15:0] n1_O_7; // @[Top.scala 46:20]
  wire  n2_clock; // @[Top.scala 49:20]
  wire  n2_reset; // @[Top.scala 49:20]
  wire  n2_valid_up; // @[Top.scala 49:20]
  wire  n2_valid_down; // @[Top.scala 49:20]
  wire [15:0] n2_I_0; // @[Top.scala 49:20]
  wire [15:0] n2_I_1; // @[Top.scala 49:20]
  wire [15:0] n2_I_2; // @[Top.scala 49:20]
  wire [15:0] n2_I_3; // @[Top.scala 49:20]
  wire [15:0] n2_I_4; // @[Top.scala 49:20]
  wire [15:0] n2_I_5; // @[Top.scala 49:20]
  wire [15:0] n2_I_6; // @[Top.scala 49:20]
  wire [15:0] n2_I_7; // @[Top.scala 49:20]
  wire [15:0] n2_O_0; // @[Top.scala 49:20]
  wire [15:0] n2_O_1; // @[Top.scala 49:20]
  wire [15:0] n2_O_2; // @[Top.scala 49:20]
  wire [15:0] n2_O_3; // @[Top.scala 49:20]
  wire [15:0] n2_O_4; // @[Top.scala 49:20]
  wire [15:0] n2_O_5; // @[Top.scala 49:20]
  wire [15:0] n2_O_6; // @[Top.scala 49:20]
  wire [15:0] n2_O_7; // @[Top.scala 49:20]
  wire  n3_clock; // @[Top.scala 52:20]
  wire  n3_reset; // @[Top.scala 52:20]
  wire  n3_valid_up; // @[Top.scala 52:20]
  wire  n3_valid_down; // @[Top.scala 52:20]
  wire [15:0] n3_I_0; // @[Top.scala 52:20]
  wire [15:0] n3_I_1; // @[Top.scala 52:20]
  wire [15:0] n3_I_2; // @[Top.scala 52:20]
  wire [15:0] n3_I_3; // @[Top.scala 52:20]
  wire [15:0] n3_I_4; // @[Top.scala 52:20]
  wire [15:0] n3_I_5; // @[Top.scala 52:20]
  wire [15:0] n3_I_6; // @[Top.scala 52:20]
  wire [15:0] n3_I_7; // @[Top.scala 52:20]
  wire [15:0] n3_O_0; // @[Top.scala 52:20]
  wire [15:0] n3_O_1; // @[Top.scala 52:20]
  wire [15:0] n3_O_2; // @[Top.scala 52:20]
  wire [15:0] n3_O_3; // @[Top.scala 52:20]
  wire [15:0] n3_O_4; // @[Top.scala 52:20]
  wire [15:0] n3_O_5; // @[Top.scala 52:20]
  wire [15:0] n3_O_6; // @[Top.scala 52:20]
  wire [15:0] n3_O_7; // @[Top.scala 52:20]
  wire  n4_clock; // @[Top.scala 55:20]
  wire  n4_valid_up; // @[Top.scala 55:20]
  wire  n4_valid_down; // @[Top.scala 55:20]
  wire [15:0] n4_I_0; // @[Top.scala 55:20]
  wire [15:0] n4_I_1; // @[Top.scala 55:20]
  wire [15:0] n4_I_2; // @[Top.scala 55:20]
  wire [15:0] n4_I_3; // @[Top.scala 55:20]
  wire [15:0] n4_I_4; // @[Top.scala 55:20]
  wire [15:0] n4_I_5; // @[Top.scala 55:20]
  wire [15:0] n4_I_6; // @[Top.scala 55:20]
  wire [15:0] n4_I_7; // @[Top.scala 55:20]
  wire [15:0] n4_O_0; // @[Top.scala 55:20]
  wire [15:0] n4_O_1; // @[Top.scala 55:20]
  wire [15:0] n4_O_2; // @[Top.scala 55:20]
  wire [15:0] n4_O_3; // @[Top.scala 55:20]
  wire [15:0] n4_O_4; // @[Top.scala 55:20]
  wire [15:0] n4_O_5; // @[Top.scala 55:20]
  wire [15:0] n4_O_6; // @[Top.scala 55:20]
  wire [15:0] n4_O_7; // @[Top.scala 55:20]
  wire  n5_clock; // @[Top.scala 58:20]
  wire  n5_valid_up; // @[Top.scala 58:20]
  wire  n5_valid_down; // @[Top.scala 58:20]
  wire [15:0] n5_I_0; // @[Top.scala 58:20]
  wire [15:0] n5_I_1; // @[Top.scala 58:20]
  wire [15:0] n5_I_2; // @[Top.scala 58:20]
  wire [15:0] n5_I_3; // @[Top.scala 58:20]
  wire [15:0] n5_I_4; // @[Top.scala 58:20]
  wire [15:0] n5_I_5; // @[Top.scala 58:20]
  wire [15:0] n5_I_6; // @[Top.scala 58:20]
  wire [15:0] n5_I_7; // @[Top.scala 58:20]
  wire [15:0] n5_O_0; // @[Top.scala 58:20]
  wire [15:0] n5_O_1; // @[Top.scala 58:20]
  wire [15:0] n5_O_2; // @[Top.scala 58:20]
  wire [15:0] n5_O_3; // @[Top.scala 58:20]
  wire [15:0] n5_O_4; // @[Top.scala 58:20]
  wire [15:0] n5_O_5; // @[Top.scala 58:20]
  wire [15:0] n5_O_6; // @[Top.scala 58:20]
  wire [15:0] n5_O_7; // @[Top.scala 58:20]
  wire  n6_valid_up; // @[Top.scala 61:20]
  wire  n6_valid_down; // @[Top.scala 61:20]
  wire [15:0] n6_I0_0; // @[Top.scala 61:20]
  wire [15:0] n6_I0_1; // @[Top.scala 61:20]
  wire [15:0] n6_I0_2; // @[Top.scala 61:20]
  wire [15:0] n6_I0_3; // @[Top.scala 61:20]
  wire [15:0] n6_I0_4; // @[Top.scala 61:20]
  wire [15:0] n6_I0_5; // @[Top.scala 61:20]
  wire [15:0] n6_I0_6; // @[Top.scala 61:20]
  wire [15:0] n6_I0_7; // @[Top.scala 61:20]
  wire [15:0] n6_I1_0; // @[Top.scala 61:20]
  wire [15:0] n6_I1_1; // @[Top.scala 61:20]
  wire [15:0] n6_I1_2; // @[Top.scala 61:20]
  wire [15:0] n6_I1_3; // @[Top.scala 61:20]
  wire [15:0] n6_I1_4; // @[Top.scala 61:20]
  wire [15:0] n6_I1_5; // @[Top.scala 61:20]
  wire [15:0] n6_I1_6; // @[Top.scala 61:20]
  wire [15:0] n6_I1_7; // @[Top.scala 61:20]
  wire [15:0] n6_O_0_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_0_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_1_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_1_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_2_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_2_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_3_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_3_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_4_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_4_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_5_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_5_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_6_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_6_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_7_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_7_1; // @[Top.scala 61:20]
  wire  n13_valid_up; // @[Top.scala 65:21]
  wire  n13_valid_down; // @[Top.scala 65:21]
  wire [15:0] n13_I0_0_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_0_1; // @[Top.scala 65:21]
  wire [15:0] n13_I0_1_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_1_1; // @[Top.scala 65:21]
  wire [15:0] n13_I0_2_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_2_1; // @[Top.scala 65:21]
  wire [15:0] n13_I0_3_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_3_1; // @[Top.scala 65:21]
  wire [15:0] n13_I0_4_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_4_1; // @[Top.scala 65:21]
  wire [15:0] n13_I0_5_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_5_1; // @[Top.scala 65:21]
  wire [15:0] n13_I0_6_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_6_1; // @[Top.scala 65:21]
  wire [15:0] n13_I0_7_0; // @[Top.scala 65:21]
  wire [15:0] n13_I0_7_1; // @[Top.scala 65:21]
  wire [15:0] n13_I1_0; // @[Top.scala 65:21]
  wire [15:0] n13_I1_1; // @[Top.scala 65:21]
  wire [15:0] n13_I1_2; // @[Top.scala 65:21]
  wire [15:0] n13_I1_3; // @[Top.scala 65:21]
  wire [15:0] n13_I1_4; // @[Top.scala 65:21]
  wire [15:0] n13_I1_5; // @[Top.scala 65:21]
  wire [15:0] n13_I1_6; // @[Top.scala 65:21]
  wire [15:0] n13_I1_7; // @[Top.scala 65:21]
  wire [15:0] n13_O_0_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_0_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_0_2; // @[Top.scala 65:21]
  wire [15:0] n13_O_1_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_1_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_1_2; // @[Top.scala 65:21]
  wire [15:0] n13_O_2_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_2_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_2_2; // @[Top.scala 65:21]
  wire [15:0] n13_O_3_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_3_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_3_2; // @[Top.scala 65:21]
  wire [15:0] n13_O_4_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_4_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_4_2; // @[Top.scala 65:21]
  wire [15:0] n13_O_5_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_5_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_5_2; // @[Top.scala 65:21]
  wire [15:0] n13_O_6_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_6_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_6_2; // @[Top.scala 65:21]
  wire [15:0] n13_O_7_0; // @[Top.scala 65:21]
  wire [15:0] n13_O_7_1; // @[Top.scala 65:21]
  wire [15:0] n13_O_7_2; // @[Top.scala 65:21]
  wire  n22_valid_up; // @[Top.scala 69:21]
  wire  n22_valid_down; // @[Top.scala 69:21]
  wire [15:0] n22_I_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_I_1_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_1_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_1_2; // @[Top.scala 69:21]
  wire [15:0] n22_I_2_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_2_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_2_2; // @[Top.scala 69:21]
  wire [15:0] n22_I_3_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_3_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_3_2; // @[Top.scala 69:21]
  wire [15:0] n22_I_4_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_4_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_4_2; // @[Top.scala 69:21]
  wire [15:0] n22_I_5_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_5_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_5_2; // @[Top.scala 69:21]
  wire [15:0] n22_I_6_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_6_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_6_2; // @[Top.scala 69:21]
  wire [15:0] n22_I_7_0; // @[Top.scala 69:21]
  wire [15:0] n22_I_7_1; // @[Top.scala 69:21]
  wire [15:0] n22_I_7_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_0_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_0_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_0_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_1_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_1_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_1_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_2_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_2_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_2_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_3_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_3_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_3_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_4_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_4_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_4_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_5_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_5_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_5_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_6_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_6_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_6_0_2; // @[Top.scala 69:21]
  wire [15:0] n22_O_7_0_0; // @[Top.scala 69:21]
  wire [15:0] n22_O_7_0_1; // @[Top.scala 69:21]
  wire [15:0] n22_O_7_0_2; // @[Top.scala 69:21]
  wire  n29_valid_up; // @[Top.scala 72:21]
  wire  n29_valid_down; // @[Top.scala 72:21]
  wire [15:0] n29_I_0_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_0_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_0_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_I_1_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_1_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_1_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_I_2_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_2_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_2_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_I_3_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_3_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_3_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_I_4_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_4_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_4_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_I_5_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_5_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_5_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_I_6_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_6_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_6_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_I_7_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_I_7_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_I_7_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_0_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_0_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_0_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_1_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_1_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_1_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_2_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_2_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_2_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_3_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_3_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_3_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_4_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_4_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_4_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_5_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_5_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_5_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_6_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_6_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_6_2; // @[Top.scala 72:21]
  wire [15:0] n29_O_7_0; // @[Top.scala 72:21]
  wire [15:0] n29_O_7_1; // @[Top.scala 72:21]
  wire [15:0] n29_O_7_2; // @[Top.scala 72:21]
  wire  n30_clock; // @[Top.scala 75:21]
  wire  n30_valid_up; // @[Top.scala 75:21]
  wire  n30_valid_down; // @[Top.scala 75:21]
  wire [15:0] n30_I_0; // @[Top.scala 75:21]
  wire [15:0] n30_I_1; // @[Top.scala 75:21]
  wire [15:0] n30_I_2; // @[Top.scala 75:21]
  wire [15:0] n30_I_3; // @[Top.scala 75:21]
  wire [15:0] n30_I_4; // @[Top.scala 75:21]
  wire [15:0] n30_I_5; // @[Top.scala 75:21]
  wire [15:0] n30_I_6; // @[Top.scala 75:21]
  wire [15:0] n30_I_7; // @[Top.scala 75:21]
  wire [15:0] n30_O_0; // @[Top.scala 75:21]
  wire [15:0] n30_O_1; // @[Top.scala 75:21]
  wire [15:0] n30_O_2; // @[Top.scala 75:21]
  wire [15:0] n30_O_3; // @[Top.scala 75:21]
  wire [15:0] n30_O_4; // @[Top.scala 75:21]
  wire [15:0] n30_O_5; // @[Top.scala 75:21]
  wire [15:0] n30_O_6; // @[Top.scala 75:21]
  wire [15:0] n30_O_7; // @[Top.scala 75:21]
  wire  n31_clock; // @[Top.scala 78:21]
  wire  n31_valid_up; // @[Top.scala 78:21]
  wire  n31_valid_down; // @[Top.scala 78:21]
  wire [15:0] n31_I_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_3; // @[Top.scala 78:21]
  wire [15:0] n31_I_4; // @[Top.scala 78:21]
  wire [15:0] n31_I_5; // @[Top.scala 78:21]
  wire [15:0] n31_I_6; // @[Top.scala 78:21]
  wire [15:0] n31_I_7; // @[Top.scala 78:21]
  wire [15:0] n31_O_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_3; // @[Top.scala 78:21]
  wire [15:0] n31_O_4; // @[Top.scala 78:21]
  wire [15:0] n31_O_5; // @[Top.scala 78:21]
  wire [15:0] n31_O_6; // @[Top.scala 78:21]
  wire [15:0] n31_O_7; // @[Top.scala 78:21]
  wire  n32_valid_up; // @[Top.scala 81:21]
  wire  n32_valid_down; // @[Top.scala 81:21]
  wire [15:0] n32_I0_0; // @[Top.scala 81:21]
  wire [15:0] n32_I0_1; // @[Top.scala 81:21]
  wire [15:0] n32_I0_2; // @[Top.scala 81:21]
  wire [15:0] n32_I0_3; // @[Top.scala 81:21]
  wire [15:0] n32_I0_4; // @[Top.scala 81:21]
  wire [15:0] n32_I0_5; // @[Top.scala 81:21]
  wire [15:0] n32_I0_6; // @[Top.scala 81:21]
  wire [15:0] n32_I0_7; // @[Top.scala 81:21]
  wire [15:0] n32_I1_0; // @[Top.scala 81:21]
  wire [15:0] n32_I1_1; // @[Top.scala 81:21]
  wire [15:0] n32_I1_2; // @[Top.scala 81:21]
  wire [15:0] n32_I1_3; // @[Top.scala 81:21]
  wire [15:0] n32_I1_4; // @[Top.scala 81:21]
  wire [15:0] n32_I1_5; // @[Top.scala 81:21]
  wire [15:0] n32_I1_6; // @[Top.scala 81:21]
  wire [15:0] n32_I1_7; // @[Top.scala 81:21]
  wire [15:0] n32_O_0_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_0_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_1_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_1_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_2_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_2_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_3_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_3_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_4_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_4_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_5_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_5_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_6_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_6_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_7_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_7_1; // @[Top.scala 81:21]
  wire  n39_valid_up; // @[Top.scala 85:21]
  wire  n39_valid_down; // @[Top.scala 85:21]
  wire [15:0] n39_I0_0_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_0_1; // @[Top.scala 85:21]
  wire [15:0] n39_I0_1_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_1_1; // @[Top.scala 85:21]
  wire [15:0] n39_I0_2_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_2_1; // @[Top.scala 85:21]
  wire [15:0] n39_I0_3_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_3_1; // @[Top.scala 85:21]
  wire [15:0] n39_I0_4_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_4_1; // @[Top.scala 85:21]
  wire [15:0] n39_I0_5_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_5_1; // @[Top.scala 85:21]
  wire [15:0] n39_I0_6_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_6_1; // @[Top.scala 85:21]
  wire [15:0] n39_I0_7_0; // @[Top.scala 85:21]
  wire [15:0] n39_I0_7_1; // @[Top.scala 85:21]
  wire [15:0] n39_I1_0; // @[Top.scala 85:21]
  wire [15:0] n39_I1_1; // @[Top.scala 85:21]
  wire [15:0] n39_I1_2; // @[Top.scala 85:21]
  wire [15:0] n39_I1_3; // @[Top.scala 85:21]
  wire [15:0] n39_I1_4; // @[Top.scala 85:21]
  wire [15:0] n39_I1_5; // @[Top.scala 85:21]
  wire [15:0] n39_I1_6; // @[Top.scala 85:21]
  wire [15:0] n39_I1_7; // @[Top.scala 85:21]
  wire [15:0] n39_O_0_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_0_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_0_2; // @[Top.scala 85:21]
  wire [15:0] n39_O_1_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_1_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_1_2; // @[Top.scala 85:21]
  wire [15:0] n39_O_2_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_2_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_2_2; // @[Top.scala 85:21]
  wire [15:0] n39_O_3_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_3_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_3_2; // @[Top.scala 85:21]
  wire [15:0] n39_O_4_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_4_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_4_2; // @[Top.scala 85:21]
  wire [15:0] n39_O_5_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_5_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_5_2; // @[Top.scala 85:21]
  wire [15:0] n39_O_6_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_6_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_6_2; // @[Top.scala 85:21]
  wire [15:0] n39_O_7_0; // @[Top.scala 85:21]
  wire [15:0] n39_O_7_1; // @[Top.scala 85:21]
  wire [15:0] n39_O_7_2; // @[Top.scala 85:21]
  wire  n48_valid_up; // @[Top.scala 89:21]
  wire  n48_valid_down; // @[Top.scala 89:21]
  wire [15:0] n48_I_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_I_1_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_1_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_1_2; // @[Top.scala 89:21]
  wire [15:0] n48_I_2_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_2_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_2_2; // @[Top.scala 89:21]
  wire [15:0] n48_I_3_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_3_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_3_2; // @[Top.scala 89:21]
  wire [15:0] n48_I_4_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_4_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_4_2; // @[Top.scala 89:21]
  wire [15:0] n48_I_5_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_5_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_5_2; // @[Top.scala 89:21]
  wire [15:0] n48_I_6_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_6_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_6_2; // @[Top.scala 89:21]
  wire [15:0] n48_I_7_0; // @[Top.scala 89:21]
  wire [15:0] n48_I_7_1; // @[Top.scala 89:21]
  wire [15:0] n48_I_7_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_0_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_0_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_0_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_1_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_1_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_1_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_2_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_2_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_2_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_3_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_3_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_3_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_4_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_4_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_4_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_5_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_5_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_5_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_6_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_6_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_6_0_2; // @[Top.scala 89:21]
  wire [15:0] n48_O_7_0_0; // @[Top.scala 89:21]
  wire [15:0] n48_O_7_0_1; // @[Top.scala 89:21]
  wire [15:0] n48_O_7_0_2; // @[Top.scala 89:21]
  wire  n55_valid_up; // @[Top.scala 92:21]
  wire  n55_valid_down; // @[Top.scala 92:21]
  wire [15:0] n55_I_0_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_0_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_0_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_I_1_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_1_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_1_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_I_2_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_2_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_2_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_I_3_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_3_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_3_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_I_4_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_4_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_4_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_I_5_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_5_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_5_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_I_6_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_6_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_6_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_I_7_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_I_7_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_I_7_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_0_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_0_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_0_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_1_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_1_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_1_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_2_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_2_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_2_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_3_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_3_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_3_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_4_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_4_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_4_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_5_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_5_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_5_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_6_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_6_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_6_2; // @[Top.scala 92:21]
  wire [15:0] n55_O_7_0; // @[Top.scala 92:21]
  wire [15:0] n55_O_7_1; // @[Top.scala 92:21]
  wire [15:0] n55_O_7_2; // @[Top.scala 92:21]
  wire  n56_valid_up; // @[Top.scala 95:21]
  wire  n56_valid_down; // @[Top.scala 95:21]
  wire [15:0] n56_I0_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_I0_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_I0_2_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_2_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_2_2; // @[Top.scala 95:21]
  wire [15:0] n56_I0_3_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_3_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_3_2; // @[Top.scala 95:21]
  wire [15:0] n56_I0_4_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_4_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_4_2; // @[Top.scala 95:21]
  wire [15:0] n56_I0_5_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_5_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_5_2; // @[Top.scala 95:21]
  wire [15:0] n56_I0_6_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_6_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_6_2; // @[Top.scala 95:21]
  wire [15:0] n56_I0_7_0; // @[Top.scala 95:21]
  wire [15:0] n56_I0_7_1; // @[Top.scala 95:21]
  wire [15:0] n56_I0_7_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_2_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_2_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_2_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_3_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_3_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_3_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_4_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_4_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_4_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_5_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_5_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_5_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_6_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_6_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_6_2; // @[Top.scala 95:21]
  wire [15:0] n56_I1_7_0; // @[Top.scala 95:21]
  wire [15:0] n56_I1_7_1; // @[Top.scala 95:21]
  wire [15:0] n56_I1_7_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_0_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_0_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_0_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_0_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_0_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_0_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_1_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_1_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_1_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_1_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_1_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_1_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_2_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_2_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_2_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_2_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_2_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_2_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_3_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_3_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_3_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_3_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_3_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_3_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_4_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_4_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_4_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_4_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_4_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_4_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_5_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_5_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_5_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_5_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_5_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_5_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_6_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_6_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_6_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_6_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_6_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_6_1_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_7_0_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_7_0_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_7_0_2; // @[Top.scala 95:21]
  wire [15:0] n56_O_7_1_0; // @[Top.scala 95:21]
  wire [15:0] n56_O_7_1_1; // @[Top.scala 95:21]
  wire [15:0] n56_O_7_1_2; // @[Top.scala 95:21]
  wire  n63_clock; // @[Top.scala 99:21]
  wire  n63_valid_up; // @[Top.scala 99:21]
  wire  n63_valid_down; // @[Top.scala 99:21]
  wire [15:0] n63_I_0; // @[Top.scala 99:21]
  wire [15:0] n63_I_1; // @[Top.scala 99:21]
  wire [15:0] n63_I_2; // @[Top.scala 99:21]
  wire [15:0] n63_I_3; // @[Top.scala 99:21]
  wire [15:0] n63_I_4; // @[Top.scala 99:21]
  wire [15:0] n63_I_5; // @[Top.scala 99:21]
  wire [15:0] n63_I_6; // @[Top.scala 99:21]
  wire [15:0] n63_I_7; // @[Top.scala 99:21]
  wire [15:0] n63_O_0; // @[Top.scala 99:21]
  wire [15:0] n63_O_1; // @[Top.scala 99:21]
  wire [15:0] n63_O_2; // @[Top.scala 99:21]
  wire [15:0] n63_O_3; // @[Top.scala 99:21]
  wire [15:0] n63_O_4; // @[Top.scala 99:21]
  wire [15:0] n63_O_5; // @[Top.scala 99:21]
  wire [15:0] n63_O_6; // @[Top.scala 99:21]
  wire [15:0] n63_O_7; // @[Top.scala 99:21]
  wire  n64_clock; // @[Top.scala 102:21]
  wire  n64_valid_up; // @[Top.scala 102:21]
  wire  n64_valid_down; // @[Top.scala 102:21]
  wire [15:0] n64_I_0; // @[Top.scala 102:21]
  wire [15:0] n64_I_1; // @[Top.scala 102:21]
  wire [15:0] n64_I_2; // @[Top.scala 102:21]
  wire [15:0] n64_I_3; // @[Top.scala 102:21]
  wire [15:0] n64_I_4; // @[Top.scala 102:21]
  wire [15:0] n64_I_5; // @[Top.scala 102:21]
  wire [15:0] n64_I_6; // @[Top.scala 102:21]
  wire [15:0] n64_I_7; // @[Top.scala 102:21]
  wire [15:0] n64_O_0; // @[Top.scala 102:21]
  wire [15:0] n64_O_1; // @[Top.scala 102:21]
  wire [15:0] n64_O_2; // @[Top.scala 102:21]
  wire [15:0] n64_O_3; // @[Top.scala 102:21]
  wire [15:0] n64_O_4; // @[Top.scala 102:21]
  wire [15:0] n64_O_5; // @[Top.scala 102:21]
  wire [15:0] n64_O_6; // @[Top.scala 102:21]
  wire [15:0] n64_O_7; // @[Top.scala 102:21]
  wire  n65_valid_up; // @[Top.scala 105:21]
  wire  n65_valid_down; // @[Top.scala 105:21]
  wire [15:0] n65_I0_0; // @[Top.scala 105:21]
  wire [15:0] n65_I0_1; // @[Top.scala 105:21]
  wire [15:0] n65_I0_2; // @[Top.scala 105:21]
  wire [15:0] n65_I0_3; // @[Top.scala 105:21]
  wire [15:0] n65_I0_4; // @[Top.scala 105:21]
  wire [15:0] n65_I0_5; // @[Top.scala 105:21]
  wire [15:0] n65_I0_6; // @[Top.scala 105:21]
  wire [15:0] n65_I0_7; // @[Top.scala 105:21]
  wire [15:0] n65_I1_0; // @[Top.scala 105:21]
  wire [15:0] n65_I1_1; // @[Top.scala 105:21]
  wire [15:0] n65_I1_2; // @[Top.scala 105:21]
  wire [15:0] n65_I1_3; // @[Top.scala 105:21]
  wire [15:0] n65_I1_4; // @[Top.scala 105:21]
  wire [15:0] n65_I1_5; // @[Top.scala 105:21]
  wire [15:0] n65_I1_6; // @[Top.scala 105:21]
  wire [15:0] n65_I1_7; // @[Top.scala 105:21]
  wire [15:0] n65_O_0_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_0_1; // @[Top.scala 105:21]
  wire [15:0] n65_O_1_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_1_1; // @[Top.scala 105:21]
  wire [15:0] n65_O_2_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_2_1; // @[Top.scala 105:21]
  wire [15:0] n65_O_3_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_3_1; // @[Top.scala 105:21]
  wire [15:0] n65_O_4_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_4_1; // @[Top.scala 105:21]
  wire [15:0] n65_O_5_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_5_1; // @[Top.scala 105:21]
  wire [15:0] n65_O_6_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_6_1; // @[Top.scala 105:21]
  wire [15:0] n65_O_7_0; // @[Top.scala 105:21]
  wire [15:0] n65_O_7_1; // @[Top.scala 105:21]
  wire  n72_valid_up; // @[Top.scala 109:21]
  wire  n72_valid_down; // @[Top.scala 109:21]
  wire [15:0] n72_I0_0_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_0_1; // @[Top.scala 109:21]
  wire [15:0] n72_I0_1_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_1_1; // @[Top.scala 109:21]
  wire [15:0] n72_I0_2_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_2_1; // @[Top.scala 109:21]
  wire [15:0] n72_I0_3_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_3_1; // @[Top.scala 109:21]
  wire [15:0] n72_I0_4_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_4_1; // @[Top.scala 109:21]
  wire [15:0] n72_I0_5_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_5_1; // @[Top.scala 109:21]
  wire [15:0] n72_I0_6_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_6_1; // @[Top.scala 109:21]
  wire [15:0] n72_I0_7_0; // @[Top.scala 109:21]
  wire [15:0] n72_I0_7_1; // @[Top.scala 109:21]
  wire [15:0] n72_I1_0; // @[Top.scala 109:21]
  wire [15:0] n72_I1_1; // @[Top.scala 109:21]
  wire [15:0] n72_I1_2; // @[Top.scala 109:21]
  wire [15:0] n72_I1_3; // @[Top.scala 109:21]
  wire [15:0] n72_I1_4; // @[Top.scala 109:21]
  wire [15:0] n72_I1_5; // @[Top.scala 109:21]
  wire [15:0] n72_I1_6; // @[Top.scala 109:21]
  wire [15:0] n72_I1_7; // @[Top.scala 109:21]
  wire [15:0] n72_O_0_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_0_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_0_2; // @[Top.scala 109:21]
  wire [15:0] n72_O_1_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_1_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_1_2; // @[Top.scala 109:21]
  wire [15:0] n72_O_2_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_2_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_2_2; // @[Top.scala 109:21]
  wire [15:0] n72_O_3_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_3_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_3_2; // @[Top.scala 109:21]
  wire [15:0] n72_O_4_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_4_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_4_2; // @[Top.scala 109:21]
  wire [15:0] n72_O_5_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_5_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_5_2; // @[Top.scala 109:21]
  wire [15:0] n72_O_6_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_6_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_6_2; // @[Top.scala 109:21]
  wire [15:0] n72_O_7_0; // @[Top.scala 109:21]
  wire [15:0] n72_O_7_1; // @[Top.scala 109:21]
  wire [15:0] n72_O_7_2; // @[Top.scala 109:21]
  wire  n81_valid_up; // @[Top.scala 113:21]
  wire  n81_valid_down; // @[Top.scala 113:21]
  wire [15:0] n81_I_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_I_1_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_1_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_1_2; // @[Top.scala 113:21]
  wire [15:0] n81_I_2_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_2_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_2_2; // @[Top.scala 113:21]
  wire [15:0] n81_I_3_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_3_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_3_2; // @[Top.scala 113:21]
  wire [15:0] n81_I_4_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_4_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_4_2; // @[Top.scala 113:21]
  wire [15:0] n81_I_5_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_5_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_5_2; // @[Top.scala 113:21]
  wire [15:0] n81_I_6_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_6_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_6_2; // @[Top.scala 113:21]
  wire [15:0] n81_I_7_0; // @[Top.scala 113:21]
  wire [15:0] n81_I_7_1; // @[Top.scala 113:21]
  wire [15:0] n81_I_7_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_0_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_0_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_0_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_1_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_1_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_1_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_2_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_2_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_2_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_3_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_3_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_3_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_4_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_4_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_4_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_5_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_5_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_5_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_6_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_6_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_6_0_2; // @[Top.scala 113:21]
  wire [15:0] n81_O_7_0_0; // @[Top.scala 113:21]
  wire [15:0] n81_O_7_0_1; // @[Top.scala 113:21]
  wire [15:0] n81_O_7_0_2; // @[Top.scala 113:21]
  wire  n88_valid_up; // @[Top.scala 116:21]
  wire  n88_valid_down; // @[Top.scala 116:21]
  wire [15:0] n88_I_0_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_0_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_0_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_I_1_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_1_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_1_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_I_2_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_2_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_2_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_I_3_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_3_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_3_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_I_4_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_4_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_4_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_I_5_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_5_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_5_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_I_6_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_6_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_6_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_I_7_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_I_7_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_I_7_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_0_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_0_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_0_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_1_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_1_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_1_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_2_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_2_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_2_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_3_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_3_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_3_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_4_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_4_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_4_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_5_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_5_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_5_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_6_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_6_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_6_2; // @[Top.scala 116:21]
  wire [15:0] n88_O_7_0; // @[Top.scala 116:21]
  wire [15:0] n88_O_7_1; // @[Top.scala 116:21]
  wire [15:0] n88_O_7_2; // @[Top.scala 116:21]
  wire  n89_valid_up; // @[Top.scala 119:21]
  wire  n89_valid_down; // @[Top.scala 119:21]
  wire [15:0] n89_I0_0_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_0_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_0_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_0_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_0_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_0_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_1_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_1_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_1_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_1_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_1_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_1_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_2_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_2_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_2_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_2_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_2_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_2_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_3_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_3_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_3_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_3_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_3_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_3_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_4_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_4_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_4_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_4_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_4_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_4_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_5_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_5_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_5_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_5_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_5_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_5_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_6_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_6_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_6_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_6_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_6_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_6_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_7_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_7_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_7_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I0_7_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I0_7_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I0_7_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_3_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_3_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_3_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_4_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_4_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_4_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_5_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_5_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_5_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_6_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_6_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_6_2; // @[Top.scala 119:21]
  wire [15:0] n89_I1_7_0; // @[Top.scala 119:21]
  wire [15:0] n89_I1_7_1; // @[Top.scala 119:21]
  wire [15:0] n89_I1_7_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_0_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_1_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_2_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_3_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_4_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_5_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_6_2_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_0_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_0_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_0_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_1_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_1_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_1_2; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_2_0; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_2_1; // @[Top.scala 119:21]
  wire [15:0] n89_O_7_2_2; // @[Top.scala 119:21]
  wire  n98_valid_up; // @[Top.scala 123:21]
  wire  n98_valid_down; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_1_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_2_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_3_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_4_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_5_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_6_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_I_7_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_0_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_1_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_2_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_3_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_4_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_5_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_6_0_2_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_0_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_0_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_0_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_1_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_1_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_1_2; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_2_0; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_2_1; // @[Top.scala 123:21]
  wire [15:0] n98_O_7_0_2_2; // @[Top.scala 123:21]
  wire  n105_valid_up; // @[Top.scala 126:22]
  wire  n105_valid_down; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_0_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_1_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_2_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_3_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_4_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_5_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_6_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_I_7_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_0_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_1_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_2_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_3_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_4_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_5_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_6_2_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_0_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_0_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_0_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_1_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_1_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_1_2; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_2_0; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_2_1; // @[Top.scala 126:22]
  wire [15:0] n105_O_7_2_2; // @[Top.scala 126:22]
  wire  n147_clock; // @[Top.scala 129:22]
  wire  n147_reset; // @[Top.scala 129:22]
  wire  n147_valid_up; // @[Top.scala 129:22]
  wire  n147_valid_down; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_0_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_1_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_2_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_3_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_4_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_5_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_6_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_0_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_0_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_1_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_1_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_1_2; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_2_0; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_2_1; // @[Top.scala 129:22]
  wire [15:0] n147_I_7_2_2; // @[Top.scala 129:22]
  wire [15:0] n147_O_0_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_O_1_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_O_2_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_O_3_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_O_4_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_O_5_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_O_6_0_0; // @[Top.scala 129:22]
  wire [15:0] n147_O_7_0_0; // @[Top.scala 129:22]
  wire  n148_valid_up; // @[Top.scala 132:22]
  wire  n148_valid_down; // @[Top.scala 132:22]
  wire [15:0] n148_I_0_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_I_1_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_I_2_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_I_3_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_I_4_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_I_5_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_I_6_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_I_7_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_0_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_1_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_2_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_3_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_4_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_5_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_6_0; // @[Top.scala 132:22]
  wire [15:0] n148_O_7_0; // @[Top.scala 132:22]
  wire  n149_valid_up; // @[Top.scala 135:22]
  wire  n149_valid_down; // @[Top.scala 135:22]
  wire [15:0] n149_I_0_0; // @[Top.scala 135:22]
  wire [15:0] n149_I_1_0; // @[Top.scala 135:22]
  wire [15:0] n149_I_2_0; // @[Top.scala 135:22]
  wire [15:0] n149_I_3_0; // @[Top.scala 135:22]
  wire [15:0] n149_I_4_0; // @[Top.scala 135:22]
  wire [15:0] n149_I_5_0; // @[Top.scala 135:22]
  wire [15:0] n149_I_6_0; // @[Top.scala 135:22]
  wire [15:0] n149_I_7_0; // @[Top.scala 135:22]
  wire [15:0] n149_O_0; // @[Top.scala 135:22]
  wire [15:0] n149_O_1; // @[Top.scala 135:22]
  wire [15:0] n149_O_2; // @[Top.scala 135:22]
  wire [15:0] n149_O_3; // @[Top.scala 135:22]
  wire [15:0] n149_O_4; // @[Top.scala 135:22]
  wire [15:0] n149_O_5; // @[Top.scala 135:22]
  wire [15:0] n149_O_6; // @[Top.scala 135:22]
  wire [15:0] n149_O_7; // @[Top.scala 135:22]
  wire  n150_clock; // @[Top.scala 138:22]
  wire  n150_reset; // @[Top.scala 138:22]
  wire  n150_valid_up; // @[Top.scala 138:22]
  wire  n150_valid_down; // @[Top.scala 138:22]
  wire [15:0] n150_I_0; // @[Top.scala 138:22]
  wire [15:0] n150_I_1; // @[Top.scala 138:22]
  wire [15:0] n150_I_2; // @[Top.scala 138:22]
  wire [15:0] n150_I_3; // @[Top.scala 138:22]
  wire [15:0] n150_I_4; // @[Top.scala 138:22]
  wire [15:0] n150_I_5; // @[Top.scala 138:22]
  wire [15:0] n150_I_6; // @[Top.scala 138:22]
  wire [15:0] n150_I_7; // @[Top.scala 138:22]
  wire [15:0] n150_O_0; // @[Top.scala 138:22]
  wire [15:0] n150_O_1; // @[Top.scala 138:22]
  wire [15:0] n150_O_2; // @[Top.scala 138:22]
  wire [15:0] n150_O_3; // @[Top.scala 138:22]
  wire [15:0] n150_O_4; // @[Top.scala 138:22]
  wire [15:0] n150_O_5; // @[Top.scala 138:22]
  wire [15:0] n150_O_6; // @[Top.scala 138:22]
  wire [15:0] n150_O_7; // @[Top.scala 138:22]
  wire  n151_clock; // @[Top.scala 141:22]
  wire  n151_reset; // @[Top.scala 141:22]
  wire  n151_valid_up; // @[Top.scala 141:22]
  wire  n151_valid_down; // @[Top.scala 141:22]
  wire [15:0] n151_I_0; // @[Top.scala 141:22]
  wire [15:0] n151_I_1; // @[Top.scala 141:22]
  wire [15:0] n151_I_2; // @[Top.scala 141:22]
  wire [15:0] n151_I_3; // @[Top.scala 141:22]
  wire [15:0] n151_I_4; // @[Top.scala 141:22]
  wire [15:0] n151_I_5; // @[Top.scala 141:22]
  wire [15:0] n151_I_6; // @[Top.scala 141:22]
  wire [15:0] n151_I_7; // @[Top.scala 141:22]
  wire [15:0] n151_O_0; // @[Top.scala 141:22]
  wire [15:0] n151_O_1; // @[Top.scala 141:22]
  wire [15:0] n151_O_2; // @[Top.scala 141:22]
  wire [15:0] n151_O_3; // @[Top.scala 141:22]
  wire [15:0] n151_O_4; // @[Top.scala 141:22]
  wire [15:0] n151_O_5; // @[Top.scala 141:22]
  wire [15:0] n151_O_6; // @[Top.scala 141:22]
  wire [15:0] n151_O_7; // @[Top.scala 141:22]
  wire  n152_clock; // @[Top.scala 144:22]
  wire  n152_reset; // @[Top.scala 144:22]
  wire  n152_valid_up; // @[Top.scala 144:22]
  wire  n152_valid_down; // @[Top.scala 144:22]
  wire [15:0] n152_I_0; // @[Top.scala 144:22]
  wire [15:0] n152_I_1; // @[Top.scala 144:22]
  wire [15:0] n152_I_2; // @[Top.scala 144:22]
  wire [15:0] n152_I_3; // @[Top.scala 144:22]
  wire [15:0] n152_I_4; // @[Top.scala 144:22]
  wire [15:0] n152_I_5; // @[Top.scala 144:22]
  wire [15:0] n152_I_6; // @[Top.scala 144:22]
  wire [15:0] n152_I_7; // @[Top.scala 144:22]
  wire [15:0] n152_O_0; // @[Top.scala 144:22]
  wire [15:0] n152_O_1; // @[Top.scala 144:22]
  wire [15:0] n152_O_2; // @[Top.scala 144:22]
  wire [15:0] n152_O_3; // @[Top.scala 144:22]
  wire [15:0] n152_O_4; // @[Top.scala 144:22]
  wire [15:0] n152_O_5; // @[Top.scala 144:22]
  wire [15:0] n152_O_6; // @[Top.scala 144:22]
  wire [15:0] n152_O_7; // @[Top.scala 144:22]
  FIFO n1 ( // @[Top.scala 46:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7)
  );
  ShiftTS n2 ( // @[Top.scala 49:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .I_2(n2_I_2),
    .I_3(n2_I_3),
    .I_4(n2_I_4),
    .I_5(n2_I_5),
    .I_6(n2_I_6),
    .I_7(n2_I_7),
    .O_0(n2_O_0),
    .O_1(n2_O_1),
    .O_2(n2_O_2),
    .O_3(n2_O_3),
    .O_4(n2_O_4),
    .O_5(n2_O_5),
    .O_6(n2_O_6),
    .O_7(n2_O_7)
  );
  ShiftTS n3 ( // @[Top.scala 52:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .I_2(n3_I_2),
    .I_3(n3_I_3),
    .I_4(n3_I_4),
    .I_5(n3_I_5),
    .I_6(n3_I_6),
    .I_7(n3_I_7),
    .O_0(n3_O_0),
    .O_1(n3_O_1),
    .O_2(n3_O_2),
    .O_3(n3_O_3),
    .O_4(n3_O_4),
    .O_5(n3_O_5),
    .O_6(n3_O_6),
    .O_7(n3_O_7)
  );
  ShiftTS_2 n4 ( // @[Top.scala 55:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .I_2(n4_I_2),
    .I_3(n4_I_3),
    .I_4(n4_I_4),
    .I_5(n4_I_5),
    .I_6(n4_I_6),
    .I_7(n4_I_7),
    .O_0(n4_O_0),
    .O_1(n4_O_1),
    .O_2(n4_O_2),
    .O_3(n4_O_3),
    .O_4(n4_O_4),
    .O_5(n4_O_5),
    .O_6(n4_O_6),
    .O_7(n4_O_7)
  );
  ShiftTS_2 n5 ( // @[Top.scala 58:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .I_2(n5_I_2),
    .I_3(n5_I_3),
    .I_4(n5_I_4),
    .I_5(n5_I_5),
    .I_6(n5_I_6),
    .I_7(n5_I_7),
    .O_0(n5_O_0),
    .O_1(n5_O_1),
    .O_2(n5_O_2),
    .O_3(n5_O_3),
    .O_4(n5_O_4),
    .O_5(n5_O_5),
    .O_6(n5_O_6),
    .O_7(n5_O_7)
  );
  Map2T n6 ( // @[Top.scala 61:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0(n6_I0_0),
    .I0_1(n6_I0_1),
    .I0_2(n6_I0_2),
    .I0_3(n6_I0_3),
    .I0_4(n6_I0_4),
    .I0_5(n6_I0_5),
    .I0_6(n6_I0_6),
    .I0_7(n6_I0_7),
    .I1_0(n6_I1_0),
    .I1_1(n6_I1_1),
    .I1_2(n6_I1_2),
    .I1_3(n6_I1_3),
    .I1_4(n6_I1_4),
    .I1_5(n6_I1_5),
    .I1_6(n6_I1_6),
    .I1_7(n6_I1_7),
    .O_0_0(n6_O_0_0),
    .O_0_1(n6_O_0_1),
    .O_1_0(n6_O_1_0),
    .O_1_1(n6_O_1_1),
    .O_2_0(n6_O_2_0),
    .O_2_1(n6_O_2_1),
    .O_3_0(n6_O_3_0),
    .O_3_1(n6_O_3_1),
    .O_4_0(n6_O_4_0),
    .O_4_1(n6_O_4_1),
    .O_5_0(n6_O_5_0),
    .O_5_1(n6_O_5_1),
    .O_6_0(n6_O_6_0),
    .O_6_1(n6_O_6_1),
    .O_7_0(n6_O_7_0),
    .O_7_1(n6_O_7_1)
  );
  Map2T_1 n13 ( // @[Top.scala 65:21]
    .valid_up(n13_valid_up),
    .valid_down(n13_valid_down),
    .I0_0_0(n13_I0_0_0),
    .I0_0_1(n13_I0_0_1),
    .I0_1_0(n13_I0_1_0),
    .I0_1_1(n13_I0_1_1),
    .I0_2_0(n13_I0_2_0),
    .I0_2_1(n13_I0_2_1),
    .I0_3_0(n13_I0_3_0),
    .I0_3_1(n13_I0_3_1),
    .I0_4_0(n13_I0_4_0),
    .I0_4_1(n13_I0_4_1),
    .I0_5_0(n13_I0_5_0),
    .I0_5_1(n13_I0_5_1),
    .I0_6_0(n13_I0_6_0),
    .I0_6_1(n13_I0_6_1),
    .I0_7_0(n13_I0_7_0),
    .I0_7_1(n13_I0_7_1),
    .I1_0(n13_I1_0),
    .I1_1(n13_I1_1),
    .I1_2(n13_I1_2),
    .I1_3(n13_I1_3),
    .I1_4(n13_I1_4),
    .I1_5(n13_I1_5),
    .I1_6(n13_I1_6),
    .I1_7(n13_I1_7),
    .O_0_0(n13_O_0_0),
    .O_0_1(n13_O_0_1),
    .O_0_2(n13_O_0_2),
    .O_1_0(n13_O_1_0),
    .O_1_1(n13_O_1_1),
    .O_1_2(n13_O_1_2),
    .O_2_0(n13_O_2_0),
    .O_2_1(n13_O_2_1),
    .O_2_2(n13_O_2_2),
    .O_3_0(n13_O_3_0),
    .O_3_1(n13_O_3_1),
    .O_3_2(n13_O_3_2),
    .O_4_0(n13_O_4_0),
    .O_4_1(n13_O_4_1),
    .O_4_2(n13_O_4_2),
    .O_5_0(n13_O_5_0),
    .O_5_1(n13_O_5_1),
    .O_5_2(n13_O_5_2),
    .O_6_0(n13_O_6_0),
    .O_6_1(n13_O_6_1),
    .O_6_2(n13_O_6_2),
    .O_7_0(n13_O_7_0),
    .O_7_1(n13_O_7_1),
    .O_7_2(n13_O_7_2)
  );
  MapT n22 ( // @[Top.scala 69:21]
    .valid_up(n22_valid_up),
    .valid_down(n22_valid_down),
    .I_0_0(n22_I_0_0),
    .I_0_1(n22_I_0_1),
    .I_0_2(n22_I_0_2),
    .I_1_0(n22_I_1_0),
    .I_1_1(n22_I_1_1),
    .I_1_2(n22_I_1_2),
    .I_2_0(n22_I_2_0),
    .I_2_1(n22_I_2_1),
    .I_2_2(n22_I_2_2),
    .I_3_0(n22_I_3_0),
    .I_3_1(n22_I_3_1),
    .I_3_2(n22_I_3_2),
    .I_4_0(n22_I_4_0),
    .I_4_1(n22_I_4_1),
    .I_4_2(n22_I_4_2),
    .I_5_0(n22_I_5_0),
    .I_5_1(n22_I_5_1),
    .I_5_2(n22_I_5_2),
    .I_6_0(n22_I_6_0),
    .I_6_1(n22_I_6_1),
    .I_6_2(n22_I_6_2),
    .I_7_0(n22_I_7_0),
    .I_7_1(n22_I_7_1),
    .I_7_2(n22_I_7_2),
    .O_0_0_0(n22_O_0_0_0),
    .O_0_0_1(n22_O_0_0_1),
    .O_0_0_2(n22_O_0_0_2),
    .O_1_0_0(n22_O_1_0_0),
    .O_1_0_1(n22_O_1_0_1),
    .O_1_0_2(n22_O_1_0_2),
    .O_2_0_0(n22_O_2_0_0),
    .O_2_0_1(n22_O_2_0_1),
    .O_2_0_2(n22_O_2_0_2),
    .O_3_0_0(n22_O_3_0_0),
    .O_3_0_1(n22_O_3_0_1),
    .O_3_0_2(n22_O_3_0_2),
    .O_4_0_0(n22_O_4_0_0),
    .O_4_0_1(n22_O_4_0_1),
    .O_4_0_2(n22_O_4_0_2),
    .O_5_0_0(n22_O_5_0_0),
    .O_5_0_1(n22_O_5_0_1),
    .O_5_0_2(n22_O_5_0_2),
    .O_6_0_0(n22_O_6_0_0),
    .O_6_0_1(n22_O_6_0_1),
    .O_6_0_2(n22_O_6_0_2),
    .O_7_0_0(n22_O_7_0_0),
    .O_7_0_1(n22_O_7_0_1),
    .O_7_0_2(n22_O_7_0_2)
  );
  MapT_1 n29 ( // @[Top.scala 72:21]
    .valid_up(n29_valid_up),
    .valid_down(n29_valid_down),
    .I_0_0_0(n29_I_0_0_0),
    .I_0_0_1(n29_I_0_0_1),
    .I_0_0_2(n29_I_0_0_2),
    .I_1_0_0(n29_I_1_0_0),
    .I_1_0_1(n29_I_1_0_1),
    .I_1_0_2(n29_I_1_0_2),
    .I_2_0_0(n29_I_2_0_0),
    .I_2_0_1(n29_I_2_0_1),
    .I_2_0_2(n29_I_2_0_2),
    .I_3_0_0(n29_I_3_0_0),
    .I_3_0_1(n29_I_3_0_1),
    .I_3_0_2(n29_I_3_0_2),
    .I_4_0_0(n29_I_4_0_0),
    .I_4_0_1(n29_I_4_0_1),
    .I_4_0_2(n29_I_4_0_2),
    .I_5_0_0(n29_I_5_0_0),
    .I_5_0_1(n29_I_5_0_1),
    .I_5_0_2(n29_I_5_0_2),
    .I_6_0_0(n29_I_6_0_0),
    .I_6_0_1(n29_I_6_0_1),
    .I_6_0_2(n29_I_6_0_2),
    .I_7_0_0(n29_I_7_0_0),
    .I_7_0_1(n29_I_7_0_1),
    .I_7_0_2(n29_I_7_0_2),
    .O_0_0(n29_O_0_0),
    .O_0_1(n29_O_0_1),
    .O_0_2(n29_O_0_2),
    .O_1_0(n29_O_1_0),
    .O_1_1(n29_O_1_1),
    .O_1_2(n29_O_1_2),
    .O_2_0(n29_O_2_0),
    .O_2_1(n29_O_2_1),
    .O_2_2(n29_O_2_2),
    .O_3_0(n29_O_3_0),
    .O_3_1(n29_O_3_1),
    .O_3_2(n29_O_3_2),
    .O_4_0(n29_O_4_0),
    .O_4_1(n29_O_4_1),
    .O_4_2(n29_O_4_2),
    .O_5_0(n29_O_5_0),
    .O_5_1(n29_O_5_1),
    .O_5_2(n29_O_5_2),
    .O_6_0(n29_O_6_0),
    .O_6_1(n29_O_6_1),
    .O_6_2(n29_O_6_2),
    .O_7_0(n29_O_7_0),
    .O_7_1(n29_O_7_1),
    .O_7_2(n29_O_7_2)
  );
  ShiftTS_2 n30 ( // @[Top.scala 75:21]
    .clock(n30_clock),
    .valid_up(n30_valid_up),
    .valid_down(n30_valid_down),
    .I_0(n30_I_0),
    .I_1(n30_I_1),
    .I_2(n30_I_2),
    .I_3(n30_I_3),
    .I_4(n30_I_4),
    .I_5(n30_I_5),
    .I_6(n30_I_6),
    .I_7(n30_I_7),
    .O_0(n30_O_0),
    .O_1(n30_O_1),
    .O_2(n30_O_2),
    .O_3(n30_O_3),
    .O_4(n30_O_4),
    .O_5(n30_O_5),
    .O_6(n30_O_6),
    .O_7(n30_O_7)
  );
  ShiftTS_2 n31 ( // @[Top.scala 78:21]
    .clock(n31_clock),
    .valid_up(n31_valid_up),
    .valid_down(n31_valid_down),
    .I_0(n31_I_0),
    .I_1(n31_I_1),
    .I_2(n31_I_2),
    .I_3(n31_I_3),
    .I_4(n31_I_4),
    .I_5(n31_I_5),
    .I_6(n31_I_6),
    .I_7(n31_I_7),
    .O_0(n31_O_0),
    .O_1(n31_O_1),
    .O_2(n31_O_2),
    .O_3(n31_O_3),
    .O_4(n31_O_4),
    .O_5(n31_O_5),
    .O_6(n31_O_6),
    .O_7(n31_O_7)
  );
  Map2T n32 ( // @[Top.scala 81:21]
    .valid_up(n32_valid_up),
    .valid_down(n32_valid_down),
    .I0_0(n32_I0_0),
    .I0_1(n32_I0_1),
    .I0_2(n32_I0_2),
    .I0_3(n32_I0_3),
    .I0_4(n32_I0_4),
    .I0_5(n32_I0_5),
    .I0_6(n32_I0_6),
    .I0_7(n32_I0_7),
    .I1_0(n32_I1_0),
    .I1_1(n32_I1_1),
    .I1_2(n32_I1_2),
    .I1_3(n32_I1_3),
    .I1_4(n32_I1_4),
    .I1_5(n32_I1_5),
    .I1_6(n32_I1_6),
    .I1_7(n32_I1_7),
    .O_0_0(n32_O_0_0),
    .O_0_1(n32_O_0_1),
    .O_1_0(n32_O_1_0),
    .O_1_1(n32_O_1_1),
    .O_2_0(n32_O_2_0),
    .O_2_1(n32_O_2_1),
    .O_3_0(n32_O_3_0),
    .O_3_1(n32_O_3_1),
    .O_4_0(n32_O_4_0),
    .O_4_1(n32_O_4_1),
    .O_5_0(n32_O_5_0),
    .O_5_1(n32_O_5_1),
    .O_6_0(n32_O_6_0),
    .O_6_1(n32_O_6_1),
    .O_7_0(n32_O_7_0),
    .O_7_1(n32_O_7_1)
  );
  Map2T_1 n39 ( // @[Top.scala 85:21]
    .valid_up(n39_valid_up),
    .valid_down(n39_valid_down),
    .I0_0_0(n39_I0_0_0),
    .I0_0_1(n39_I0_0_1),
    .I0_1_0(n39_I0_1_0),
    .I0_1_1(n39_I0_1_1),
    .I0_2_0(n39_I0_2_0),
    .I0_2_1(n39_I0_2_1),
    .I0_3_0(n39_I0_3_0),
    .I0_3_1(n39_I0_3_1),
    .I0_4_0(n39_I0_4_0),
    .I0_4_1(n39_I0_4_1),
    .I0_5_0(n39_I0_5_0),
    .I0_5_1(n39_I0_5_1),
    .I0_6_0(n39_I0_6_0),
    .I0_6_1(n39_I0_6_1),
    .I0_7_0(n39_I0_7_0),
    .I0_7_1(n39_I0_7_1),
    .I1_0(n39_I1_0),
    .I1_1(n39_I1_1),
    .I1_2(n39_I1_2),
    .I1_3(n39_I1_3),
    .I1_4(n39_I1_4),
    .I1_5(n39_I1_5),
    .I1_6(n39_I1_6),
    .I1_7(n39_I1_7),
    .O_0_0(n39_O_0_0),
    .O_0_1(n39_O_0_1),
    .O_0_2(n39_O_0_2),
    .O_1_0(n39_O_1_0),
    .O_1_1(n39_O_1_1),
    .O_1_2(n39_O_1_2),
    .O_2_0(n39_O_2_0),
    .O_2_1(n39_O_2_1),
    .O_2_2(n39_O_2_2),
    .O_3_0(n39_O_3_0),
    .O_3_1(n39_O_3_1),
    .O_3_2(n39_O_3_2),
    .O_4_0(n39_O_4_0),
    .O_4_1(n39_O_4_1),
    .O_4_2(n39_O_4_2),
    .O_5_0(n39_O_5_0),
    .O_5_1(n39_O_5_1),
    .O_5_2(n39_O_5_2),
    .O_6_0(n39_O_6_0),
    .O_6_1(n39_O_6_1),
    .O_6_2(n39_O_6_2),
    .O_7_0(n39_O_7_0),
    .O_7_1(n39_O_7_1),
    .O_7_2(n39_O_7_2)
  );
  MapT n48 ( // @[Top.scala 89:21]
    .valid_up(n48_valid_up),
    .valid_down(n48_valid_down),
    .I_0_0(n48_I_0_0),
    .I_0_1(n48_I_0_1),
    .I_0_2(n48_I_0_2),
    .I_1_0(n48_I_1_0),
    .I_1_1(n48_I_1_1),
    .I_1_2(n48_I_1_2),
    .I_2_0(n48_I_2_0),
    .I_2_1(n48_I_2_1),
    .I_2_2(n48_I_2_2),
    .I_3_0(n48_I_3_0),
    .I_3_1(n48_I_3_1),
    .I_3_2(n48_I_3_2),
    .I_4_0(n48_I_4_0),
    .I_4_1(n48_I_4_1),
    .I_4_2(n48_I_4_2),
    .I_5_0(n48_I_5_0),
    .I_5_1(n48_I_5_1),
    .I_5_2(n48_I_5_2),
    .I_6_0(n48_I_6_0),
    .I_6_1(n48_I_6_1),
    .I_6_2(n48_I_6_2),
    .I_7_0(n48_I_7_0),
    .I_7_1(n48_I_7_1),
    .I_7_2(n48_I_7_2),
    .O_0_0_0(n48_O_0_0_0),
    .O_0_0_1(n48_O_0_0_1),
    .O_0_0_2(n48_O_0_0_2),
    .O_1_0_0(n48_O_1_0_0),
    .O_1_0_1(n48_O_1_0_1),
    .O_1_0_2(n48_O_1_0_2),
    .O_2_0_0(n48_O_2_0_0),
    .O_2_0_1(n48_O_2_0_1),
    .O_2_0_2(n48_O_2_0_2),
    .O_3_0_0(n48_O_3_0_0),
    .O_3_0_1(n48_O_3_0_1),
    .O_3_0_2(n48_O_3_0_2),
    .O_4_0_0(n48_O_4_0_0),
    .O_4_0_1(n48_O_4_0_1),
    .O_4_0_2(n48_O_4_0_2),
    .O_5_0_0(n48_O_5_0_0),
    .O_5_0_1(n48_O_5_0_1),
    .O_5_0_2(n48_O_5_0_2),
    .O_6_0_0(n48_O_6_0_0),
    .O_6_0_1(n48_O_6_0_1),
    .O_6_0_2(n48_O_6_0_2),
    .O_7_0_0(n48_O_7_0_0),
    .O_7_0_1(n48_O_7_0_1),
    .O_7_0_2(n48_O_7_0_2)
  );
  MapT_1 n55 ( // @[Top.scala 92:21]
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I_0_0_0(n55_I_0_0_0),
    .I_0_0_1(n55_I_0_0_1),
    .I_0_0_2(n55_I_0_0_2),
    .I_1_0_0(n55_I_1_0_0),
    .I_1_0_1(n55_I_1_0_1),
    .I_1_0_2(n55_I_1_0_2),
    .I_2_0_0(n55_I_2_0_0),
    .I_2_0_1(n55_I_2_0_1),
    .I_2_0_2(n55_I_2_0_2),
    .I_3_0_0(n55_I_3_0_0),
    .I_3_0_1(n55_I_3_0_1),
    .I_3_0_2(n55_I_3_0_2),
    .I_4_0_0(n55_I_4_0_0),
    .I_4_0_1(n55_I_4_0_1),
    .I_4_0_2(n55_I_4_0_2),
    .I_5_0_0(n55_I_5_0_0),
    .I_5_0_1(n55_I_5_0_1),
    .I_5_0_2(n55_I_5_0_2),
    .I_6_0_0(n55_I_6_0_0),
    .I_6_0_1(n55_I_6_0_1),
    .I_6_0_2(n55_I_6_0_2),
    .I_7_0_0(n55_I_7_0_0),
    .I_7_0_1(n55_I_7_0_1),
    .I_7_0_2(n55_I_7_0_2),
    .O_0_0(n55_O_0_0),
    .O_0_1(n55_O_0_1),
    .O_0_2(n55_O_0_2),
    .O_1_0(n55_O_1_0),
    .O_1_1(n55_O_1_1),
    .O_1_2(n55_O_1_2),
    .O_2_0(n55_O_2_0),
    .O_2_1(n55_O_2_1),
    .O_2_2(n55_O_2_2),
    .O_3_0(n55_O_3_0),
    .O_3_1(n55_O_3_1),
    .O_3_2(n55_O_3_2),
    .O_4_0(n55_O_4_0),
    .O_4_1(n55_O_4_1),
    .O_4_2(n55_O_4_2),
    .O_5_0(n55_O_5_0),
    .O_5_1(n55_O_5_1),
    .O_5_2(n55_O_5_2),
    .O_6_0(n55_O_6_0),
    .O_6_1(n55_O_6_1),
    .O_6_2(n55_O_6_2),
    .O_7_0(n55_O_7_0),
    .O_7_1(n55_O_7_1),
    .O_7_2(n55_O_7_2)
  );
  Map2T_4 n56 ( // @[Top.scala 95:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0(n56_I0_0_0),
    .I0_0_1(n56_I0_0_1),
    .I0_0_2(n56_I0_0_2),
    .I0_1_0(n56_I0_1_0),
    .I0_1_1(n56_I0_1_1),
    .I0_1_2(n56_I0_1_2),
    .I0_2_0(n56_I0_2_0),
    .I0_2_1(n56_I0_2_1),
    .I0_2_2(n56_I0_2_2),
    .I0_3_0(n56_I0_3_0),
    .I0_3_1(n56_I0_3_1),
    .I0_3_2(n56_I0_3_2),
    .I0_4_0(n56_I0_4_0),
    .I0_4_1(n56_I0_4_1),
    .I0_4_2(n56_I0_4_2),
    .I0_5_0(n56_I0_5_0),
    .I0_5_1(n56_I0_5_1),
    .I0_5_2(n56_I0_5_2),
    .I0_6_0(n56_I0_6_0),
    .I0_6_1(n56_I0_6_1),
    .I0_6_2(n56_I0_6_2),
    .I0_7_0(n56_I0_7_0),
    .I0_7_1(n56_I0_7_1),
    .I0_7_2(n56_I0_7_2),
    .I1_0_0(n56_I1_0_0),
    .I1_0_1(n56_I1_0_1),
    .I1_0_2(n56_I1_0_2),
    .I1_1_0(n56_I1_1_0),
    .I1_1_1(n56_I1_1_1),
    .I1_1_2(n56_I1_1_2),
    .I1_2_0(n56_I1_2_0),
    .I1_2_1(n56_I1_2_1),
    .I1_2_2(n56_I1_2_2),
    .I1_3_0(n56_I1_3_0),
    .I1_3_1(n56_I1_3_1),
    .I1_3_2(n56_I1_3_2),
    .I1_4_0(n56_I1_4_0),
    .I1_4_1(n56_I1_4_1),
    .I1_4_2(n56_I1_4_2),
    .I1_5_0(n56_I1_5_0),
    .I1_5_1(n56_I1_5_1),
    .I1_5_2(n56_I1_5_2),
    .I1_6_0(n56_I1_6_0),
    .I1_6_1(n56_I1_6_1),
    .I1_6_2(n56_I1_6_2),
    .I1_7_0(n56_I1_7_0),
    .I1_7_1(n56_I1_7_1),
    .I1_7_2(n56_I1_7_2),
    .O_0_0_0(n56_O_0_0_0),
    .O_0_0_1(n56_O_0_0_1),
    .O_0_0_2(n56_O_0_0_2),
    .O_0_1_0(n56_O_0_1_0),
    .O_0_1_1(n56_O_0_1_1),
    .O_0_1_2(n56_O_0_1_2),
    .O_1_0_0(n56_O_1_0_0),
    .O_1_0_1(n56_O_1_0_1),
    .O_1_0_2(n56_O_1_0_2),
    .O_1_1_0(n56_O_1_1_0),
    .O_1_1_1(n56_O_1_1_1),
    .O_1_1_2(n56_O_1_1_2),
    .O_2_0_0(n56_O_2_0_0),
    .O_2_0_1(n56_O_2_0_1),
    .O_2_0_2(n56_O_2_0_2),
    .O_2_1_0(n56_O_2_1_0),
    .O_2_1_1(n56_O_2_1_1),
    .O_2_1_2(n56_O_2_1_2),
    .O_3_0_0(n56_O_3_0_0),
    .O_3_0_1(n56_O_3_0_1),
    .O_3_0_2(n56_O_3_0_2),
    .O_3_1_0(n56_O_3_1_0),
    .O_3_1_1(n56_O_3_1_1),
    .O_3_1_2(n56_O_3_1_2),
    .O_4_0_0(n56_O_4_0_0),
    .O_4_0_1(n56_O_4_0_1),
    .O_4_0_2(n56_O_4_0_2),
    .O_4_1_0(n56_O_4_1_0),
    .O_4_1_1(n56_O_4_1_1),
    .O_4_1_2(n56_O_4_1_2),
    .O_5_0_0(n56_O_5_0_0),
    .O_5_0_1(n56_O_5_0_1),
    .O_5_0_2(n56_O_5_0_2),
    .O_5_1_0(n56_O_5_1_0),
    .O_5_1_1(n56_O_5_1_1),
    .O_5_1_2(n56_O_5_1_2),
    .O_6_0_0(n56_O_6_0_0),
    .O_6_0_1(n56_O_6_0_1),
    .O_6_0_2(n56_O_6_0_2),
    .O_6_1_0(n56_O_6_1_0),
    .O_6_1_1(n56_O_6_1_1),
    .O_6_1_2(n56_O_6_1_2),
    .O_7_0_0(n56_O_7_0_0),
    .O_7_0_1(n56_O_7_0_1),
    .O_7_0_2(n56_O_7_0_2),
    .O_7_1_0(n56_O_7_1_0),
    .O_7_1_1(n56_O_7_1_1),
    .O_7_1_2(n56_O_7_1_2)
  );
  ShiftTS_2 n63 ( // @[Top.scala 99:21]
    .clock(n63_clock),
    .valid_up(n63_valid_up),
    .valid_down(n63_valid_down),
    .I_0(n63_I_0),
    .I_1(n63_I_1),
    .I_2(n63_I_2),
    .I_3(n63_I_3),
    .I_4(n63_I_4),
    .I_5(n63_I_5),
    .I_6(n63_I_6),
    .I_7(n63_I_7),
    .O_0(n63_O_0),
    .O_1(n63_O_1),
    .O_2(n63_O_2),
    .O_3(n63_O_3),
    .O_4(n63_O_4),
    .O_5(n63_O_5),
    .O_6(n63_O_6),
    .O_7(n63_O_7)
  );
  ShiftTS_2 n64 ( // @[Top.scala 102:21]
    .clock(n64_clock),
    .valid_up(n64_valid_up),
    .valid_down(n64_valid_down),
    .I_0(n64_I_0),
    .I_1(n64_I_1),
    .I_2(n64_I_2),
    .I_3(n64_I_3),
    .I_4(n64_I_4),
    .I_5(n64_I_5),
    .I_6(n64_I_6),
    .I_7(n64_I_7),
    .O_0(n64_O_0),
    .O_1(n64_O_1),
    .O_2(n64_O_2),
    .O_3(n64_O_3),
    .O_4(n64_O_4),
    .O_5(n64_O_5),
    .O_6(n64_O_6),
    .O_7(n64_O_7)
  );
  Map2T n65 ( // @[Top.scala 105:21]
    .valid_up(n65_valid_up),
    .valid_down(n65_valid_down),
    .I0_0(n65_I0_0),
    .I0_1(n65_I0_1),
    .I0_2(n65_I0_2),
    .I0_3(n65_I0_3),
    .I0_4(n65_I0_4),
    .I0_5(n65_I0_5),
    .I0_6(n65_I0_6),
    .I0_7(n65_I0_7),
    .I1_0(n65_I1_0),
    .I1_1(n65_I1_1),
    .I1_2(n65_I1_2),
    .I1_3(n65_I1_3),
    .I1_4(n65_I1_4),
    .I1_5(n65_I1_5),
    .I1_6(n65_I1_6),
    .I1_7(n65_I1_7),
    .O_0_0(n65_O_0_0),
    .O_0_1(n65_O_0_1),
    .O_1_0(n65_O_1_0),
    .O_1_1(n65_O_1_1),
    .O_2_0(n65_O_2_0),
    .O_2_1(n65_O_2_1),
    .O_3_0(n65_O_3_0),
    .O_3_1(n65_O_3_1),
    .O_4_0(n65_O_4_0),
    .O_4_1(n65_O_4_1),
    .O_5_0(n65_O_5_0),
    .O_5_1(n65_O_5_1),
    .O_6_0(n65_O_6_0),
    .O_6_1(n65_O_6_1),
    .O_7_0(n65_O_7_0),
    .O_7_1(n65_O_7_1)
  );
  Map2T_1 n72 ( // @[Top.scala 109:21]
    .valid_up(n72_valid_up),
    .valid_down(n72_valid_down),
    .I0_0_0(n72_I0_0_0),
    .I0_0_1(n72_I0_0_1),
    .I0_1_0(n72_I0_1_0),
    .I0_1_1(n72_I0_1_1),
    .I0_2_0(n72_I0_2_0),
    .I0_2_1(n72_I0_2_1),
    .I0_3_0(n72_I0_3_0),
    .I0_3_1(n72_I0_3_1),
    .I0_4_0(n72_I0_4_0),
    .I0_4_1(n72_I0_4_1),
    .I0_5_0(n72_I0_5_0),
    .I0_5_1(n72_I0_5_1),
    .I0_6_0(n72_I0_6_0),
    .I0_6_1(n72_I0_6_1),
    .I0_7_0(n72_I0_7_0),
    .I0_7_1(n72_I0_7_1),
    .I1_0(n72_I1_0),
    .I1_1(n72_I1_1),
    .I1_2(n72_I1_2),
    .I1_3(n72_I1_3),
    .I1_4(n72_I1_4),
    .I1_5(n72_I1_5),
    .I1_6(n72_I1_6),
    .I1_7(n72_I1_7),
    .O_0_0(n72_O_0_0),
    .O_0_1(n72_O_0_1),
    .O_0_2(n72_O_0_2),
    .O_1_0(n72_O_1_0),
    .O_1_1(n72_O_1_1),
    .O_1_2(n72_O_1_2),
    .O_2_0(n72_O_2_0),
    .O_2_1(n72_O_2_1),
    .O_2_2(n72_O_2_2),
    .O_3_0(n72_O_3_0),
    .O_3_1(n72_O_3_1),
    .O_3_2(n72_O_3_2),
    .O_4_0(n72_O_4_0),
    .O_4_1(n72_O_4_1),
    .O_4_2(n72_O_4_2),
    .O_5_0(n72_O_5_0),
    .O_5_1(n72_O_5_1),
    .O_5_2(n72_O_5_2),
    .O_6_0(n72_O_6_0),
    .O_6_1(n72_O_6_1),
    .O_6_2(n72_O_6_2),
    .O_7_0(n72_O_7_0),
    .O_7_1(n72_O_7_1),
    .O_7_2(n72_O_7_2)
  );
  MapT n81 ( // @[Top.scala 113:21]
    .valid_up(n81_valid_up),
    .valid_down(n81_valid_down),
    .I_0_0(n81_I_0_0),
    .I_0_1(n81_I_0_1),
    .I_0_2(n81_I_0_2),
    .I_1_0(n81_I_1_0),
    .I_1_1(n81_I_1_1),
    .I_1_2(n81_I_1_2),
    .I_2_0(n81_I_2_0),
    .I_2_1(n81_I_2_1),
    .I_2_2(n81_I_2_2),
    .I_3_0(n81_I_3_0),
    .I_3_1(n81_I_3_1),
    .I_3_2(n81_I_3_2),
    .I_4_0(n81_I_4_0),
    .I_4_1(n81_I_4_1),
    .I_4_2(n81_I_4_2),
    .I_5_0(n81_I_5_0),
    .I_5_1(n81_I_5_1),
    .I_5_2(n81_I_5_2),
    .I_6_0(n81_I_6_0),
    .I_6_1(n81_I_6_1),
    .I_6_2(n81_I_6_2),
    .I_7_0(n81_I_7_0),
    .I_7_1(n81_I_7_1),
    .I_7_2(n81_I_7_2),
    .O_0_0_0(n81_O_0_0_0),
    .O_0_0_1(n81_O_0_0_1),
    .O_0_0_2(n81_O_0_0_2),
    .O_1_0_0(n81_O_1_0_0),
    .O_1_0_1(n81_O_1_0_1),
    .O_1_0_2(n81_O_1_0_2),
    .O_2_0_0(n81_O_2_0_0),
    .O_2_0_1(n81_O_2_0_1),
    .O_2_0_2(n81_O_2_0_2),
    .O_3_0_0(n81_O_3_0_0),
    .O_3_0_1(n81_O_3_0_1),
    .O_3_0_2(n81_O_3_0_2),
    .O_4_0_0(n81_O_4_0_0),
    .O_4_0_1(n81_O_4_0_1),
    .O_4_0_2(n81_O_4_0_2),
    .O_5_0_0(n81_O_5_0_0),
    .O_5_0_1(n81_O_5_0_1),
    .O_5_0_2(n81_O_5_0_2),
    .O_6_0_0(n81_O_6_0_0),
    .O_6_0_1(n81_O_6_0_1),
    .O_6_0_2(n81_O_6_0_2),
    .O_7_0_0(n81_O_7_0_0),
    .O_7_0_1(n81_O_7_0_1),
    .O_7_0_2(n81_O_7_0_2)
  );
  MapT_1 n88 ( // @[Top.scala 116:21]
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_0_0_1(n88_I_0_0_1),
    .I_0_0_2(n88_I_0_0_2),
    .I_1_0_0(n88_I_1_0_0),
    .I_1_0_1(n88_I_1_0_1),
    .I_1_0_2(n88_I_1_0_2),
    .I_2_0_0(n88_I_2_0_0),
    .I_2_0_1(n88_I_2_0_1),
    .I_2_0_2(n88_I_2_0_2),
    .I_3_0_0(n88_I_3_0_0),
    .I_3_0_1(n88_I_3_0_1),
    .I_3_0_2(n88_I_3_0_2),
    .I_4_0_0(n88_I_4_0_0),
    .I_4_0_1(n88_I_4_0_1),
    .I_4_0_2(n88_I_4_0_2),
    .I_5_0_0(n88_I_5_0_0),
    .I_5_0_1(n88_I_5_0_1),
    .I_5_0_2(n88_I_5_0_2),
    .I_6_0_0(n88_I_6_0_0),
    .I_6_0_1(n88_I_6_0_1),
    .I_6_0_2(n88_I_6_0_2),
    .I_7_0_0(n88_I_7_0_0),
    .I_7_0_1(n88_I_7_0_1),
    .I_7_0_2(n88_I_7_0_2),
    .O_0_0(n88_O_0_0),
    .O_0_1(n88_O_0_1),
    .O_0_2(n88_O_0_2),
    .O_1_0(n88_O_1_0),
    .O_1_1(n88_O_1_1),
    .O_1_2(n88_O_1_2),
    .O_2_0(n88_O_2_0),
    .O_2_1(n88_O_2_1),
    .O_2_2(n88_O_2_2),
    .O_3_0(n88_O_3_0),
    .O_3_1(n88_O_3_1),
    .O_3_2(n88_O_3_2),
    .O_4_0(n88_O_4_0),
    .O_4_1(n88_O_4_1),
    .O_4_2(n88_O_4_2),
    .O_5_0(n88_O_5_0),
    .O_5_1(n88_O_5_1),
    .O_5_2(n88_O_5_2),
    .O_6_0(n88_O_6_0),
    .O_6_1(n88_O_6_1),
    .O_6_2(n88_O_6_2),
    .O_7_0(n88_O_7_0),
    .O_7_1(n88_O_7_1),
    .O_7_2(n88_O_7_2)
  );
  Map2T_7 n89 ( // @[Top.scala 119:21]
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I0_0_0_0(n89_I0_0_0_0),
    .I0_0_0_1(n89_I0_0_0_1),
    .I0_0_0_2(n89_I0_0_0_2),
    .I0_0_1_0(n89_I0_0_1_0),
    .I0_0_1_1(n89_I0_0_1_1),
    .I0_0_1_2(n89_I0_0_1_2),
    .I0_1_0_0(n89_I0_1_0_0),
    .I0_1_0_1(n89_I0_1_0_1),
    .I0_1_0_2(n89_I0_1_0_2),
    .I0_1_1_0(n89_I0_1_1_0),
    .I0_1_1_1(n89_I0_1_1_1),
    .I0_1_1_2(n89_I0_1_1_2),
    .I0_2_0_0(n89_I0_2_0_0),
    .I0_2_0_1(n89_I0_2_0_1),
    .I0_2_0_2(n89_I0_2_0_2),
    .I0_2_1_0(n89_I0_2_1_0),
    .I0_2_1_1(n89_I0_2_1_1),
    .I0_2_1_2(n89_I0_2_1_2),
    .I0_3_0_0(n89_I0_3_0_0),
    .I0_3_0_1(n89_I0_3_0_1),
    .I0_3_0_2(n89_I0_3_0_2),
    .I0_3_1_0(n89_I0_3_1_0),
    .I0_3_1_1(n89_I0_3_1_1),
    .I0_3_1_2(n89_I0_3_1_2),
    .I0_4_0_0(n89_I0_4_0_0),
    .I0_4_0_1(n89_I0_4_0_1),
    .I0_4_0_2(n89_I0_4_0_2),
    .I0_4_1_0(n89_I0_4_1_0),
    .I0_4_1_1(n89_I0_4_1_1),
    .I0_4_1_2(n89_I0_4_1_2),
    .I0_5_0_0(n89_I0_5_0_0),
    .I0_5_0_1(n89_I0_5_0_1),
    .I0_5_0_2(n89_I0_5_0_2),
    .I0_5_1_0(n89_I0_5_1_0),
    .I0_5_1_1(n89_I0_5_1_1),
    .I0_5_1_2(n89_I0_5_1_2),
    .I0_6_0_0(n89_I0_6_0_0),
    .I0_6_0_1(n89_I0_6_0_1),
    .I0_6_0_2(n89_I0_6_0_2),
    .I0_6_1_0(n89_I0_6_1_0),
    .I0_6_1_1(n89_I0_6_1_1),
    .I0_6_1_2(n89_I0_6_1_2),
    .I0_7_0_0(n89_I0_7_0_0),
    .I0_7_0_1(n89_I0_7_0_1),
    .I0_7_0_2(n89_I0_7_0_2),
    .I0_7_1_0(n89_I0_7_1_0),
    .I0_7_1_1(n89_I0_7_1_1),
    .I0_7_1_2(n89_I0_7_1_2),
    .I1_0_0(n89_I1_0_0),
    .I1_0_1(n89_I1_0_1),
    .I1_0_2(n89_I1_0_2),
    .I1_1_0(n89_I1_1_0),
    .I1_1_1(n89_I1_1_1),
    .I1_1_2(n89_I1_1_2),
    .I1_2_0(n89_I1_2_0),
    .I1_2_1(n89_I1_2_1),
    .I1_2_2(n89_I1_2_2),
    .I1_3_0(n89_I1_3_0),
    .I1_3_1(n89_I1_3_1),
    .I1_3_2(n89_I1_3_2),
    .I1_4_0(n89_I1_4_0),
    .I1_4_1(n89_I1_4_1),
    .I1_4_2(n89_I1_4_2),
    .I1_5_0(n89_I1_5_0),
    .I1_5_1(n89_I1_5_1),
    .I1_5_2(n89_I1_5_2),
    .I1_6_0(n89_I1_6_0),
    .I1_6_1(n89_I1_6_1),
    .I1_6_2(n89_I1_6_2),
    .I1_7_0(n89_I1_7_0),
    .I1_7_1(n89_I1_7_1),
    .I1_7_2(n89_I1_7_2),
    .O_0_0_0(n89_O_0_0_0),
    .O_0_0_1(n89_O_0_0_1),
    .O_0_0_2(n89_O_0_0_2),
    .O_0_1_0(n89_O_0_1_0),
    .O_0_1_1(n89_O_0_1_1),
    .O_0_1_2(n89_O_0_1_2),
    .O_0_2_0(n89_O_0_2_0),
    .O_0_2_1(n89_O_0_2_1),
    .O_0_2_2(n89_O_0_2_2),
    .O_1_0_0(n89_O_1_0_0),
    .O_1_0_1(n89_O_1_0_1),
    .O_1_0_2(n89_O_1_0_2),
    .O_1_1_0(n89_O_1_1_0),
    .O_1_1_1(n89_O_1_1_1),
    .O_1_1_2(n89_O_1_1_2),
    .O_1_2_0(n89_O_1_2_0),
    .O_1_2_1(n89_O_1_2_1),
    .O_1_2_2(n89_O_1_2_2),
    .O_2_0_0(n89_O_2_0_0),
    .O_2_0_1(n89_O_2_0_1),
    .O_2_0_2(n89_O_2_0_2),
    .O_2_1_0(n89_O_2_1_0),
    .O_2_1_1(n89_O_2_1_1),
    .O_2_1_2(n89_O_2_1_2),
    .O_2_2_0(n89_O_2_2_0),
    .O_2_2_1(n89_O_2_2_1),
    .O_2_2_2(n89_O_2_2_2),
    .O_3_0_0(n89_O_3_0_0),
    .O_3_0_1(n89_O_3_0_1),
    .O_3_0_2(n89_O_3_0_2),
    .O_3_1_0(n89_O_3_1_0),
    .O_3_1_1(n89_O_3_1_1),
    .O_3_1_2(n89_O_3_1_2),
    .O_3_2_0(n89_O_3_2_0),
    .O_3_2_1(n89_O_3_2_1),
    .O_3_2_2(n89_O_3_2_2),
    .O_4_0_0(n89_O_4_0_0),
    .O_4_0_1(n89_O_4_0_1),
    .O_4_0_2(n89_O_4_0_2),
    .O_4_1_0(n89_O_4_1_0),
    .O_4_1_1(n89_O_4_1_1),
    .O_4_1_2(n89_O_4_1_2),
    .O_4_2_0(n89_O_4_2_0),
    .O_4_2_1(n89_O_4_2_1),
    .O_4_2_2(n89_O_4_2_2),
    .O_5_0_0(n89_O_5_0_0),
    .O_5_0_1(n89_O_5_0_1),
    .O_5_0_2(n89_O_5_0_2),
    .O_5_1_0(n89_O_5_1_0),
    .O_5_1_1(n89_O_5_1_1),
    .O_5_1_2(n89_O_5_1_2),
    .O_5_2_0(n89_O_5_2_0),
    .O_5_2_1(n89_O_5_2_1),
    .O_5_2_2(n89_O_5_2_2),
    .O_6_0_0(n89_O_6_0_0),
    .O_6_0_1(n89_O_6_0_1),
    .O_6_0_2(n89_O_6_0_2),
    .O_6_1_0(n89_O_6_1_0),
    .O_6_1_1(n89_O_6_1_1),
    .O_6_1_2(n89_O_6_1_2),
    .O_6_2_0(n89_O_6_2_0),
    .O_6_2_1(n89_O_6_2_1),
    .O_6_2_2(n89_O_6_2_2),
    .O_7_0_0(n89_O_7_0_0),
    .O_7_0_1(n89_O_7_0_1),
    .O_7_0_2(n89_O_7_0_2),
    .O_7_1_0(n89_O_7_1_0),
    .O_7_1_1(n89_O_7_1_1),
    .O_7_1_2(n89_O_7_1_2),
    .O_7_2_0(n89_O_7_2_0),
    .O_7_2_1(n89_O_7_2_1),
    .O_7_2_2(n89_O_7_2_2)
  );
  MapT_6 n98 ( // @[Top.scala 123:21]
    .valid_up(n98_valid_up),
    .valid_down(n98_valid_down),
    .I_0_0_0(n98_I_0_0_0),
    .I_0_0_1(n98_I_0_0_1),
    .I_0_0_2(n98_I_0_0_2),
    .I_0_1_0(n98_I_0_1_0),
    .I_0_1_1(n98_I_0_1_1),
    .I_0_1_2(n98_I_0_1_2),
    .I_0_2_0(n98_I_0_2_0),
    .I_0_2_1(n98_I_0_2_1),
    .I_0_2_2(n98_I_0_2_2),
    .I_1_0_0(n98_I_1_0_0),
    .I_1_0_1(n98_I_1_0_1),
    .I_1_0_2(n98_I_1_0_2),
    .I_1_1_0(n98_I_1_1_0),
    .I_1_1_1(n98_I_1_1_1),
    .I_1_1_2(n98_I_1_1_2),
    .I_1_2_0(n98_I_1_2_0),
    .I_1_2_1(n98_I_1_2_1),
    .I_1_2_2(n98_I_1_2_2),
    .I_2_0_0(n98_I_2_0_0),
    .I_2_0_1(n98_I_2_0_1),
    .I_2_0_2(n98_I_2_0_2),
    .I_2_1_0(n98_I_2_1_0),
    .I_2_1_1(n98_I_2_1_1),
    .I_2_1_2(n98_I_2_1_2),
    .I_2_2_0(n98_I_2_2_0),
    .I_2_2_1(n98_I_2_2_1),
    .I_2_2_2(n98_I_2_2_2),
    .I_3_0_0(n98_I_3_0_0),
    .I_3_0_1(n98_I_3_0_1),
    .I_3_0_2(n98_I_3_0_2),
    .I_3_1_0(n98_I_3_1_0),
    .I_3_1_1(n98_I_3_1_1),
    .I_3_1_2(n98_I_3_1_2),
    .I_3_2_0(n98_I_3_2_0),
    .I_3_2_1(n98_I_3_2_1),
    .I_3_2_2(n98_I_3_2_2),
    .I_4_0_0(n98_I_4_0_0),
    .I_4_0_1(n98_I_4_0_1),
    .I_4_0_2(n98_I_4_0_2),
    .I_4_1_0(n98_I_4_1_0),
    .I_4_1_1(n98_I_4_1_1),
    .I_4_1_2(n98_I_4_1_2),
    .I_4_2_0(n98_I_4_2_0),
    .I_4_2_1(n98_I_4_2_1),
    .I_4_2_2(n98_I_4_2_2),
    .I_5_0_0(n98_I_5_0_0),
    .I_5_0_1(n98_I_5_0_1),
    .I_5_0_2(n98_I_5_0_2),
    .I_5_1_0(n98_I_5_1_0),
    .I_5_1_1(n98_I_5_1_1),
    .I_5_1_2(n98_I_5_1_2),
    .I_5_2_0(n98_I_5_2_0),
    .I_5_2_1(n98_I_5_2_1),
    .I_5_2_2(n98_I_5_2_2),
    .I_6_0_0(n98_I_6_0_0),
    .I_6_0_1(n98_I_6_0_1),
    .I_6_0_2(n98_I_6_0_2),
    .I_6_1_0(n98_I_6_1_0),
    .I_6_1_1(n98_I_6_1_1),
    .I_6_1_2(n98_I_6_1_2),
    .I_6_2_0(n98_I_6_2_0),
    .I_6_2_1(n98_I_6_2_1),
    .I_6_2_2(n98_I_6_2_2),
    .I_7_0_0(n98_I_7_0_0),
    .I_7_0_1(n98_I_7_0_1),
    .I_7_0_2(n98_I_7_0_2),
    .I_7_1_0(n98_I_7_1_0),
    .I_7_1_1(n98_I_7_1_1),
    .I_7_1_2(n98_I_7_1_2),
    .I_7_2_0(n98_I_7_2_0),
    .I_7_2_1(n98_I_7_2_1),
    .I_7_2_2(n98_I_7_2_2),
    .O_0_0_0_0(n98_O_0_0_0_0),
    .O_0_0_0_1(n98_O_0_0_0_1),
    .O_0_0_0_2(n98_O_0_0_0_2),
    .O_0_0_1_0(n98_O_0_0_1_0),
    .O_0_0_1_1(n98_O_0_0_1_1),
    .O_0_0_1_2(n98_O_0_0_1_2),
    .O_0_0_2_0(n98_O_0_0_2_0),
    .O_0_0_2_1(n98_O_0_0_2_1),
    .O_0_0_2_2(n98_O_0_0_2_2),
    .O_1_0_0_0(n98_O_1_0_0_0),
    .O_1_0_0_1(n98_O_1_0_0_1),
    .O_1_0_0_2(n98_O_1_0_0_2),
    .O_1_0_1_0(n98_O_1_0_1_0),
    .O_1_0_1_1(n98_O_1_0_1_1),
    .O_1_0_1_2(n98_O_1_0_1_2),
    .O_1_0_2_0(n98_O_1_0_2_0),
    .O_1_0_2_1(n98_O_1_0_2_1),
    .O_1_0_2_2(n98_O_1_0_2_2),
    .O_2_0_0_0(n98_O_2_0_0_0),
    .O_2_0_0_1(n98_O_2_0_0_1),
    .O_2_0_0_2(n98_O_2_0_0_2),
    .O_2_0_1_0(n98_O_2_0_1_0),
    .O_2_0_1_1(n98_O_2_0_1_1),
    .O_2_0_1_2(n98_O_2_0_1_2),
    .O_2_0_2_0(n98_O_2_0_2_0),
    .O_2_0_2_1(n98_O_2_0_2_1),
    .O_2_0_2_2(n98_O_2_0_2_2),
    .O_3_0_0_0(n98_O_3_0_0_0),
    .O_3_0_0_1(n98_O_3_0_0_1),
    .O_3_0_0_2(n98_O_3_0_0_2),
    .O_3_0_1_0(n98_O_3_0_1_0),
    .O_3_0_1_1(n98_O_3_0_1_1),
    .O_3_0_1_2(n98_O_3_0_1_2),
    .O_3_0_2_0(n98_O_3_0_2_0),
    .O_3_0_2_1(n98_O_3_0_2_1),
    .O_3_0_2_2(n98_O_3_0_2_2),
    .O_4_0_0_0(n98_O_4_0_0_0),
    .O_4_0_0_1(n98_O_4_0_0_1),
    .O_4_0_0_2(n98_O_4_0_0_2),
    .O_4_0_1_0(n98_O_4_0_1_0),
    .O_4_0_1_1(n98_O_4_0_1_1),
    .O_4_0_1_2(n98_O_4_0_1_2),
    .O_4_0_2_0(n98_O_4_0_2_0),
    .O_4_0_2_1(n98_O_4_0_2_1),
    .O_4_0_2_2(n98_O_4_0_2_2),
    .O_5_0_0_0(n98_O_5_0_0_0),
    .O_5_0_0_1(n98_O_5_0_0_1),
    .O_5_0_0_2(n98_O_5_0_0_2),
    .O_5_0_1_0(n98_O_5_0_1_0),
    .O_5_0_1_1(n98_O_5_0_1_1),
    .O_5_0_1_2(n98_O_5_0_1_2),
    .O_5_0_2_0(n98_O_5_0_2_0),
    .O_5_0_2_1(n98_O_5_0_2_1),
    .O_5_0_2_2(n98_O_5_0_2_2),
    .O_6_0_0_0(n98_O_6_0_0_0),
    .O_6_0_0_1(n98_O_6_0_0_1),
    .O_6_0_0_2(n98_O_6_0_0_2),
    .O_6_0_1_0(n98_O_6_0_1_0),
    .O_6_0_1_1(n98_O_6_0_1_1),
    .O_6_0_1_2(n98_O_6_0_1_2),
    .O_6_0_2_0(n98_O_6_0_2_0),
    .O_6_0_2_1(n98_O_6_0_2_1),
    .O_6_0_2_2(n98_O_6_0_2_2),
    .O_7_0_0_0(n98_O_7_0_0_0),
    .O_7_0_0_1(n98_O_7_0_0_1),
    .O_7_0_0_2(n98_O_7_0_0_2),
    .O_7_0_1_0(n98_O_7_0_1_0),
    .O_7_0_1_1(n98_O_7_0_1_1),
    .O_7_0_1_2(n98_O_7_0_1_2),
    .O_7_0_2_0(n98_O_7_0_2_0),
    .O_7_0_2_1(n98_O_7_0_2_1),
    .O_7_0_2_2(n98_O_7_0_2_2)
  );
  MapT_7 n105 ( // @[Top.scala 126:22]
    .valid_up(n105_valid_up),
    .valid_down(n105_valid_down),
    .I_0_0_0_0(n105_I_0_0_0_0),
    .I_0_0_0_1(n105_I_0_0_0_1),
    .I_0_0_0_2(n105_I_0_0_0_2),
    .I_0_0_1_0(n105_I_0_0_1_0),
    .I_0_0_1_1(n105_I_0_0_1_1),
    .I_0_0_1_2(n105_I_0_0_1_2),
    .I_0_0_2_0(n105_I_0_0_2_0),
    .I_0_0_2_1(n105_I_0_0_2_1),
    .I_0_0_2_2(n105_I_0_0_2_2),
    .I_1_0_0_0(n105_I_1_0_0_0),
    .I_1_0_0_1(n105_I_1_0_0_1),
    .I_1_0_0_2(n105_I_1_0_0_2),
    .I_1_0_1_0(n105_I_1_0_1_0),
    .I_1_0_1_1(n105_I_1_0_1_1),
    .I_1_0_1_2(n105_I_1_0_1_2),
    .I_1_0_2_0(n105_I_1_0_2_0),
    .I_1_0_2_1(n105_I_1_0_2_1),
    .I_1_0_2_2(n105_I_1_0_2_2),
    .I_2_0_0_0(n105_I_2_0_0_0),
    .I_2_0_0_1(n105_I_2_0_0_1),
    .I_2_0_0_2(n105_I_2_0_0_2),
    .I_2_0_1_0(n105_I_2_0_1_0),
    .I_2_0_1_1(n105_I_2_0_1_1),
    .I_2_0_1_2(n105_I_2_0_1_2),
    .I_2_0_2_0(n105_I_2_0_2_0),
    .I_2_0_2_1(n105_I_2_0_2_1),
    .I_2_0_2_2(n105_I_2_0_2_2),
    .I_3_0_0_0(n105_I_3_0_0_0),
    .I_3_0_0_1(n105_I_3_0_0_1),
    .I_3_0_0_2(n105_I_3_0_0_2),
    .I_3_0_1_0(n105_I_3_0_1_0),
    .I_3_0_1_1(n105_I_3_0_1_1),
    .I_3_0_1_2(n105_I_3_0_1_2),
    .I_3_0_2_0(n105_I_3_0_2_0),
    .I_3_0_2_1(n105_I_3_0_2_1),
    .I_3_0_2_2(n105_I_3_0_2_2),
    .I_4_0_0_0(n105_I_4_0_0_0),
    .I_4_0_0_1(n105_I_4_0_0_1),
    .I_4_0_0_2(n105_I_4_0_0_2),
    .I_4_0_1_0(n105_I_4_0_1_0),
    .I_4_0_1_1(n105_I_4_0_1_1),
    .I_4_0_1_2(n105_I_4_0_1_2),
    .I_4_0_2_0(n105_I_4_0_2_0),
    .I_4_0_2_1(n105_I_4_0_2_1),
    .I_4_0_2_2(n105_I_4_0_2_2),
    .I_5_0_0_0(n105_I_5_0_0_0),
    .I_5_0_0_1(n105_I_5_0_0_1),
    .I_5_0_0_2(n105_I_5_0_0_2),
    .I_5_0_1_0(n105_I_5_0_1_0),
    .I_5_0_1_1(n105_I_5_0_1_1),
    .I_5_0_1_2(n105_I_5_0_1_2),
    .I_5_0_2_0(n105_I_5_0_2_0),
    .I_5_0_2_1(n105_I_5_0_2_1),
    .I_5_0_2_2(n105_I_5_0_2_2),
    .I_6_0_0_0(n105_I_6_0_0_0),
    .I_6_0_0_1(n105_I_6_0_0_1),
    .I_6_0_0_2(n105_I_6_0_0_2),
    .I_6_0_1_0(n105_I_6_0_1_0),
    .I_6_0_1_1(n105_I_6_0_1_1),
    .I_6_0_1_2(n105_I_6_0_1_2),
    .I_6_0_2_0(n105_I_6_0_2_0),
    .I_6_0_2_1(n105_I_6_0_2_1),
    .I_6_0_2_2(n105_I_6_0_2_2),
    .I_7_0_0_0(n105_I_7_0_0_0),
    .I_7_0_0_1(n105_I_7_0_0_1),
    .I_7_0_0_2(n105_I_7_0_0_2),
    .I_7_0_1_0(n105_I_7_0_1_0),
    .I_7_0_1_1(n105_I_7_0_1_1),
    .I_7_0_1_2(n105_I_7_0_1_2),
    .I_7_0_2_0(n105_I_7_0_2_0),
    .I_7_0_2_1(n105_I_7_0_2_1),
    .I_7_0_2_2(n105_I_7_0_2_2),
    .O_0_0_0(n105_O_0_0_0),
    .O_0_0_1(n105_O_0_0_1),
    .O_0_0_2(n105_O_0_0_2),
    .O_0_1_0(n105_O_0_1_0),
    .O_0_1_1(n105_O_0_1_1),
    .O_0_1_2(n105_O_0_1_2),
    .O_0_2_0(n105_O_0_2_0),
    .O_0_2_1(n105_O_0_2_1),
    .O_0_2_2(n105_O_0_2_2),
    .O_1_0_0(n105_O_1_0_0),
    .O_1_0_1(n105_O_1_0_1),
    .O_1_0_2(n105_O_1_0_2),
    .O_1_1_0(n105_O_1_1_0),
    .O_1_1_1(n105_O_1_1_1),
    .O_1_1_2(n105_O_1_1_2),
    .O_1_2_0(n105_O_1_2_0),
    .O_1_2_1(n105_O_1_2_1),
    .O_1_2_2(n105_O_1_2_2),
    .O_2_0_0(n105_O_2_0_0),
    .O_2_0_1(n105_O_2_0_1),
    .O_2_0_2(n105_O_2_0_2),
    .O_2_1_0(n105_O_2_1_0),
    .O_2_1_1(n105_O_2_1_1),
    .O_2_1_2(n105_O_2_1_2),
    .O_2_2_0(n105_O_2_2_0),
    .O_2_2_1(n105_O_2_2_1),
    .O_2_2_2(n105_O_2_2_2),
    .O_3_0_0(n105_O_3_0_0),
    .O_3_0_1(n105_O_3_0_1),
    .O_3_0_2(n105_O_3_0_2),
    .O_3_1_0(n105_O_3_1_0),
    .O_3_1_1(n105_O_3_1_1),
    .O_3_1_2(n105_O_3_1_2),
    .O_3_2_0(n105_O_3_2_0),
    .O_3_2_1(n105_O_3_2_1),
    .O_3_2_2(n105_O_3_2_2),
    .O_4_0_0(n105_O_4_0_0),
    .O_4_0_1(n105_O_4_0_1),
    .O_4_0_2(n105_O_4_0_2),
    .O_4_1_0(n105_O_4_1_0),
    .O_4_1_1(n105_O_4_1_1),
    .O_4_1_2(n105_O_4_1_2),
    .O_4_2_0(n105_O_4_2_0),
    .O_4_2_1(n105_O_4_2_1),
    .O_4_2_2(n105_O_4_2_2),
    .O_5_0_0(n105_O_5_0_0),
    .O_5_0_1(n105_O_5_0_1),
    .O_5_0_2(n105_O_5_0_2),
    .O_5_1_0(n105_O_5_1_0),
    .O_5_1_1(n105_O_5_1_1),
    .O_5_1_2(n105_O_5_1_2),
    .O_5_2_0(n105_O_5_2_0),
    .O_5_2_1(n105_O_5_2_1),
    .O_5_2_2(n105_O_5_2_2),
    .O_6_0_0(n105_O_6_0_0),
    .O_6_0_1(n105_O_6_0_1),
    .O_6_0_2(n105_O_6_0_2),
    .O_6_1_0(n105_O_6_1_0),
    .O_6_1_1(n105_O_6_1_1),
    .O_6_1_2(n105_O_6_1_2),
    .O_6_2_0(n105_O_6_2_0),
    .O_6_2_1(n105_O_6_2_1),
    .O_6_2_2(n105_O_6_2_2),
    .O_7_0_0(n105_O_7_0_0),
    .O_7_0_1(n105_O_7_0_1),
    .O_7_0_2(n105_O_7_0_2),
    .O_7_1_0(n105_O_7_1_0),
    .O_7_1_1(n105_O_7_1_1),
    .O_7_1_2(n105_O_7_1_2),
    .O_7_2_0(n105_O_7_2_0),
    .O_7_2_1(n105_O_7_2_1),
    .O_7_2_2(n105_O_7_2_2)
  );
  MapT_8 n147 ( // @[Top.scala 129:22]
    .clock(n147_clock),
    .reset(n147_reset),
    .valid_up(n147_valid_up),
    .valid_down(n147_valid_down),
    .I_0_0_0(n147_I_0_0_0),
    .I_0_0_1(n147_I_0_0_1),
    .I_0_0_2(n147_I_0_0_2),
    .I_0_1_0(n147_I_0_1_0),
    .I_0_1_1(n147_I_0_1_1),
    .I_0_1_2(n147_I_0_1_2),
    .I_0_2_0(n147_I_0_2_0),
    .I_0_2_1(n147_I_0_2_1),
    .I_0_2_2(n147_I_0_2_2),
    .I_1_0_0(n147_I_1_0_0),
    .I_1_0_1(n147_I_1_0_1),
    .I_1_0_2(n147_I_1_0_2),
    .I_1_1_0(n147_I_1_1_0),
    .I_1_1_1(n147_I_1_1_1),
    .I_1_1_2(n147_I_1_1_2),
    .I_1_2_0(n147_I_1_2_0),
    .I_1_2_1(n147_I_1_2_1),
    .I_1_2_2(n147_I_1_2_2),
    .I_2_0_0(n147_I_2_0_0),
    .I_2_0_1(n147_I_2_0_1),
    .I_2_0_2(n147_I_2_0_2),
    .I_2_1_0(n147_I_2_1_0),
    .I_2_1_1(n147_I_2_1_1),
    .I_2_1_2(n147_I_2_1_2),
    .I_2_2_0(n147_I_2_2_0),
    .I_2_2_1(n147_I_2_2_1),
    .I_2_2_2(n147_I_2_2_2),
    .I_3_0_0(n147_I_3_0_0),
    .I_3_0_1(n147_I_3_0_1),
    .I_3_0_2(n147_I_3_0_2),
    .I_3_1_0(n147_I_3_1_0),
    .I_3_1_1(n147_I_3_1_1),
    .I_3_1_2(n147_I_3_1_2),
    .I_3_2_0(n147_I_3_2_0),
    .I_3_2_1(n147_I_3_2_1),
    .I_3_2_2(n147_I_3_2_2),
    .I_4_0_0(n147_I_4_0_0),
    .I_4_0_1(n147_I_4_0_1),
    .I_4_0_2(n147_I_4_0_2),
    .I_4_1_0(n147_I_4_1_0),
    .I_4_1_1(n147_I_4_1_1),
    .I_4_1_2(n147_I_4_1_2),
    .I_4_2_0(n147_I_4_2_0),
    .I_4_2_1(n147_I_4_2_1),
    .I_4_2_2(n147_I_4_2_2),
    .I_5_0_0(n147_I_5_0_0),
    .I_5_0_1(n147_I_5_0_1),
    .I_5_0_2(n147_I_5_0_2),
    .I_5_1_0(n147_I_5_1_0),
    .I_5_1_1(n147_I_5_1_1),
    .I_5_1_2(n147_I_5_1_2),
    .I_5_2_0(n147_I_5_2_0),
    .I_5_2_1(n147_I_5_2_1),
    .I_5_2_2(n147_I_5_2_2),
    .I_6_0_0(n147_I_6_0_0),
    .I_6_0_1(n147_I_6_0_1),
    .I_6_0_2(n147_I_6_0_2),
    .I_6_1_0(n147_I_6_1_0),
    .I_6_1_1(n147_I_6_1_1),
    .I_6_1_2(n147_I_6_1_2),
    .I_6_2_0(n147_I_6_2_0),
    .I_6_2_1(n147_I_6_2_1),
    .I_6_2_2(n147_I_6_2_2),
    .I_7_0_0(n147_I_7_0_0),
    .I_7_0_1(n147_I_7_0_1),
    .I_7_0_2(n147_I_7_0_2),
    .I_7_1_0(n147_I_7_1_0),
    .I_7_1_1(n147_I_7_1_1),
    .I_7_1_2(n147_I_7_1_2),
    .I_7_2_0(n147_I_7_2_0),
    .I_7_2_1(n147_I_7_2_1),
    .I_7_2_2(n147_I_7_2_2),
    .O_0_0_0(n147_O_0_0_0),
    .O_1_0_0(n147_O_1_0_0),
    .O_2_0_0(n147_O_2_0_0),
    .O_3_0_0(n147_O_3_0_0),
    .O_4_0_0(n147_O_4_0_0),
    .O_5_0_0(n147_O_5_0_0),
    .O_6_0_0(n147_O_6_0_0),
    .O_7_0_0(n147_O_7_0_0)
  );
  Passthrough n148 ( // @[Top.scala 132:22]
    .valid_up(n148_valid_up),
    .valid_down(n148_valid_down),
    .I_0_0_0(n148_I_0_0_0),
    .I_1_0_0(n148_I_1_0_0),
    .I_2_0_0(n148_I_2_0_0),
    .I_3_0_0(n148_I_3_0_0),
    .I_4_0_0(n148_I_4_0_0),
    .I_5_0_0(n148_I_5_0_0),
    .I_6_0_0(n148_I_6_0_0),
    .I_7_0_0(n148_I_7_0_0),
    .O_0_0(n148_O_0_0),
    .O_1_0(n148_O_1_0),
    .O_2_0(n148_O_2_0),
    .O_3_0(n148_O_3_0),
    .O_4_0(n148_O_4_0),
    .O_5_0(n148_O_5_0),
    .O_6_0(n148_O_6_0),
    .O_7_0(n148_O_7_0)
  );
  Passthrough_1 n149 ( // @[Top.scala 135:22]
    .valid_up(n149_valid_up),
    .valid_down(n149_valid_down),
    .I_0_0(n149_I_0_0),
    .I_1_0(n149_I_1_0),
    .I_2_0(n149_I_2_0),
    .I_3_0(n149_I_3_0),
    .I_4_0(n149_I_4_0),
    .I_5_0(n149_I_5_0),
    .I_6_0(n149_I_6_0),
    .I_7_0(n149_I_7_0),
    .O_0(n149_O_0),
    .O_1(n149_O_1),
    .O_2(n149_O_2),
    .O_3(n149_O_3),
    .O_4(n149_O_4),
    .O_5(n149_O_5),
    .O_6(n149_O_6),
    .O_7(n149_O_7)
  );
  FIFO n150 ( // @[Top.scala 138:22]
    .clock(n150_clock),
    .reset(n150_reset),
    .valid_up(n150_valid_up),
    .valid_down(n150_valid_down),
    .I_0(n150_I_0),
    .I_1(n150_I_1),
    .I_2(n150_I_2),
    .I_3(n150_I_3),
    .I_4(n150_I_4),
    .I_5(n150_I_5),
    .I_6(n150_I_6),
    .I_7(n150_I_7),
    .O_0(n150_O_0),
    .O_1(n150_O_1),
    .O_2(n150_O_2),
    .O_3(n150_O_3),
    .O_4(n150_O_4),
    .O_5(n150_O_5),
    .O_6(n150_O_6),
    .O_7(n150_O_7)
  );
  FIFO n151 ( // @[Top.scala 141:22]
    .clock(n151_clock),
    .reset(n151_reset),
    .valid_up(n151_valid_up),
    .valid_down(n151_valid_down),
    .I_0(n151_I_0),
    .I_1(n151_I_1),
    .I_2(n151_I_2),
    .I_3(n151_I_3),
    .I_4(n151_I_4),
    .I_5(n151_I_5),
    .I_6(n151_I_6),
    .I_7(n151_I_7),
    .O_0(n151_O_0),
    .O_1(n151_O_1),
    .O_2(n151_O_2),
    .O_3(n151_O_3),
    .O_4(n151_O_4),
    .O_5(n151_O_5),
    .O_6(n151_O_6),
    .O_7(n151_O_7)
  );
  FIFO n152 ( // @[Top.scala 144:22]
    .clock(n152_clock),
    .reset(n152_reset),
    .valid_up(n152_valid_up),
    .valid_down(n152_valid_down),
    .I_0(n152_I_0),
    .I_1(n152_I_1),
    .I_2(n152_I_2),
    .I_3(n152_I_3),
    .I_4(n152_I_4),
    .I_5(n152_I_5),
    .I_6(n152_I_6),
    .I_7(n152_I_7),
    .O_0(n152_O_0),
    .O_1(n152_O_1),
    .O_2(n152_O_2),
    .O_3(n152_O_3),
    .O_4(n152_O_4),
    .O_5(n152_O_5),
    .O_6(n152_O_6),
    .O_7(n152_O_7)
  );
  assign valid_down = n152_valid_down; // @[Top.scala 148:16]
  assign O_0 = n152_O_0; // @[Top.scala 147:7]
  assign O_1 = n152_O_1; // @[Top.scala 147:7]
  assign O_2 = n152_O_2; // @[Top.scala 147:7]
  assign O_3 = n152_O_3; // @[Top.scala 147:7]
  assign O_4 = n152_O_4; // @[Top.scala 147:7]
  assign O_5 = n152_O_5; // @[Top.scala 147:7]
  assign O_6 = n152_O_6; // @[Top.scala 147:7]
  assign O_7 = n152_O_7; // @[Top.scala 147:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 48:17]
  assign n1_I_0 = I_0; // @[Top.scala 47:10]
  assign n1_I_1 = I_1; // @[Top.scala 47:10]
  assign n1_I_2 = I_2; // @[Top.scala 47:10]
  assign n1_I_3 = I_3; // @[Top.scala 47:10]
  assign n1_I_4 = I_4; // @[Top.scala 47:10]
  assign n1_I_5 = I_5; // @[Top.scala 47:10]
  assign n1_I_6 = I_6; // @[Top.scala 47:10]
  assign n1_I_7 = I_7; // @[Top.scala 47:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 51:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 50:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 50:10]
  assign n2_I_2 = n1_O_2; // @[Top.scala 50:10]
  assign n2_I_3 = n1_O_3; // @[Top.scala 50:10]
  assign n2_I_4 = n1_O_4; // @[Top.scala 50:10]
  assign n2_I_5 = n1_O_5; // @[Top.scala 50:10]
  assign n2_I_6 = n1_O_6; // @[Top.scala 50:10]
  assign n2_I_7 = n1_O_7; // @[Top.scala 50:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 54:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 53:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 53:10]
  assign n3_I_2 = n2_O_2; // @[Top.scala 53:10]
  assign n3_I_3 = n2_O_3; // @[Top.scala 53:10]
  assign n3_I_4 = n2_O_4; // @[Top.scala 53:10]
  assign n3_I_5 = n2_O_5; // @[Top.scala 53:10]
  assign n3_I_6 = n2_O_6; // @[Top.scala 53:10]
  assign n3_I_7 = n2_O_7; // @[Top.scala 53:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 57:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 56:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 56:10]
  assign n4_I_2 = n3_O_2; // @[Top.scala 56:10]
  assign n4_I_3 = n3_O_3; // @[Top.scala 56:10]
  assign n4_I_4 = n3_O_4; // @[Top.scala 56:10]
  assign n4_I_5 = n3_O_5; // @[Top.scala 56:10]
  assign n4_I_6 = n3_O_6; // @[Top.scala 56:10]
  assign n4_I_7 = n3_O_7; // @[Top.scala 56:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 60:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 59:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 59:10]
  assign n5_I_2 = n4_O_2; // @[Top.scala 59:10]
  assign n5_I_3 = n4_O_3; // @[Top.scala 59:10]
  assign n5_I_4 = n4_O_4; // @[Top.scala 59:10]
  assign n5_I_5 = n4_O_5; // @[Top.scala 59:10]
  assign n5_I_6 = n4_O_6; // @[Top.scala 59:10]
  assign n5_I_7 = n4_O_7; // @[Top.scala 59:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 64:17]
  assign n6_I0_0 = n5_O_0; // @[Top.scala 62:11]
  assign n6_I0_1 = n5_O_1; // @[Top.scala 62:11]
  assign n6_I0_2 = n5_O_2; // @[Top.scala 62:11]
  assign n6_I0_3 = n5_O_3; // @[Top.scala 62:11]
  assign n6_I0_4 = n5_O_4; // @[Top.scala 62:11]
  assign n6_I0_5 = n5_O_5; // @[Top.scala 62:11]
  assign n6_I0_6 = n5_O_6; // @[Top.scala 62:11]
  assign n6_I0_7 = n5_O_7; // @[Top.scala 62:11]
  assign n6_I1_0 = n4_O_0; // @[Top.scala 63:11]
  assign n6_I1_1 = n4_O_1; // @[Top.scala 63:11]
  assign n6_I1_2 = n4_O_2; // @[Top.scala 63:11]
  assign n6_I1_3 = n4_O_3; // @[Top.scala 63:11]
  assign n6_I1_4 = n4_O_4; // @[Top.scala 63:11]
  assign n6_I1_5 = n4_O_5; // @[Top.scala 63:11]
  assign n6_I1_6 = n4_O_6; // @[Top.scala 63:11]
  assign n6_I1_7 = n4_O_7; // @[Top.scala 63:11]
  assign n13_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 68:18]
  assign n13_I0_0_0 = n6_O_0_0; // @[Top.scala 66:12]
  assign n13_I0_0_1 = n6_O_0_1; // @[Top.scala 66:12]
  assign n13_I0_1_0 = n6_O_1_0; // @[Top.scala 66:12]
  assign n13_I0_1_1 = n6_O_1_1; // @[Top.scala 66:12]
  assign n13_I0_2_0 = n6_O_2_0; // @[Top.scala 66:12]
  assign n13_I0_2_1 = n6_O_2_1; // @[Top.scala 66:12]
  assign n13_I0_3_0 = n6_O_3_0; // @[Top.scala 66:12]
  assign n13_I0_3_1 = n6_O_3_1; // @[Top.scala 66:12]
  assign n13_I0_4_0 = n6_O_4_0; // @[Top.scala 66:12]
  assign n13_I0_4_1 = n6_O_4_1; // @[Top.scala 66:12]
  assign n13_I0_5_0 = n6_O_5_0; // @[Top.scala 66:12]
  assign n13_I0_5_1 = n6_O_5_1; // @[Top.scala 66:12]
  assign n13_I0_6_0 = n6_O_6_0; // @[Top.scala 66:12]
  assign n13_I0_6_1 = n6_O_6_1; // @[Top.scala 66:12]
  assign n13_I0_7_0 = n6_O_7_0; // @[Top.scala 66:12]
  assign n13_I0_7_1 = n6_O_7_1; // @[Top.scala 66:12]
  assign n13_I1_0 = n3_O_0; // @[Top.scala 67:12]
  assign n13_I1_1 = n3_O_1; // @[Top.scala 67:12]
  assign n13_I1_2 = n3_O_2; // @[Top.scala 67:12]
  assign n13_I1_3 = n3_O_3; // @[Top.scala 67:12]
  assign n13_I1_4 = n3_O_4; // @[Top.scala 67:12]
  assign n13_I1_5 = n3_O_5; // @[Top.scala 67:12]
  assign n13_I1_6 = n3_O_6; // @[Top.scala 67:12]
  assign n13_I1_7 = n3_O_7; // @[Top.scala 67:12]
  assign n22_valid_up = n13_valid_down; // @[Top.scala 71:18]
  assign n22_I_0_0 = n13_O_0_0; // @[Top.scala 70:11]
  assign n22_I_0_1 = n13_O_0_1; // @[Top.scala 70:11]
  assign n22_I_0_2 = n13_O_0_2; // @[Top.scala 70:11]
  assign n22_I_1_0 = n13_O_1_0; // @[Top.scala 70:11]
  assign n22_I_1_1 = n13_O_1_1; // @[Top.scala 70:11]
  assign n22_I_1_2 = n13_O_1_2; // @[Top.scala 70:11]
  assign n22_I_2_0 = n13_O_2_0; // @[Top.scala 70:11]
  assign n22_I_2_1 = n13_O_2_1; // @[Top.scala 70:11]
  assign n22_I_2_2 = n13_O_2_2; // @[Top.scala 70:11]
  assign n22_I_3_0 = n13_O_3_0; // @[Top.scala 70:11]
  assign n22_I_3_1 = n13_O_3_1; // @[Top.scala 70:11]
  assign n22_I_3_2 = n13_O_3_2; // @[Top.scala 70:11]
  assign n22_I_4_0 = n13_O_4_0; // @[Top.scala 70:11]
  assign n22_I_4_1 = n13_O_4_1; // @[Top.scala 70:11]
  assign n22_I_4_2 = n13_O_4_2; // @[Top.scala 70:11]
  assign n22_I_5_0 = n13_O_5_0; // @[Top.scala 70:11]
  assign n22_I_5_1 = n13_O_5_1; // @[Top.scala 70:11]
  assign n22_I_5_2 = n13_O_5_2; // @[Top.scala 70:11]
  assign n22_I_6_0 = n13_O_6_0; // @[Top.scala 70:11]
  assign n22_I_6_1 = n13_O_6_1; // @[Top.scala 70:11]
  assign n22_I_6_2 = n13_O_6_2; // @[Top.scala 70:11]
  assign n22_I_7_0 = n13_O_7_0; // @[Top.scala 70:11]
  assign n22_I_7_1 = n13_O_7_1; // @[Top.scala 70:11]
  assign n22_I_7_2 = n13_O_7_2; // @[Top.scala 70:11]
  assign n29_valid_up = n22_valid_down; // @[Top.scala 74:18]
  assign n29_I_0_0_0 = n22_O_0_0_0; // @[Top.scala 73:11]
  assign n29_I_0_0_1 = n22_O_0_0_1; // @[Top.scala 73:11]
  assign n29_I_0_0_2 = n22_O_0_0_2; // @[Top.scala 73:11]
  assign n29_I_1_0_0 = n22_O_1_0_0; // @[Top.scala 73:11]
  assign n29_I_1_0_1 = n22_O_1_0_1; // @[Top.scala 73:11]
  assign n29_I_1_0_2 = n22_O_1_0_2; // @[Top.scala 73:11]
  assign n29_I_2_0_0 = n22_O_2_0_0; // @[Top.scala 73:11]
  assign n29_I_2_0_1 = n22_O_2_0_1; // @[Top.scala 73:11]
  assign n29_I_2_0_2 = n22_O_2_0_2; // @[Top.scala 73:11]
  assign n29_I_3_0_0 = n22_O_3_0_0; // @[Top.scala 73:11]
  assign n29_I_3_0_1 = n22_O_3_0_1; // @[Top.scala 73:11]
  assign n29_I_3_0_2 = n22_O_3_0_2; // @[Top.scala 73:11]
  assign n29_I_4_0_0 = n22_O_4_0_0; // @[Top.scala 73:11]
  assign n29_I_4_0_1 = n22_O_4_0_1; // @[Top.scala 73:11]
  assign n29_I_4_0_2 = n22_O_4_0_2; // @[Top.scala 73:11]
  assign n29_I_5_0_0 = n22_O_5_0_0; // @[Top.scala 73:11]
  assign n29_I_5_0_1 = n22_O_5_0_1; // @[Top.scala 73:11]
  assign n29_I_5_0_2 = n22_O_5_0_2; // @[Top.scala 73:11]
  assign n29_I_6_0_0 = n22_O_6_0_0; // @[Top.scala 73:11]
  assign n29_I_6_0_1 = n22_O_6_0_1; // @[Top.scala 73:11]
  assign n29_I_6_0_2 = n22_O_6_0_2; // @[Top.scala 73:11]
  assign n29_I_7_0_0 = n22_O_7_0_0; // @[Top.scala 73:11]
  assign n29_I_7_0_1 = n22_O_7_0_1; // @[Top.scala 73:11]
  assign n29_I_7_0_2 = n22_O_7_0_2; // @[Top.scala 73:11]
  assign n30_clock = clock;
  assign n30_valid_up = n2_valid_down; // @[Top.scala 77:18]
  assign n30_I_0 = n2_O_0; // @[Top.scala 76:11]
  assign n30_I_1 = n2_O_1; // @[Top.scala 76:11]
  assign n30_I_2 = n2_O_2; // @[Top.scala 76:11]
  assign n30_I_3 = n2_O_3; // @[Top.scala 76:11]
  assign n30_I_4 = n2_O_4; // @[Top.scala 76:11]
  assign n30_I_5 = n2_O_5; // @[Top.scala 76:11]
  assign n30_I_6 = n2_O_6; // @[Top.scala 76:11]
  assign n30_I_7 = n2_O_7; // @[Top.scala 76:11]
  assign n31_clock = clock;
  assign n31_valid_up = n30_valid_down; // @[Top.scala 80:18]
  assign n31_I_0 = n30_O_0; // @[Top.scala 79:11]
  assign n31_I_1 = n30_O_1; // @[Top.scala 79:11]
  assign n31_I_2 = n30_O_2; // @[Top.scala 79:11]
  assign n31_I_3 = n30_O_3; // @[Top.scala 79:11]
  assign n31_I_4 = n30_O_4; // @[Top.scala 79:11]
  assign n31_I_5 = n30_O_5; // @[Top.scala 79:11]
  assign n31_I_6 = n30_O_6; // @[Top.scala 79:11]
  assign n31_I_7 = n30_O_7; // @[Top.scala 79:11]
  assign n32_valid_up = n31_valid_down & n30_valid_down; // @[Top.scala 84:18]
  assign n32_I0_0 = n31_O_0; // @[Top.scala 82:12]
  assign n32_I0_1 = n31_O_1; // @[Top.scala 82:12]
  assign n32_I0_2 = n31_O_2; // @[Top.scala 82:12]
  assign n32_I0_3 = n31_O_3; // @[Top.scala 82:12]
  assign n32_I0_4 = n31_O_4; // @[Top.scala 82:12]
  assign n32_I0_5 = n31_O_5; // @[Top.scala 82:12]
  assign n32_I0_6 = n31_O_6; // @[Top.scala 82:12]
  assign n32_I0_7 = n31_O_7; // @[Top.scala 82:12]
  assign n32_I1_0 = n30_O_0; // @[Top.scala 83:12]
  assign n32_I1_1 = n30_O_1; // @[Top.scala 83:12]
  assign n32_I1_2 = n30_O_2; // @[Top.scala 83:12]
  assign n32_I1_3 = n30_O_3; // @[Top.scala 83:12]
  assign n32_I1_4 = n30_O_4; // @[Top.scala 83:12]
  assign n32_I1_5 = n30_O_5; // @[Top.scala 83:12]
  assign n32_I1_6 = n30_O_6; // @[Top.scala 83:12]
  assign n32_I1_7 = n30_O_7; // @[Top.scala 83:12]
  assign n39_valid_up = n32_valid_down & n2_valid_down; // @[Top.scala 88:18]
  assign n39_I0_0_0 = n32_O_0_0; // @[Top.scala 86:12]
  assign n39_I0_0_1 = n32_O_0_1; // @[Top.scala 86:12]
  assign n39_I0_1_0 = n32_O_1_0; // @[Top.scala 86:12]
  assign n39_I0_1_1 = n32_O_1_1; // @[Top.scala 86:12]
  assign n39_I0_2_0 = n32_O_2_0; // @[Top.scala 86:12]
  assign n39_I0_2_1 = n32_O_2_1; // @[Top.scala 86:12]
  assign n39_I0_3_0 = n32_O_3_0; // @[Top.scala 86:12]
  assign n39_I0_3_1 = n32_O_3_1; // @[Top.scala 86:12]
  assign n39_I0_4_0 = n32_O_4_0; // @[Top.scala 86:12]
  assign n39_I0_4_1 = n32_O_4_1; // @[Top.scala 86:12]
  assign n39_I0_5_0 = n32_O_5_0; // @[Top.scala 86:12]
  assign n39_I0_5_1 = n32_O_5_1; // @[Top.scala 86:12]
  assign n39_I0_6_0 = n32_O_6_0; // @[Top.scala 86:12]
  assign n39_I0_6_1 = n32_O_6_1; // @[Top.scala 86:12]
  assign n39_I0_7_0 = n32_O_7_0; // @[Top.scala 86:12]
  assign n39_I0_7_1 = n32_O_7_1; // @[Top.scala 86:12]
  assign n39_I1_0 = n2_O_0; // @[Top.scala 87:12]
  assign n39_I1_1 = n2_O_1; // @[Top.scala 87:12]
  assign n39_I1_2 = n2_O_2; // @[Top.scala 87:12]
  assign n39_I1_3 = n2_O_3; // @[Top.scala 87:12]
  assign n39_I1_4 = n2_O_4; // @[Top.scala 87:12]
  assign n39_I1_5 = n2_O_5; // @[Top.scala 87:12]
  assign n39_I1_6 = n2_O_6; // @[Top.scala 87:12]
  assign n39_I1_7 = n2_O_7; // @[Top.scala 87:12]
  assign n48_valid_up = n39_valid_down; // @[Top.scala 91:18]
  assign n48_I_0_0 = n39_O_0_0; // @[Top.scala 90:11]
  assign n48_I_0_1 = n39_O_0_1; // @[Top.scala 90:11]
  assign n48_I_0_2 = n39_O_0_2; // @[Top.scala 90:11]
  assign n48_I_1_0 = n39_O_1_0; // @[Top.scala 90:11]
  assign n48_I_1_1 = n39_O_1_1; // @[Top.scala 90:11]
  assign n48_I_1_2 = n39_O_1_2; // @[Top.scala 90:11]
  assign n48_I_2_0 = n39_O_2_0; // @[Top.scala 90:11]
  assign n48_I_2_1 = n39_O_2_1; // @[Top.scala 90:11]
  assign n48_I_2_2 = n39_O_2_2; // @[Top.scala 90:11]
  assign n48_I_3_0 = n39_O_3_0; // @[Top.scala 90:11]
  assign n48_I_3_1 = n39_O_3_1; // @[Top.scala 90:11]
  assign n48_I_3_2 = n39_O_3_2; // @[Top.scala 90:11]
  assign n48_I_4_0 = n39_O_4_0; // @[Top.scala 90:11]
  assign n48_I_4_1 = n39_O_4_1; // @[Top.scala 90:11]
  assign n48_I_4_2 = n39_O_4_2; // @[Top.scala 90:11]
  assign n48_I_5_0 = n39_O_5_0; // @[Top.scala 90:11]
  assign n48_I_5_1 = n39_O_5_1; // @[Top.scala 90:11]
  assign n48_I_5_2 = n39_O_5_2; // @[Top.scala 90:11]
  assign n48_I_6_0 = n39_O_6_0; // @[Top.scala 90:11]
  assign n48_I_6_1 = n39_O_6_1; // @[Top.scala 90:11]
  assign n48_I_6_2 = n39_O_6_2; // @[Top.scala 90:11]
  assign n48_I_7_0 = n39_O_7_0; // @[Top.scala 90:11]
  assign n48_I_7_1 = n39_O_7_1; // @[Top.scala 90:11]
  assign n48_I_7_2 = n39_O_7_2; // @[Top.scala 90:11]
  assign n55_valid_up = n48_valid_down; // @[Top.scala 94:18]
  assign n55_I_0_0_0 = n48_O_0_0_0; // @[Top.scala 93:11]
  assign n55_I_0_0_1 = n48_O_0_0_1; // @[Top.scala 93:11]
  assign n55_I_0_0_2 = n48_O_0_0_2; // @[Top.scala 93:11]
  assign n55_I_1_0_0 = n48_O_1_0_0; // @[Top.scala 93:11]
  assign n55_I_1_0_1 = n48_O_1_0_1; // @[Top.scala 93:11]
  assign n55_I_1_0_2 = n48_O_1_0_2; // @[Top.scala 93:11]
  assign n55_I_2_0_0 = n48_O_2_0_0; // @[Top.scala 93:11]
  assign n55_I_2_0_1 = n48_O_2_0_1; // @[Top.scala 93:11]
  assign n55_I_2_0_2 = n48_O_2_0_2; // @[Top.scala 93:11]
  assign n55_I_3_0_0 = n48_O_3_0_0; // @[Top.scala 93:11]
  assign n55_I_3_0_1 = n48_O_3_0_1; // @[Top.scala 93:11]
  assign n55_I_3_0_2 = n48_O_3_0_2; // @[Top.scala 93:11]
  assign n55_I_4_0_0 = n48_O_4_0_0; // @[Top.scala 93:11]
  assign n55_I_4_0_1 = n48_O_4_0_1; // @[Top.scala 93:11]
  assign n55_I_4_0_2 = n48_O_4_0_2; // @[Top.scala 93:11]
  assign n55_I_5_0_0 = n48_O_5_0_0; // @[Top.scala 93:11]
  assign n55_I_5_0_1 = n48_O_5_0_1; // @[Top.scala 93:11]
  assign n55_I_5_0_2 = n48_O_5_0_2; // @[Top.scala 93:11]
  assign n55_I_6_0_0 = n48_O_6_0_0; // @[Top.scala 93:11]
  assign n55_I_6_0_1 = n48_O_6_0_1; // @[Top.scala 93:11]
  assign n55_I_6_0_2 = n48_O_6_0_2; // @[Top.scala 93:11]
  assign n55_I_7_0_0 = n48_O_7_0_0; // @[Top.scala 93:11]
  assign n55_I_7_0_1 = n48_O_7_0_1; // @[Top.scala 93:11]
  assign n55_I_7_0_2 = n48_O_7_0_2; // @[Top.scala 93:11]
  assign n56_valid_up = n29_valid_down & n55_valid_down; // @[Top.scala 98:18]
  assign n56_I0_0_0 = n29_O_0_0; // @[Top.scala 96:12]
  assign n56_I0_0_1 = n29_O_0_1; // @[Top.scala 96:12]
  assign n56_I0_0_2 = n29_O_0_2; // @[Top.scala 96:12]
  assign n56_I0_1_0 = n29_O_1_0; // @[Top.scala 96:12]
  assign n56_I0_1_1 = n29_O_1_1; // @[Top.scala 96:12]
  assign n56_I0_1_2 = n29_O_1_2; // @[Top.scala 96:12]
  assign n56_I0_2_0 = n29_O_2_0; // @[Top.scala 96:12]
  assign n56_I0_2_1 = n29_O_2_1; // @[Top.scala 96:12]
  assign n56_I0_2_2 = n29_O_2_2; // @[Top.scala 96:12]
  assign n56_I0_3_0 = n29_O_3_0; // @[Top.scala 96:12]
  assign n56_I0_3_1 = n29_O_3_1; // @[Top.scala 96:12]
  assign n56_I0_3_2 = n29_O_3_2; // @[Top.scala 96:12]
  assign n56_I0_4_0 = n29_O_4_0; // @[Top.scala 96:12]
  assign n56_I0_4_1 = n29_O_4_1; // @[Top.scala 96:12]
  assign n56_I0_4_2 = n29_O_4_2; // @[Top.scala 96:12]
  assign n56_I0_5_0 = n29_O_5_0; // @[Top.scala 96:12]
  assign n56_I0_5_1 = n29_O_5_1; // @[Top.scala 96:12]
  assign n56_I0_5_2 = n29_O_5_2; // @[Top.scala 96:12]
  assign n56_I0_6_0 = n29_O_6_0; // @[Top.scala 96:12]
  assign n56_I0_6_1 = n29_O_6_1; // @[Top.scala 96:12]
  assign n56_I0_6_2 = n29_O_6_2; // @[Top.scala 96:12]
  assign n56_I0_7_0 = n29_O_7_0; // @[Top.scala 96:12]
  assign n56_I0_7_1 = n29_O_7_1; // @[Top.scala 96:12]
  assign n56_I0_7_2 = n29_O_7_2; // @[Top.scala 96:12]
  assign n56_I1_0_0 = n55_O_0_0; // @[Top.scala 97:12]
  assign n56_I1_0_1 = n55_O_0_1; // @[Top.scala 97:12]
  assign n56_I1_0_2 = n55_O_0_2; // @[Top.scala 97:12]
  assign n56_I1_1_0 = n55_O_1_0; // @[Top.scala 97:12]
  assign n56_I1_1_1 = n55_O_1_1; // @[Top.scala 97:12]
  assign n56_I1_1_2 = n55_O_1_2; // @[Top.scala 97:12]
  assign n56_I1_2_0 = n55_O_2_0; // @[Top.scala 97:12]
  assign n56_I1_2_1 = n55_O_2_1; // @[Top.scala 97:12]
  assign n56_I1_2_2 = n55_O_2_2; // @[Top.scala 97:12]
  assign n56_I1_3_0 = n55_O_3_0; // @[Top.scala 97:12]
  assign n56_I1_3_1 = n55_O_3_1; // @[Top.scala 97:12]
  assign n56_I1_3_2 = n55_O_3_2; // @[Top.scala 97:12]
  assign n56_I1_4_0 = n55_O_4_0; // @[Top.scala 97:12]
  assign n56_I1_4_1 = n55_O_4_1; // @[Top.scala 97:12]
  assign n56_I1_4_2 = n55_O_4_2; // @[Top.scala 97:12]
  assign n56_I1_5_0 = n55_O_5_0; // @[Top.scala 97:12]
  assign n56_I1_5_1 = n55_O_5_1; // @[Top.scala 97:12]
  assign n56_I1_5_2 = n55_O_5_2; // @[Top.scala 97:12]
  assign n56_I1_6_0 = n55_O_6_0; // @[Top.scala 97:12]
  assign n56_I1_6_1 = n55_O_6_1; // @[Top.scala 97:12]
  assign n56_I1_6_2 = n55_O_6_2; // @[Top.scala 97:12]
  assign n56_I1_7_0 = n55_O_7_0; // @[Top.scala 97:12]
  assign n56_I1_7_1 = n55_O_7_1; // @[Top.scala 97:12]
  assign n56_I1_7_2 = n55_O_7_2; // @[Top.scala 97:12]
  assign n63_clock = clock;
  assign n63_valid_up = n1_valid_down; // @[Top.scala 101:18]
  assign n63_I_0 = n1_O_0; // @[Top.scala 100:11]
  assign n63_I_1 = n1_O_1; // @[Top.scala 100:11]
  assign n63_I_2 = n1_O_2; // @[Top.scala 100:11]
  assign n63_I_3 = n1_O_3; // @[Top.scala 100:11]
  assign n63_I_4 = n1_O_4; // @[Top.scala 100:11]
  assign n63_I_5 = n1_O_5; // @[Top.scala 100:11]
  assign n63_I_6 = n1_O_6; // @[Top.scala 100:11]
  assign n63_I_7 = n1_O_7; // @[Top.scala 100:11]
  assign n64_clock = clock;
  assign n64_valid_up = n63_valid_down; // @[Top.scala 104:18]
  assign n64_I_0 = n63_O_0; // @[Top.scala 103:11]
  assign n64_I_1 = n63_O_1; // @[Top.scala 103:11]
  assign n64_I_2 = n63_O_2; // @[Top.scala 103:11]
  assign n64_I_3 = n63_O_3; // @[Top.scala 103:11]
  assign n64_I_4 = n63_O_4; // @[Top.scala 103:11]
  assign n64_I_5 = n63_O_5; // @[Top.scala 103:11]
  assign n64_I_6 = n63_O_6; // @[Top.scala 103:11]
  assign n64_I_7 = n63_O_7; // @[Top.scala 103:11]
  assign n65_valid_up = n64_valid_down & n63_valid_down; // @[Top.scala 108:18]
  assign n65_I0_0 = n64_O_0; // @[Top.scala 106:12]
  assign n65_I0_1 = n64_O_1; // @[Top.scala 106:12]
  assign n65_I0_2 = n64_O_2; // @[Top.scala 106:12]
  assign n65_I0_3 = n64_O_3; // @[Top.scala 106:12]
  assign n65_I0_4 = n64_O_4; // @[Top.scala 106:12]
  assign n65_I0_5 = n64_O_5; // @[Top.scala 106:12]
  assign n65_I0_6 = n64_O_6; // @[Top.scala 106:12]
  assign n65_I0_7 = n64_O_7; // @[Top.scala 106:12]
  assign n65_I1_0 = n63_O_0; // @[Top.scala 107:12]
  assign n65_I1_1 = n63_O_1; // @[Top.scala 107:12]
  assign n65_I1_2 = n63_O_2; // @[Top.scala 107:12]
  assign n65_I1_3 = n63_O_3; // @[Top.scala 107:12]
  assign n65_I1_4 = n63_O_4; // @[Top.scala 107:12]
  assign n65_I1_5 = n63_O_5; // @[Top.scala 107:12]
  assign n65_I1_6 = n63_O_6; // @[Top.scala 107:12]
  assign n65_I1_7 = n63_O_7; // @[Top.scala 107:12]
  assign n72_valid_up = n65_valid_down & n1_valid_down; // @[Top.scala 112:18]
  assign n72_I0_0_0 = n65_O_0_0; // @[Top.scala 110:12]
  assign n72_I0_0_1 = n65_O_0_1; // @[Top.scala 110:12]
  assign n72_I0_1_0 = n65_O_1_0; // @[Top.scala 110:12]
  assign n72_I0_1_1 = n65_O_1_1; // @[Top.scala 110:12]
  assign n72_I0_2_0 = n65_O_2_0; // @[Top.scala 110:12]
  assign n72_I0_2_1 = n65_O_2_1; // @[Top.scala 110:12]
  assign n72_I0_3_0 = n65_O_3_0; // @[Top.scala 110:12]
  assign n72_I0_3_1 = n65_O_3_1; // @[Top.scala 110:12]
  assign n72_I0_4_0 = n65_O_4_0; // @[Top.scala 110:12]
  assign n72_I0_4_1 = n65_O_4_1; // @[Top.scala 110:12]
  assign n72_I0_5_0 = n65_O_5_0; // @[Top.scala 110:12]
  assign n72_I0_5_1 = n65_O_5_1; // @[Top.scala 110:12]
  assign n72_I0_6_0 = n65_O_6_0; // @[Top.scala 110:12]
  assign n72_I0_6_1 = n65_O_6_1; // @[Top.scala 110:12]
  assign n72_I0_7_0 = n65_O_7_0; // @[Top.scala 110:12]
  assign n72_I0_7_1 = n65_O_7_1; // @[Top.scala 110:12]
  assign n72_I1_0 = n1_O_0; // @[Top.scala 111:12]
  assign n72_I1_1 = n1_O_1; // @[Top.scala 111:12]
  assign n72_I1_2 = n1_O_2; // @[Top.scala 111:12]
  assign n72_I1_3 = n1_O_3; // @[Top.scala 111:12]
  assign n72_I1_4 = n1_O_4; // @[Top.scala 111:12]
  assign n72_I1_5 = n1_O_5; // @[Top.scala 111:12]
  assign n72_I1_6 = n1_O_6; // @[Top.scala 111:12]
  assign n72_I1_7 = n1_O_7; // @[Top.scala 111:12]
  assign n81_valid_up = n72_valid_down; // @[Top.scala 115:18]
  assign n81_I_0_0 = n72_O_0_0; // @[Top.scala 114:11]
  assign n81_I_0_1 = n72_O_0_1; // @[Top.scala 114:11]
  assign n81_I_0_2 = n72_O_0_2; // @[Top.scala 114:11]
  assign n81_I_1_0 = n72_O_1_0; // @[Top.scala 114:11]
  assign n81_I_1_1 = n72_O_1_1; // @[Top.scala 114:11]
  assign n81_I_1_2 = n72_O_1_2; // @[Top.scala 114:11]
  assign n81_I_2_0 = n72_O_2_0; // @[Top.scala 114:11]
  assign n81_I_2_1 = n72_O_2_1; // @[Top.scala 114:11]
  assign n81_I_2_2 = n72_O_2_2; // @[Top.scala 114:11]
  assign n81_I_3_0 = n72_O_3_0; // @[Top.scala 114:11]
  assign n81_I_3_1 = n72_O_3_1; // @[Top.scala 114:11]
  assign n81_I_3_2 = n72_O_3_2; // @[Top.scala 114:11]
  assign n81_I_4_0 = n72_O_4_0; // @[Top.scala 114:11]
  assign n81_I_4_1 = n72_O_4_1; // @[Top.scala 114:11]
  assign n81_I_4_2 = n72_O_4_2; // @[Top.scala 114:11]
  assign n81_I_5_0 = n72_O_5_0; // @[Top.scala 114:11]
  assign n81_I_5_1 = n72_O_5_1; // @[Top.scala 114:11]
  assign n81_I_5_2 = n72_O_5_2; // @[Top.scala 114:11]
  assign n81_I_6_0 = n72_O_6_0; // @[Top.scala 114:11]
  assign n81_I_6_1 = n72_O_6_1; // @[Top.scala 114:11]
  assign n81_I_6_2 = n72_O_6_2; // @[Top.scala 114:11]
  assign n81_I_7_0 = n72_O_7_0; // @[Top.scala 114:11]
  assign n81_I_7_1 = n72_O_7_1; // @[Top.scala 114:11]
  assign n81_I_7_2 = n72_O_7_2; // @[Top.scala 114:11]
  assign n88_valid_up = n81_valid_down; // @[Top.scala 118:18]
  assign n88_I_0_0_0 = n81_O_0_0_0; // @[Top.scala 117:11]
  assign n88_I_0_0_1 = n81_O_0_0_1; // @[Top.scala 117:11]
  assign n88_I_0_0_2 = n81_O_0_0_2; // @[Top.scala 117:11]
  assign n88_I_1_0_0 = n81_O_1_0_0; // @[Top.scala 117:11]
  assign n88_I_1_0_1 = n81_O_1_0_1; // @[Top.scala 117:11]
  assign n88_I_1_0_2 = n81_O_1_0_2; // @[Top.scala 117:11]
  assign n88_I_2_0_0 = n81_O_2_0_0; // @[Top.scala 117:11]
  assign n88_I_2_0_1 = n81_O_2_0_1; // @[Top.scala 117:11]
  assign n88_I_2_0_2 = n81_O_2_0_2; // @[Top.scala 117:11]
  assign n88_I_3_0_0 = n81_O_3_0_0; // @[Top.scala 117:11]
  assign n88_I_3_0_1 = n81_O_3_0_1; // @[Top.scala 117:11]
  assign n88_I_3_0_2 = n81_O_3_0_2; // @[Top.scala 117:11]
  assign n88_I_4_0_0 = n81_O_4_0_0; // @[Top.scala 117:11]
  assign n88_I_4_0_1 = n81_O_4_0_1; // @[Top.scala 117:11]
  assign n88_I_4_0_2 = n81_O_4_0_2; // @[Top.scala 117:11]
  assign n88_I_5_0_0 = n81_O_5_0_0; // @[Top.scala 117:11]
  assign n88_I_5_0_1 = n81_O_5_0_1; // @[Top.scala 117:11]
  assign n88_I_5_0_2 = n81_O_5_0_2; // @[Top.scala 117:11]
  assign n88_I_6_0_0 = n81_O_6_0_0; // @[Top.scala 117:11]
  assign n88_I_6_0_1 = n81_O_6_0_1; // @[Top.scala 117:11]
  assign n88_I_6_0_2 = n81_O_6_0_2; // @[Top.scala 117:11]
  assign n88_I_7_0_0 = n81_O_7_0_0; // @[Top.scala 117:11]
  assign n88_I_7_0_1 = n81_O_7_0_1; // @[Top.scala 117:11]
  assign n88_I_7_0_2 = n81_O_7_0_2; // @[Top.scala 117:11]
  assign n89_valid_up = n56_valid_down & n88_valid_down; // @[Top.scala 122:18]
  assign n89_I0_0_0_0 = n56_O_0_0_0; // @[Top.scala 120:12]
  assign n89_I0_0_0_1 = n56_O_0_0_1; // @[Top.scala 120:12]
  assign n89_I0_0_0_2 = n56_O_0_0_2; // @[Top.scala 120:12]
  assign n89_I0_0_1_0 = n56_O_0_1_0; // @[Top.scala 120:12]
  assign n89_I0_0_1_1 = n56_O_0_1_1; // @[Top.scala 120:12]
  assign n89_I0_0_1_2 = n56_O_0_1_2; // @[Top.scala 120:12]
  assign n89_I0_1_0_0 = n56_O_1_0_0; // @[Top.scala 120:12]
  assign n89_I0_1_0_1 = n56_O_1_0_1; // @[Top.scala 120:12]
  assign n89_I0_1_0_2 = n56_O_1_0_2; // @[Top.scala 120:12]
  assign n89_I0_1_1_0 = n56_O_1_1_0; // @[Top.scala 120:12]
  assign n89_I0_1_1_1 = n56_O_1_1_1; // @[Top.scala 120:12]
  assign n89_I0_1_1_2 = n56_O_1_1_2; // @[Top.scala 120:12]
  assign n89_I0_2_0_0 = n56_O_2_0_0; // @[Top.scala 120:12]
  assign n89_I0_2_0_1 = n56_O_2_0_1; // @[Top.scala 120:12]
  assign n89_I0_2_0_2 = n56_O_2_0_2; // @[Top.scala 120:12]
  assign n89_I0_2_1_0 = n56_O_2_1_0; // @[Top.scala 120:12]
  assign n89_I0_2_1_1 = n56_O_2_1_1; // @[Top.scala 120:12]
  assign n89_I0_2_1_2 = n56_O_2_1_2; // @[Top.scala 120:12]
  assign n89_I0_3_0_0 = n56_O_3_0_0; // @[Top.scala 120:12]
  assign n89_I0_3_0_1 = n56_O_3_0_1; // @[Top.scala 120:12]
  assign n89_I0_3_0_2 = n56_O_3_0_2; // @[Top.scala 120:12]
  assign n89_I0_3_1_0 = n56_O_3_1_0; // @[Top.scala 120:12]
  assign n89_I0_3_1_1 = n56_O_3_1_1; // @[Top.scala 120:12]
  assign n89_I0_3_1_2 = n56_O_3_1_2; // @[Top.scala 120:12]
  assign n89_I0_4_0_0 = n56_O_4_0_0; // @[Top.scala 120:12]
  assign n89_I0_4_0_1 = n56_O_4_0_1; // @[Top.scala 120:12]
  assign n89_I0_4_0_2 = n56_O_4_0_2; // @[Top.scala 120:12]
  assign n89_I0_4_1_0 = n56_O_4_1_0; // @[Top.scala 120:12]
  assign n89_I0_4_1_1 = n56_O_4_1_1; // @[Top.scala 120:12]
  assign n89_I0_4_1_2 = n56_O_4_1_2; // @[Top.scala 120:12]
  assign n89_I0_5_0_0 = n56_O_5_0_0; // @[Top.scala 120:12]
  assign n89_I0_5_0_1 = n56_O_5_0_1; // @[Top.scala 120:12]
  assign n89_I0_5_0_2 = n56_O_5_0_2; // @[Top.scala 120:12]
  assign n89_I0_5_1_0 = n56_O_5_1_0; // @[Top.scala 120:12]
  assign n89_I0_5_1_1 = n56_O_5_1_1; // @[Top.scala 120:12]
  assign n89_I0_5_1_2 = n56_O_5_1_2; // @[Top.scala 120:12]
  assign n89_I0_6_0_0 = n56_O_6_0_0; // @[Top.scala 120:12]
  assign n89_I0_6_0_1 = n56_O_6_0_1; // @[Top.scala 120:12]
  assign n89_I0_6_0_2 = n56_O_6_0_2; // @[Top.scala 120:12]
  assign n89_I0_6_1_0 = n56_O_6_1_0; // @[Top.scala 120:12]
  assign n89_I0_6_1_1 = n56_O_6_1_1; // @[Top.scala 120:12]
  assign n89_I0_6_1_2 = n56_O_6_1_2; // @[Top.scala 120:12]
  assign n89_I0_7_0_0 = n56_O_7_0_0; // @[Top.scala 120:12]
  assign n89_I0_7_0_1 = n56_O_7_0_1; // @[Top.scala 120:12]
  assign n89_I0_7_0_2 = n56_O_7_0_2; // @[Top.scala 120:12]
  assign n89_I0_7_1_0 = n56_O_7_1_0; // @[Top.scala 120:12]
  assign n89_I0_7_1_1 = n56_O_7_1_1; // @[Top.scala 120:12]
  assign n89_I0_7_1_2 = n56_O_7_1_2; // @[Top.scala 120:12]
  assign n89_I1_0_0 = n88_O_0_0; // @[Top.scala 121:12]
  assign n89_I1_0_1 = n88_O_0_1; // @[Top.scala 121:12]
  assign n89_I1_0_2 = n88_O_0_2; // @[Top.scala 121:12]
  assign n89_I1_1_0 = n88_O_1_0; // @[Top.scala 121:12]
  assign n89_I1_1_1 = n88_O_1_1; // @[Top.scala 121:12]
  assign n89_I1_1_2 = n88_O_1_2; // @[Top.scala 121:12]
  assign n89_I1_2_0 = n88_O_2_0; // @[Top.scala 121:12]
  assign n89_I1_2_1 = n88_O_2_1; // @[Top.scala 121:12]
  assign n89_I1_2_2 = n88_O_2_2; // @[Top.scala 121:12]
  assign n89_I1_3_0 = n88_O_3_0; // @[Top.scala 121:12]
  assign n89_I1_3_1 = n88_O_3_1; // @[Top.scala 121:12]
  assign n89_I1_3_2 = n88_O_3_2; // @[Top.scala 121:12]
  assign n89_I1_4_0 = n88_O_4_0; // @[Top.scala 121:12]
  assign n89_I1_4_1 = n88_O_4_1; // @[Top.scala 121:12]
  assign n89_I1_4_2 = n88_O_4_2; // @[Top.scala 121:12]
  assign n89_I1_5_0 = n88_O_5_0; // @[Top.scala 121:12]
  assign n89_I1_5_1 = n88_O_5_1; // @[Top.scala 121:12]
  assign n89_I1_5_2 = n88_O_5_2; // @[Top.scala 121:12]
  assign n89_I1_6_0 = n88_O_6_0; // @[Top.scala 121:12]
  assign n89_I1_6_1 = n88_O_6_1; // @[Top.scala 121:12]
  assign n89_I1_6_2 = n88_O_6_2; // @[Top.scala 121:12]
  assign n89_I1_7_0 = n88_O_7_0; // @[Top.scala 121:12]
  assign n89_I1_7_1 = n88_O_7_1; // @[Top.scala 121:12]
  assign n89_I1_7_2 = n88_O_7_2; // @[Top.scala 121:12]
  assign n98_valid_up = n89_valid_down; // @[Top.scala 125:18]
  assign n98_I_0_0_0 = n89_O_0_0_0; // @[Top.scala 124:11]
  assign n98_I_0_0_1 = n89_O_0_0_1; // @[Top.scala 124:11]
  assign n98_I_0_0_2 = n89_O_0_0_2; // @[Top.scala 124:11]
  assign n98_I_0_1_0 = n89_O_0_1_0; // @[Top.scala 124:11]
  assign n98_I_0_1_1 = n89_O_0_1_1; // @[Top.scala 124:11]
  assign n98_I_0_1_2 = n89_O_0_1_2; // @[Top.scala 124:11]
  assign n98_I_0_2_0 = n89_O_0_2_0; // @[Top.scala 124:11]
  assign n98_I_0_2_1 = n89_O_0_2_1; // @[Top.scala 124:11]
  assign n98_I_0_2_2 = n89_O_0_2_2; // @[Top.scala 124:11]
  assign n98_I_1_0_0 = n89_O_1_0_0; // @[Top.scala 124:11]
  assign n98_I_1_0_1 = n89_O_1_0_1; // @[Top.scala 124:11]
  assign n98_I_1_0_2 = n89_O_1_0_2; // @[Top.scala 124:11]
  assign n98_I_1_1_0 = n89_O_1_1_0; // @[Top.scala 124:11]
  assign n98_I_1_1_1 = n89_O_1_1_1; // @[Top.scala 124:11]
  assign n98_I_1_1_2 = n89_O_1_1_2; // @[Top.scala 124:11]
  assign n98_I_1_2_0 = n89_O_1_2_0; // @[Top.scala 124:11]
  assign n98_I_1_2_1 = n89_O_1_2_1; // @[Top.scala 124:11]
  assign n98_I_1_2_2 = n89_O_1_2_2; // @[Top.scala 124:11]
  assign n98_I_2_0_0 = n89_O_2_0_0; // @[Top.scala 124:11]
  assign n98_I_2_0_1 = n89_O_2_0_1; // @[Top.scala 124:11]
  assign n98_I_2_0_2 = n89_O_2_0_2; // @[Top.scala 124:11]
  assign n98_I_2_1_0 = n89_O_2_1_0; // @[Top.scala 124:11]
  assign n98_I_2_1_1 = n89_O_2_1_1; // @[Top.scala 124:11]
  assign n98_I_2_1_2 = n89_O_2_1_2; // @[Top.scala 124:11]
  assign n98_I_2_2_0 = n89_O_2_2_0; // @[Top.scala 124:11]
  assign n98_I_2_2_1 = n89_O_2_2_1; // @[Top.scala 124:11]
  assign n98_I_2_2_2 = n89_O_2_2_2; // @[Top.scala 124:11]
  assign n98_I_3_0_0 = n89_O_3_0_0; // @[Top.scala 124:11]
  assign n98_I_3_0_1 = n89_O_3_0_1; // @[Top.scala 124:11]
  assign n98_I_3_0_2 = n89_O_3_0_2; // @[Top.scala 124:11]
  assign n98_I_3_1_0 = n89_O_3_1_0; // @[Top.scala 124:11]
  assign n98_I_3_1_1 = n89_O_3_1_1; // @[Top.scala 124:11]
  assign n98_I_3_1_2 = n89_O_3_1_2; // @[Top.scala 124:11]
  assign n98_I_3_2_0 = n89_O_3_2_0; // @[Top.scala 124:11]
  assign n98_I_3_2_1 = n89_O_3_2_1; // @[Top.scala 124:11]
  assign n98_I_3_2_2 = n89_O_3_2_2; // @[Top.scala 124:11]
  assign n98_I_4_0_0 = n89_O_4_0_0; // @[Top.scala 124:11]
  assign n98_I_4_0_1 = n89_O_4_0_1; // @[Top.scala 124:11]
  assign n98_I_4_0_2 = n89_O_4_0_2; // @[Top.scala 124:11]
  assign n98_I_4_1_0 = n89_O_4_1_0; // @[Top.scala 124:11]
  assign n98_I_4_1_1 = n89_O_4_1_1; // @[Top.scala 124:11]
  assign n98_I_4_1_2 = n89_O_4_1_2; // @[Top.scala 124:11]
  assign n98_I_4_2_0 = n89_O_4_2_0; // @[Top.scala 124:11]
  assign n98_I_4_2_1 = n89_O_4_2_1; // @[Top.scala 124:11]
  assign n98_I_4_2_2 = n89_O_4_2_2; // @[Top.scala 124:11]
  assign n98_I_5_0_0 = n89_O_5_0_0; // @[Top.scala 124:11]
  assign n98_I_5_0_1 = n89_O_5_0_1; // @[Top.scala 124:11]
  assign n98_I_5_0_2 = n89_O_5_0_2; // @[Top.scala 124:11]
  assign n98_I_5_1_0 = n89_O_5_1_0; // @[Top.scala 124:11]
  assign n98_I_5_1_1 = n89_O_5_1_1; // @[Top.scala 124:11]
  assign n98_I_5_1_2 = n89_O_5_1_2; // @[Top.scala 124:11]
  assign n98_I_5_2_0 = n89_O_5_2_0; // @[Top.scala 124:11]
  assign n98_I_5_2_1 = n89_O_5_2_1; // @[Top.scala 124:11]
  assign n98_I_5_2_2 = n89_O_5_2_2; // @[Top.scala 124:11]
  assign n98_I_6_0_0 = n89_O_6_0_0; // @[Top.scala 124:11]
  assign n98_I_6_0_1 = n89_O_6_0_1; // @[Top.scala 124:11]
  assign n98_I_6_0_2 = n89_O_6_0_2; // @[Top.scala 124:11]
  assign n98_I_6_1_0 = n89_O_6_1_0; // @[Top.scala 124:11]
  assign n98_I_6_1_1 = n89_O_6_1_1; // @[Top.scala 124:11]
  assign n98_I_6_1_2 = n89_O_6_1_2; // @[Top.scala 124:11]
  assign n98_I_6_2_0 = n89_O_6_2_0; // @[Top.scala 124:11]
  assign n98_I_6_2_1 = n89_O_6_2_1; // @[Top.scala 124:11]
  assign n98_I_6_2_2 = n89_O_6_2_2; // @[Top.scala 124:11]
  assign n98_I_7_0_0 = n89_O_7_0_0; // @[Top.scala 124:11]
  assign n98_I_7_0_1 = n89_O_7_0_1; // @[Top.scala 124:11]
  assign n98_I_7_0_2 = n89_O_7_0_2; // @[Top.scala 124:11]
  assign n98_I_7_1_0 = n89_O_7_1_0; // @[Top.scala 124:11]
  assign n98_I_7_1_1 = n89_O_7_1_1; // @[Top.scala 124:11]
  assign n98_I_7_1_2 = n89_O_7_1_2; // @[Top.scala 124:11]
  assign n98_I_7_2_0 = n89_O_7_2_0; // @[Top.scala 124:11]
  assign n98_I_7_2_1 = n89_O_7_2_1; // @[Top.scala 124:11]
  assign n98_I_7_2_2 = n89_O_7_2_2; // @[Top.scala 124:11]
  assign n105_valid_up = n98_valid_down; // @[Top.scala 128:19]
  assign n105_I_0_0_0_0 = n98_O_0_0_0_0; // @[Top.scala 127:12]
  assign n105_I_0_0_0_1 = n98_O_0_0_0_1; // @[Top.scala 127:12]
  assign n105_I_0_0_0_2 = n98_O_0_0_0_2; // @[Top.scala 127:12]
  assign n105_I_0_0_1_0 = n98_O_0_0_1_0; // @[Top.scala 127:12]
  assign n105_I_0_0_1_1 = n98_O_0_0_1_1; // @[Top.scala 127:12]
  assign n105_I_0_0_1_2 = n98_O_0_0_1_2; // @[Top.scala 127:12]
  assign n105_I_0_0_2_0 = n98_O_0_0_2_0; // @[Top.scala 127:12]
  assign n105_I_0_0_2_1 = n98_O_0_0_2_1; // @[Top.scala 127:12]
  assign n105_I_0_0_2_2 = n98_O_0_0_2_2; // @[Top.scala 127:12]
  assign n105_I_1_0_0_0 = n98_O_1_0_0_0; // @[Top.scala 127:12]
  assign n105_I_1_0_0_1 = n98_O_1_0_0_1; // @[Top.scala 127:12]
  assign n105_I_1_0_0_2 = n98_O_1_0_0_2; // @[Top.scala 127:12]
  assign n105_I_1_0_1_0 = n98_O_1_0_1_0; // @[Top.scala 127:12]
  assign n105_I_1_0_1_1 = n98_O_1_0_1_1; // @[Top.scala 127:12]
  assign n105_I_1_0_1_2 = n98_O_1_0_1_2; // @[Top.scala 127:12]
  assign n105_I_1_0_2_0 = n98_O_1_0_2_0; // @[Top.scala 127:12]
  assign n105_I_1_0_2_1 = n98_O_1_0_2_1; // @[Top.scala 127:12]
  assign n105_I_1_0_2_2 = n98_O_1_0_2_2; // @[Top.scala 127:12]
  assign n105_I_2_0_0_0 = n98_O_2_0_0_0; // @[Top.scala 127:12]
  assign n105_I_2_0_0_1 = n98_O_2_0_0_1; // @[Top.scala 127:12]
  assign n105_I_2_0_0_2 = n98_O_2_0_0_2; // @[Top.scala 127:12]
  assign n105_I_2_0_1_0 = n98_O_2_0_1_0; // @[Top.scala 127:12]
  assign n105_I_2_0_1_1 = n98_O_2_0_1_1; // @[Top.scala 127:12]
  assign n105_I_2_0_1_2 = n98_O_2_0_1_2; // @[Top.scala 127:12]
  assign n105_I_2_0_2_0 = n98_O_2_0_2_0; // @[Top.scala 127:12]
  assign n105_I_2_0_2_1 = n98_O_2_0_2_1; // @[Top.scala 127:12]
  assign n105_I_2_0_2_2 = n98_O_2_0_2_2; // @[Top.scala 127:12]
  assign n105_I_3_0_0_0 = n98_O_3_0_0_0; // @[Top.scala 127:12]
  assign n105_I_3_0_0_1 = n98_O_3_0_0_1; // @[Top.scala 127:12]
  assign n105_I_3_0_0_2 = n98_O_3_0_0_2; // @[Top.scala 127:12]
  assign n105_I_3_0_1_0 = n98_O_3_0_1_0; // @[Top.scala 127:12]
  assign n105_I_3_0_1_1 = n98_O_3_0_1_1; // @[Top.scala 127:12]
  assign n105_I_3_0_1_2 = n98_O_3_0_1_2; // @[Top.scala 127:12]
  assign n105_I_3_0_2_0 = n98_O_3_0_2_0; // @[Top.scala 127:12]
  assign n105_I_3_0_2_1 = n98_O_3_0_2_1; // @[Top.scala 127:12]
  assign n105_I_3_0_2_2 = n98_O_3_0_2_2; // @[Top.scala 127:12]
  assign n105_I_4_0_0_0 = n98_O_4_0_0_0; // @[Top.scala 127:12]
  assign n105_I_4_0_0_1 = n98_O_4_0_0_1; // @[Top.scala 127:12]
  assign n105_I_4_0_0_2 = n98_O_4_0_0_2; // @[Top.scala 127:12]
  assign n105_I_4_0_1_0 = n98_O_4_0_1_0; // @[Top.scala 127:12]
  assign n105_I_4_0_1_1 = n98_O_4_0_1_1; // @[Top.scala 127:12]
  assign n105_I_4_0_1_2 = n98_O_4_0_1_2; // @[Top.scala 127:12]
  assign n105_I_4_0_2_0 = n98_O_4_0_2_0; // @[Top.scala 127:12]
  assign n105_I_4_0_2_1 = n98_O_4_0_2_1; // @[Top.scala 127:12]
  assign n105_I_4_0_2_2 = n98_O_4_0_2_2; // @[Top.scala 127:12]
  assign n105_I_5_0_0_0 = n98_O_5_0_0_0; // @[Top.scala 127:12]
  assign n105_I_5_0_0_1 = n98_O_5_0_0_1; // @[Top.scala 127:12]
  assign n105_I_5_0_0_2 = n98_O_5_0_0_2; // @[Top.scala 127:12]
  assign n105_I_5_0_1_0 = n98_O_5_0_1_0; // @[Top.scala 127:12]
  assign n105_I_5_0_1_1 = n98_O_5_0_1_1; // @[Top.scala 127:12]
  assign n105_I_5_0_1_2 = n98_O_5_0_1_2; // @[Top.scala 127:12]
  assign n105_I_5_0_2_0 = n98_O_5_0_2_0; // @[Top.scala 127:12]
  assign n105_I_5_0_2_1 = n98_O_5_0_2_1; // @[Top.scala 127:12]
  assign n105_I_5_0_2_2 = n98_O_5_0_2_2; // @[Top.scala 127:12]
  assign n105_I_6_0_0_0 = n98_O_6_0_0_0; // @[Top.scala 127:12]
  assign n105_I_6_0_0_1 = n98_O_6_0_0_1; // @[Top.scala 127:12]
  assign n105_I_6_0_0_2 = n98_O_6_0_0_2; // @[Top.scala 127:12]
  assign n105_I_6_0_1_0 = n98_O_6_0_1_0; // @[Top.scala 127:12]
  assign n105_I_6_0_1_1 = n98_O_6_0_1_1; // @[Top.scala 127:12]
  assign n105_I_6_0_1_2 = n98_O_6_0_1_2; // @[Top.scala 127:12]
  assign n105_I_6_0_2_0 = n98_O_6_0_2_0; // @[Top.scala 127:12]
  assign n105_I_6_0_2_1 = n98_O_6_0_2_1; // @[Top.scala 127:12]
  assign n105_I_6_0_2_2 = n98_O_6_0_2_2; // @[Top.scala 127:12]
  assign n105_I_7_0_0_0 = n98_O_7_0_0_0; // @[Top.scala 127:12]
  assign n105_I_7_0_0_1 = n98_O_7_0_0_1; // @[Top.scala 127:12]
  assign n105_I_7_0_0_2 = n98_O_7_0_0_2; // @[Top.scala 127:12]
  assign n105_I_7_0_1_0 = n98_O_7_0_1_0; // @[Top.scala 127:12]
  assign n105_I_7_0_1_1 = n98_O_7_0_1_1; // @[Top.scala 127:12]
  assign n105_I_7_0_1_2 = n98_O_7_0_1_2; // @[Top.scala 127:12]
  assign n105_I_7_0_2_0 = n98_O_7_0_2_0; // @[Top.scala 127:12]
  assign n105_I_7_0_2_1 = n98_O_7_0_2_1; // @[Top.scala 127:12]
  assign n105_I_7_0_2_2 = n98_O_7_0_2_2; // @[Top.scala 127:12]
  assign n147_clock = clock;
  assign n147_reset = reset;
  assign n147_valid_up = n105_valid_down; // @[Top.scala 131:19]
  assign n147_I_0_0_0 = n105_O_0_0_0; // @[Top.scala 130:12]
  assign n147_I_0_0_1 = n105_O_0_0_1; // @[Top.scala 130:12]
  assign n147_I_0_0_2 = n105_O_0_0_2; // @[Top.scala 130:12]
  assign n147_I_0_1_0 = n105_O_0_1_0; // @[Top.scala 130:12]
  assign n147_I_0_1_1 = n105_O_0_1_1; // @[Top.scala 130:12]
  assign n147_I_0_1_2 = n105_O_0_1_2; // @[Top.scala 130:12]
  assign n147_I_0_2_0 = n105_O_0_2_0; // @[Top.scala 130:12]
  assign n147_I_0_2_1 = n105_O_0_2_1; // @[Top.scala 130:12]
  assign n147_I_0_2_2 = n105_O_0_2_2; // @[Top.scala 130:12]
  assign n147_I_1_0_0 = n105_O_1_0_0; // @[Top.scala 130:12]
  assign n147_I_1_0_1 = n105_O_1_0_1; // @[Top.scala 130:12]
  assign n147_I_1_0_2 = n105_O_1_0_2; // @[Top.scala 130:12]
  assign n147_I_1_1_0 = n105_O_1_1_0; // @[Top.scala 130:12]
  assign n147_I_1_1_1 = n105_O_1_1_1; // @[Top.scala 130:12]
  assign n147_I_1_1_2 = n105_O_1_1_2; // @[Top.scala 130:12]
  assign n147_I_1_2_0 = n105_O_1_2_0; // @[Top.scala 130:12]
  assign n147_I_1_2_1 = n105_O_1_2_1; // @[Top.scala 130:12]
  assign n147_I_1_2_2 = n105_O_1_2_2; // @[Top.scala 130:12]
  assign n147_I_2_0_0 = n105_O_2_0_0; // @[Top.scala 130:12]
  assign n147_I_2_0_1 = n105_O_2_0_1; // @[Top.scala 130:12]
  assign n147_I_2_0_2 = n105_O_2_0_2; // @[Top.scala 130:12]
  assign n147_I_2_1_0 = n105_O_2_1_0; // @[Top.scala 130:12]
  assign n147_I_2_1_1 = n105_O_2_1_1; // @[Top.scala 130:12]
  assign n147_I_2_1_2 = n105_O_2_1_2; // @[Top.scala 130:12]
  assign n147_I_2_2_0 = n105_O_2_2_0; // @[Top.scala 130:12]
  assign n147_I_2_2_1 = n105_O_2_2_1; // @[Top.scala 130:12]
  assign n147_I_2_2_2 = n105_O_2_2_2; // @[Top.scala 130:12]
  assign n147_I_3_0_0 = n105_O_3_0_0; // @[Top.scala 130:12]
  assign n147_I_3_0_1 = n105_O_3_0_1; // @[Top.scala 130:12]
  assign n147_I_3_0_2 = n105_O_3_0_2; // @[Top.scala 130:12]
  assign n147_I_3_1_0 = n105_O_3_1_0; // @[Top.scala 130:12]
  assign n147_I_3_1_1 = n105_O_3_1_1; // @[Top.scala 130:12]
  assign n147_I_3_1_2 = n105_O_3_1_2; // @[Top.scala 130:12]
  assign n147_I_3_2_0 = n105_O_3_2_0; // @[Top.scala 130:12]
  assign n147_I_3_2_1 = n105_O_3_2_1; // @[Top.scala 130:12]
  assign n147_I_3_2_2 = n105_O_3_2_2; // @[Top.scala 130:12]
  assign n147_I_4_0_0 = n105_O_4_0_0; // @[Top.scala 130:12]
  assign n147_I_4_0_1 = n105_O_4_0_1; // @[Top.scala 130:12]
  assign n147_I_4_0_2 = n105_O_4_0_2; // @[Top.scala 130:12]
  assign n147_I_4_1_0 = n105_O_4_1_0; // @[Top.scala 130:12]
  assign n147_I_4_1_1 = n105_O_4_1_1; // @[Top.scala 130:12]
  assign n147_I_4_1_2 = n105_O_4_1_2; // @[Top.scala 130:12]
  assign n147_I_4_2_0 = n105_O_4_2_0; // @[Top.scala 130:12]
  assign n147_I_4_2_1 = n105_O_4_2_1; // @[Top.scala 130:12]
  assign n147_I_4_2_2 = n105_O_4_2_2; // @[Top.scala 130:12]
  assign n147_I_5_0_0 = n105_O_5_0_0; // @[Top.scala 130:12]
  assign n147_I_5_0_1 = n105_O_5_0_1; // @[Top.scala 130:12]
  assign n147_I_5_0_2 = n105_O_5_0_2; // @[Top.scala 130:12]
  assign n147_I_5_1_0 = n105_O_5_1_0; // @[Top.scala 130:12]
  assign n147_I_5_1_1 = n105_O_5_1_1; // @[Top.scala 130:12]
  assign n147_I_5_1_2 = n105_O_5_1_2; // @[Top.scala 130:12]
  assign n147_I_5_2_0 = n105_O_5_2_0; // @[Top.scala 130:12]
  assign n147_I_5_2_1 = n105_O_5_2_1; // @[Top.scala 130:12]
  assign n147_I_5_2_2 = n105_O_5_2_2; // @[Top.scala 130:12]
  assign n147_I_6_0_0 = n105_O_6_0_0; // @[Top.scala 130:12]
  assign n147_I_6_0_1 = n105_O_6_0_1; // @[Top.scala 130:12]
  assign n147_I_6_0_2 = n105_O_6_0_2; // @[Top.scala 130:12]
  assign n147_I_6_1_0 = n105_O_6_1_0; // @[Top.scala 130:12]
  assign n147_I_6_1_1 = n105_O_6_1_1; // @[Top.scala 130:12]
  assign n147_I_6_1_2 = n105_O_6_1_2; // @[Top.scala 130:12]
  assign n147_I_6_2_0 = n105_O_6_2_0; // @[Top.scala 130:12]
  assign n147_I_6_2_1 = n105_O_6_2_1; // @[Top.scala 130:12]
  assign n147_I_6_2_2 = n105_O_6_2_2; // @[Top.scala 130:12]
  assign n147_I_7_0_0 = n105_O_7_0_0; // @[Top.scala 130:12]
  assign n147_I_7_0_1 = n105_O_7_0_1; // @[Top.scala 130:12]
  assign n147_I_7_0_2 = n105_O_7_0_2; // @[Top.scala 130:12]
  assign n147_I_7_1_0 = n105_O_7_1_0; // @[Top.scala 130:12]
  assign n147_I_7_1_1 = n105_O_7_1_1; // @[Top.scala 130:12]
  assign n147_I_7_1_2 = n105_O_7_1_2; // @[Top.scala 130:12]
  assign n147_I_7_2_0 = n105_O_7_2_0; // @[Top.scala 130:12]
  assign n147_I_7_2_1 = n105_O_7_2_1; // @[Top.scala 130:12]
  assign n147_I_7_2_2 = n105_O_7_2_2; // @[Top.scala 130:12]
  assign n148_valid_up = n147_valid_down; // @[Top.scala 134:19]
  assign n148_I_0_0_0 = n147_O_0_0_0; // @[Top.scala 133:12]
  assign n148_I_1_0_0 = n147_O_1_0_0; // @[Top.scala 133:12]
  assign n148_I_2_0_0 = n147_O_2_0_0; // @[Top.scala 133:12]
  assign n148_I_3_0_0 = n147_O_3_0_0; // @[Top.scala 133:12]
  assign n148_I_4_0_0 = n147_O_4_0_0; // @[Top.scala 133:12]
  assign n148_I_5_0_0 = n147_O_5_0_0; // @[Top.scala 133:12]
  assign n148_I_6_0_0 = n147_O_6_0_0; // @[Top.scala 133:12]
  assign n148_I_7_0_0 = n147_O_7_0_0; // @[Top.scala 133:12]
  assign n149_valid_up = n148_valid_down; // @[Top.scala 137:19]
  assign n149_I_0_0 = n148_O_0_0; // @[Top.scala 136:12]
  assign n149_I_1_0 = n148_O_1_0; // @[Top.scala 136:12]
  assign n149_I_2_0 = n148_O_2_0; // @[Top.scala 136:12]
  assign n149_I_3_0 = n148_O_3_0; // @[Top.scala 136:12]
  assign n149_I_4_0 = n148_O_4_0; // @[Top.scala 136:12]
  assign n149_I_5_0 = n148_O_5_0; // @[Top.scala 136:12]
  assign n149_I_6_0 = n148_O_6_0; // @[Top.scala 136:12]
  assign n149_I_7_0 = n148_O_7_0; // @[Top.scala 136:12]
  assign n150_clock = clock;
  assign n150_reset = reset;
  assign n150_valid_up = n149_valid_down; // @[Top.scala 140:19]
  assign n150_I_0 = n149_O_0; // @[Top.scala 139:12]
  assign n150_I_1 = n149_O_1; // @[Top.scala 139:12]
  assign n150_I_2 = n149_O_2; // @[Top.scala 139:12]
  assign n150_I_3 = n149_O_3; // @[Top.scala 139:12]
  assign n150_I_4 = n149_O_4; // @[Top.scala 139:12]
  assign n150_I_5 = n149_O_5; // @[Top.scala 139:12]
  assign n150_I_6 = n149_O_6; // @[Top.scala 139:12]
  assign n150_I_7 = n149_O_7; // @[Top.scala 139:12]
  assign n151_clock = clock;
  assign n151_reset = reset;
  assign n151_valid_up = n150_valid_down; // @[Top.scala 143:19]
  assign n151_I_0 = n150_O_0; // @[Top.scala 142:12]
  assign n151_I_1 = n150_O_1; // @[Top.scala 142:12]
  assign n151_I_2 = n150_O_2; // @[Top.scala 142:12]
  assign n151_I_3 = n150_O_3; // @[Top.scala 142:12]
  assign n151_I_4 = n150_O_4; // @[Top.scala 142:12]
  assign n151_I_5 = n150_O_5; // @[Top.scala 142:12]
  assign n151_I_6 = n150_O_6; // @[Top.scala 142:12]
  assign n151_I_7 = n150_O_7; // @[Top.scala 142:12]
  assign n152_clock = clock;
  assign n152_reset = reset;
  assign n152_valid_up = n151_valid_down; // @[Top.scala 146:19]
  assign n152_I_0 = n151_O_0; // @[Top.scala 145:12]
  assign n152_I_1 = n151_O_1; // @[Top.scala 145:12]
  assign n152_I_2 = n151_O_2; // @[Top.scala 145:12]
  assign n152_I_3 = n151_O_3; // @[Top.scala 145:12]
  assign n152_I_4 = n151_O_4; // @[Top.scala 145:12]
  assign n152_I_5 = n151_O_5; // @[Top.scala 145:12]
  assign n152_I_6 = n151_O_6; // @[Top.scala 145:12]
  assign n152_I_7 = n151_O_7; // @[Top.scala 145:12]
endmodule
