module stupleToSSeq_tInt_n3 (input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O_0 = I_0;
assign O_1 = I_1;
assign O_2 = I_2;
assign valid_down = valid_up;
endmodule

module sseqTupleCreator_tSSeq_3_Int_ (input [7:0] I0_0/*verilator public*/, input [7:0] I0_1/*verilator public*/, input [7:0] I0_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output [7:0] O_1_0/*verilator public*/, output [7:0] O_1_1/*verilator public*/, output [7:0] O_1_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O_0_0 = I0_0;
assign O_0_1 = I0_1;
assign O_0_2 = I0_2;
assign O_1_0 = I1_0;
assign O_1_1 = I1_1;
assign O_1_2 = I1_2;
assign valid_down = valid_up;
endmodule

module sseqTupleCreator_tInt (input [7:0] I0/*verilator public*/, input [7:0] I1/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O_0 = I0;
assign O_1 = I1;
assign valid_down = valid_up;
endmodule

module sseqTupleAppender_tSSeq_3_Int__n2 (input [7:0] I0_0_0/*verilator public*/, input [7:0] I0_0_1/*verilator public*/, input [7:0] I0_0_2/*verilator public*/, input [7:0] I0_1_0/*verilator public*/, input [7:0] I0_1_1/*verilator public*/, input [7:0] I0_1_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output [7:0] O_1_0/*verilator public*/, output [7:0] O_1_1/*verilator public*/, output [7:0] O_1_2/*verilator public*/, output [7:0] O_2_0/*verilator public*/, output [7:0] O_2_1/*verilator public*/, output [7:0] O_2_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O_0_0 = I0_0_0;
assign O_0_1 = I0_0_1;
assign O_0_2 = I0_0_2;
assign O_1_0 = I0_1_0;
assign O_1_1 = I0_1_1;
assign O_1_2 = I0_1_2;
assign O_2_0 = I1_0;
assign O_2_1 = I1_1;
assign O_2_2 = I1_2;
assign valid_down = valid_up;
endmodule

module sseqTupleAppender_tInt_n2 (input [7:0] I0_0/*verilator public*/, input [7:0] I0_1/*verilator public*/, input [7:0] I1/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O_0 = I0_0;
assign O_1 = I0_1;
assign O_2 = I1;
assign valid_down = valid_up;
endmodule

module corebit_xor (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 ^ in1;
endmodule

module corebit_term (input in/*verilator public*/);

endmodule

module corebit_not (input in/*verilator public*/, output out/*verilator public*/);
  assign out = ~in;
endmodule

module corebit_eq (input I0/*verilator public*/, input I1/*verilator public*/, output O/*verilator public*/);
wire not_inst0_out;
wire xor_inst0_out;
corebit_not not_inst0(.in(xor_inst0_out), .out(not_inst0_out));
corebit_xor xor_inst0(.in0(I0), .in1(I1), .out(xor_inst0_out));
assign O = not_inst0_out;
endmodule

module corebit_const #(parameter value = 1) (output out/*verilator public*/);
  assign out = value;
endmodule

module corebit_and (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 & in1;
endmodule

module atomTupleCreator_t0Int_t1Int (input [7:0] I0/*verilator public*/, input [7:0] I1/*verilator public*/, output [7:0] O__0/*verilator public*/, output [7:0] O__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O__0 = I0;
assign O__1 = I1;
assign valid_down = valid_up;
endmodule

module coreir_ult #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 < in1;
endmodule

module coreir_term #(parameter width = 1) (input [width-1:0] in/*verilator public*/);

endmodule

module coreir_slice #(parameter hi = 1, parameter lo = 0, parameter width = 1) (input [width-1:0] in/*verilator public*/, output [hi-lo-1:0] out/*verilator public*/);
  assign out = in[hi-1:lo];
endmodule

module coreir_shl #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = in0 << in1;
endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk/*verilator public*/, input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  reg [width-1:0] outReg/*verilator public*/=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_mux #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, input sel/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = sel ? in1 : in0;
endmodule

module coreir_mem #(parameter has_init = 0, parameter depth = 1, parameter width = 1) (input clk/*verilator public*/, input [width-1:0] wdata/*verilator public*/, input [$clog2(depth)-1:0] waddr/*verilator public*/, input wen/*verilator public*/, output [width-1:0] rdata/*verilator public*/, input [$clog2(depth)-1:0] raddr/*verilator public*/);
  reg [width-1:0] data[depth-1:0] /*verilator public*/;
  always @(posedge clk) begin
    if (wen) begin
      data[waddr] <= wdata;
    end
  end
  assign rdata = data[raddr];
endmodule

module coreir_lshr #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = in0 >> in1;
endmodule

module coreir_eq #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 == in1;
endmodule

module coreir_const #(parameter width = 1, parameter value = 1) (output [width-1:0] out/*verilator public*/);
  assign out = value;
endmodule

module coreir_add #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = in0 + in1;
endmodule

module \commonlib_muxn__N2__width8 (input [7:0] in_data_0/*verilator public*/, input [7:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [7:0] out/*verilator public*/);
wire [7:0] _join_out;
coreir_mux #(.width(8)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module \commonlib_muxn__N4__width8 (input [7:0] in_data_0/*verilator public*/, input [7:0] in_data_1/*verilator public*/, input [7:0] in_data_2/*verilator public*/, input [7:0] in_data_3/*verilator public*/, input [1:0] in_sel/*verilator public*/, output [7:0] out/*verilator public*/);
wire [7:0] _join_out;
wire [7:0] muxN_0_out;
wire [7:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(.width(8)) _join(.in0(muxN_0_out), .in1(muxN_1_out), .out(_join_out), .sel(in_sel[1]));
\commonlib_muxn__N2__width8 muxN_0(.in_data_0(in_data_0), .in_data_1(in_data_1), .in_sel(sel_slice0_out), .out(muxN_0_out));
\commonlib_muxn__N2__width8 muxN_1(.in_data_0(in_data_2), .in_data_1(in_data_3), .in_sel(sel_slice1_out), .out(muxN_1_out));
coreir_slice #(.hi(1), .lo(0), .width(2)) sel_slice0(.in(in_sel), .out(sel_slice0_out));
coreir_slice #(.hi(1), .lo(0), .width(2)) sel_slice1(.in(in_sel), .out(sel_slice1_out));
assign out = _join_out;
endmodule

module \commonlib_muxn__N2__width4 (input [3:0] in_data_0/*verilator public*/, input [3:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [3:0] out/*verilator public*/);
wire [3:0] _join_out;
coreir_mux #(.width(4)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module \commonlib_muxn__N2__width3 (input [2:0] in_data_0/*verilator public*/, input [2:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [2:0] out/*verilator public*/);
wire [2:0] _join_out;
coreir_mux #(.width(3)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module \commonlib_muxn__N2__width24 (input [23:0] in_data_0/*verilator public*/, input [23:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [23:0] out/*verilator public*/);
wire [23:0] _join_out;
coreir_mux #(.width(24)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module \commonlib_muxn__N2__width2 (input [1:0] in_data_0/*verilator public*/, input [1:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [1:0] out/*verilator public*/);
wire [1:0] _join_out;
coreir_mux #(.width(2)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module \commonlib_muxn__N2__width1 (input [0:0] in_data_0/*verilator public*/, input [0:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [0:0] out/*verilator public*/);
wire [0:0] _join_out;
coreir_mux #(.width(1)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module \commonlib_muxn__N1__width24 (input [23:0] in_data_0/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [23:0] out/*verilator public*/);
corebit_term term_sel(.in(in_sel[0]));
assign out = in_data_0;
endmodule

module \commonlib_muxn__N3__width24 (input [23:0] in_data_0/*verilator public*/, input [23:0] in_data_1/*verilator public*/, input [23:0] in_data_2/*verilator public*/, input [1:0] in_sel/*verilator public*/, output [23:0] out/*verilator public*/);
wire [23:0] _join_out;
wire [23:0] muxN_0_out;
wire [23:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(.width(24)) _join(.in0(muxN_0_out), .in1(muxN_1_out), .out(_join_out), .sel(in_sel[1]));
\commonlib_muxn__N2__width24 muxN_0(.in_data_0(in_data_0), .in_data_1(in_data_1), .in_sel(sel_slice0_out), .out(muxN_0_out));
\commonlib_muxn__N1__width24 muxN_1(.in_data_0(in_data_2), .in_sel(sel_slice1_out), .out(muxN_1_out));
coreir_slice #(.hi(1), .lo(0), .width(2)) sel_slice0(.in(in_sel), .out(sel_slice0_out));
coreir_slice #(.hi(1), .lo(0), .width(2)) sel_slice1(.in(in_sel), .out(sel_slice1_out));
assign out = _join_out;
endmodule

module lutN #(parameter N = 1, parameter init = 1) (input [N-1:0] in/*verilator public*/, output out/*verilator public*/);
  assign out = init[in];
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit83 (input [23:0] in/*verilator public*/, output [7:0] out_0/*verilator public*/, output [7:0] out_1/*verilator public*/, output [7:0] out_2/*verilator public*/);
assign out_0 = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
assign out_1 = {in[15],in[14],in[13],in[12],in[11],in[10],in[9],in[8]};
assign out_2 = {in[23],in[22],in[21],in[20],in[19],in[18],in[17],in[16]};
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit81 (input [7:0] in/*verilator public*/, output [7:0] out_0/*verilator public*/);
assign out_0 = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit83 (input [7:0] in_0/*verilator public*/, input [7:0] in_1/*verilator public*/, input [7:0] in_2/*verilator public*/, output [23:0] out/*verilator public*/);
assign out = {in_2[7],in_2[6],in_2[5],in_2[4],in_2[3],in_2[2],in_2[1],in_2[0],in_1[7],in_1[6],in_1[5],in_1[4],in_1[3],in_1[2],in_1[1],in_1[0],in_0[7],in_0[6],in_0[5],in_0[4],in_0[3],in_0[2],in_0[1],in_0[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit81 (input [7:0] in_0/*verilator public*/, output [7:0] out/*verilator public*/);
assign out = {in_0[7],in_0[6],in_0[5],in_0[4],in_0[3],in_0[2],in_0[1],in_0[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit2 (input [1:0] in/*verilator public*/, output [1:0] out/*verilator public*/);
assign out = {in[1],in[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit1 (input [0:0] in/*verilator public*/, output [0:0] out/*verilator public*/);
assign out = in[0];
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit (input in/*verilator public*/, output [0:0] out/*verilator public*/);
assign out = in;
endmodule

module Term_Bitt (input I/*verilator public*/);
wire [0:0] dehydrate_tBit_inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
coreir_term #(.width(1)) term_w1_inst0(.in(dehydrate_tBit_inst0_out));
endmodule

module Term_Bits_1_t (input [0:0] I/*verilator public*/);
wire [0:0] dehydrate_tBits_1__inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit1 dehydrate_tBits_1__inst0(.in(I), .out(dehydrate_tBits_1__inst0_out));
coreir_term #(.width(1)) term_w1_inst0(.in(dehydrate_tBits_1__inst0_out));
endmodule

module Term_Array_2_Bit_t (input [1:0] I/*verilator public*/);
wire [1:0] dehydrate_tArray_2_Bit__inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit2 dehydrate_tArray_2_Bit__inst0(.in(I), .out(dehydrate_tArray_2_Bit__inst0_out));
coreir_term #(.width(2)) term_w2_inst0(.in(dehydrate_tArray_2_Bit__inst0_out));
endmodule

module SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/);
wire [0:0] const_0_1_out;
Term_Bitt Term_Bitt_inst0(.I(CE));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
assign O = const_0_1_out;
endmodule

module Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ (input [7:0] I_0_0/*verilator public*/, input [7:0] I_0_1/*verilator public*/, input [7:0] I_0_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] stupleToSSeq_tInt_n3_inst0_O_0;
wire [7:0] stupleToSSeq_tInt_n3_inst0_O_1;
wire [7:0] stupleToSSeq_tInt_n3_inst0_O_2;
wire stupleToSSeq_tInt_n3_inst0_valid_down;
stupleToSSeq_tInt_n3 stupleToSSeq_tInt_n3_inst0(.I_0(I_0_0), .I_1(I_0_1), .I_2(I_0_2), .O_0(stupleToSSeq_tInt_n3_inst0_O_0), .O_1(stupleToSSeq_tInt_n3_inst0_O_1), .O_2(stupleToSSeq_tInt_n3_inst0_O_2), .valid_down(stupleToSSeq_tInt_n3_inst0_valid_down), .valid_up(valid_up));
assign O_0 = stupleToSSeq_tInt_n3_inst0_O_0;
assign O_1 = stupleToSSeq_tInt_n3_inst0_O_1;
assign O_2 = stupleToSSeq_tInt_n3_inst0_O_2;
assign valid_down = stupleToSSeq_tInt_n3_inst0_valid_down;
endmodule

module RShift_Atom (input [7:0] I__0/*verilator public*/, input [7:0] I__1/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] lshr8_inst0_out;
coreir_lshr #(.width(8)) lshr8_inst0(.in0(I__0), .in1(I__1), .out(lshr8_inst0_out));
assign O = lshr8_inst0_out;
assign valid_down = valid_up;
endmodule

module RAM1x8 (input CLK/*verilator public*/, input [0:0] RADDR/*verilator public*/, output [7:0] RDATA/*verilator public*/, input [0:0] WADDR/*verilator public*/, input [7:0] WDATA/*verilator public*/, input WE/*verilator public*/);
wire [7:0] coreir_mem1x8_inst0_rdata;
coreir_mem #(.depth(1), .has_init(0), .width(8)) coreir_mem1x8_inst0(.clk(CLK), .raddr(RADDR), .rdata(coreir_mem1x8_inst0_rdata), .waddr(WADDR), .wdata(WDATA), .wen(WE));
assign RDATA = coreir_mem1x8_inst0_rdata;
endmodule

module RAM_Array_1_Array_8_Bit__t_1n (input CLK/*verilator public*/, input [0:0] RADDR/*verilator public*/, output [7:0] RDATA_0/*verilator public*/, input [0:0] WADDR/*verilator public*/, input [7:0] WDATA_0/*verilator public*/, input WE/*verilator public*/);
wire [7:0] RAM1x8_inst0_RDATA;
wire [7:0] dehydrate_tArray_1_Array_8_Bit___inst0_out;
wire [7:0] hydrate_tArray_1_Array_8_Bit___inst0_out_0;
RAM1x8 RAM1x8_inst0(.CLK(CLK), .RADDR(RADDR), .RDATA(RAM1x8_inst0_RDATA), .WADDR(WADDR), .WDATA(dehydrate_tArray_1_Array_8_Bit___inst0_out), .WE(WE));
\aetherlinglib_dehydrate__hydratedTypeBit81 dehydrate_tArray_1_Array_8_Bit___inst0(.in_0(WDATA_0), .out(dehydrate_tArray_1_Array_8_Bit___inst0_out));
\aetherlinglib_hydrate__hydratedTypeBit81 hydrate_tArray_1_Array_8_Bit___inst0(.in(RAM1x8_inst0_RDATA), .out_0(hydrate_tArray_1_Array_8_Bit___inst0_out_0));
assign RDATA_0 = hydrate_tArray_1_Array_8_Bit___inst0_out_0;
endmodule

module NestedCounters_Int_hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output last/*verilator public*/, output valid/*verilator public*/);
wire [0:0] coreir_const11_inst0_out;
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign last = coreir_const11_inst0_out[0];
assign valid = CE;
endmodule

module NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output last/*verilator public*/, output valid/*verilator public*/);
wire NestedCounters_Int_hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_Int_hasCETrue_hasResetFalse_inst0_valid;
NestedCounters_Int_hasCETrue_hasResetFalse NestedCounters_Int_hasCETrue_hasResetFalse_inst0(.CE(CE), .CLK(CLK), .last(NestedCounters_Int_hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_Int_hasCETrue_hasResetFalse_inst0_valid));
assign last = NestedCounters_Int_hasCETrue_hasResetFalse_inst0_last;
assign valid = NestedCounters_Int_hasCETrue_hasResetFalse_inst0_valid;
endmodule

module NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit___ (input [7:0] I_0_0/*verilator public*/, input [7:0] I_1_0/*verilator public*/, input [7:0] I_2_0/*verilator public*/, input [7:0] I_3_0/*verilator public*/, output [7:0] out_0/*verilator public*/, output [7:0] out_1/*verilator public*/, output [7:0] out_2/*verilator public*/, output [7:0] out_3/*verilator public*/);
wire [7:0] dehydrate_tArray_1_Array_8_Bit___inst0_out;
wire [7:0] dehydrate_tArray_1_Array_8_Bit___inst1_out;
wire [7:0] dehydrate_tArray_1_Array_8_Bit___inst2_out;
wire [7:0] dehydrate_tArray_1_Array_8_Bit___inst3_out;
\aetherlinglib_dehydrate__hydratedTypeBit81 dehydrate_tArray_1_Array_8_Bit___inst0(.in_0(I_0_0), .out(dehydrate_tArray_1_Array_8_Bit___inst0_out));
\aetherlinglib_dehydrate__hydratedTypeBit81 dehydrate_tArray_1_Array_8_Bit___inst1(.in_0(I_1_0), .out(dehydrate_tArray_1_Array_8_Bit___inst1_out));
\aetherlinglib_dehydrate__hydratedTypeBit81 dehydrate_tArray_1_Array_8_Bit___inst2(.in_0(I_2_0), .out(dehydrate_tArray_1_Array_8_Bit___inst2_out));
\aetherlinglib_dehydrate__hydratedTypeBit81 dehydrate_tArray_1_Array_8_Bit___inst3(.in_0(I_3_0), .out(dehydrate_tArray_1_Array_8_Bit___inst3_out));
assign out_0 = dehydrate_tArray_1_Array_8_Bit___inst0_out;
assign out_1 = dehydrate_tArray_1_Array_8_Bit___inst1_out;
assign out_2 = dehydrate_tArray_1_Array_8_Bit___inst2_out;
assign out_3 = dehydrate_tArray_1_Array_8_Bit___inst3_out;
endmodule

module NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit___ (input [7:0] I_0_0/*verilator public*/, input [7:0] I_0_1/*verilator public*/, input [7:0] I_0_2/*verilator public*/, input [7:0] I_1_0/*verilator public*/, input [7:0] I_1_1/*verilator public*/, input [7:0] I_1_2/*verilator public*/, input [7:0] I_2_0/*verilator public*/, input [7:0] I_2_1/*verilator public*/, input [7:0] I_2_2/*verilator public*/, output [23:0] out_0/*verilator public*/, output [23:0] out_1/*verilator public*/, output [23:0] out_2/*verilator public*/);
wire [23:0] dehydrate_tArray_3_Array_8_Bit___inst0_out;
wire [23:0] dehydrate_tArray_3_Array_8_Bit___inst1_out;
wire [23:0] dehydrate_tArray_3_Array_8_Bit___inst2_out;
\aetherlinglib_dehydrate__hydratedTypeBit83 dehydrate_tArray_3_Array_8_Bit___inst0(.in_0(I_0_0), .in_1(I_0_1), .in_2(I_0_2), .out(dehydrate_tArray_3_Array_8_Bit___inst0_out));
\aetherlinglib_dehydrate__hydratedTypeBit83 dehydrate_tArray_3_Array_8_Bit___inst1(.in_0(I_1_0), .in_1(I_1_1), .in_2(I_1_2), .out(dehydrate_tArray_3_Array_8_Bit___inst1_out));
\aetherlinglib_dehydrate__hydratedTypeBit83 dehydrate_tArray_3_Array_8_Bit___inst2(.in_0(I_2_0), .in_1(I_2_1), .in_2(I_2_2), .out(dehydrate_tArray_3_Array_8_Bit___inst2_out));
assign out_0 = dehydrate_tArray_3_Array_8_Bit___inst0_out;
assign out_1 = dehydrate_tArray_3_Array_8_Bit___inst1_out;
assign out_2 = dehydrate_tArray_3_Array_8_Bit___inst2_out;
endmodule

module NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ (input [7:0] I0_0/*verilator public*/, input [7:0] I0_1/*verilator public*/, input [7:0] I0_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0__0/*verilator public*/, output [7:0] O_0__1/*verilator public*/, output [7:0] O_1__0/*verilator public*/, output [7:0] O_1__1/*verilator public*/, output [7:0] O_2__0/*verilator public*/, output [7:0] O_2__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire and_inst0_out;
wire and_inst1_out;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst1_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst1_O__1;
wire atomTupleCreator_t0Int_t1Int_inst1_valid_down;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst2_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst2_O__1;
wire atomTupleCreator_t0Int_t1Int_inst2_valid_down;
corebit_and and_inst0(.in0(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .in1(atomTupleCreator_t0Int_t1Int_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(atomTupleCreator_t0Int_t1Int_inst2_valid_down), .out(and_inst1_out));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I0_0), .I1(I1_0), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(valid_up));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst1(.I0(I0_1), .I1(I1_1), .O__0(atomTupleCreator_t0Int_t1Int_inst1_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst1_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst1_valid_down), .valid_up(valid_up));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst2(.I0(I0_2), .I1(I1_2), .O__0(atomTupleCreator_t0Int_t1Int_inst2_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst2_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst2_valid_down), .valid_up(valid_up));
assign O_0__0 = atomTupleCreator_t0Int_t1Int_inst0_O__0;
assign O_0__1 = atomTupleCreator_t0Int_t1Int_inst0_O__1;
assign O_1__0 = atomTupleCreator_t0Int_t1Int_inst1_O__0;
assign O_1__1 = atomTupleCreator_t0Int_t1Int_inst1_O__1;
assign O_2__0 = atomTupleCreator_t0Int_t1Int_inst2_O__0;
assign O_2__1 = atomTupleCreator_t0Int_t1Int_inst2_O__1;
assign valid_down = and_inst1_out;
endmodule

module NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit___ (input [7:0] I_0_0/*verilator public*/, input [7:0] I_0_1/*verilator public*/, input [7:0] I_0_2/*verilator public*/, input [7:0] I_1_0/*verilator public*/, input [7:0] I_1_1/*verilator public*/, input [7:0] I_1_2/*verilator public*/, output [23:0] out_0/*verilator public*/, output [23:0] out_1/*verilator public*/);
wire [23:0] dehydrate_tArray_3_Array_8_Bit___inst0_out;
wire [23:0] dehydrate_tArray_3_Array_8_Bit___inst1_out;
\aetherlinglib_dehydrate__hydratedTypeBit83 dehydrate_tArray_3_Array_8_Bit___inst0(.in_0(I_0_0), .in_1(I_0_1), .in_2(I_0_2), .out(dehydrate_tArray_3_Array_8_Bit___inst0_out));
\aetherlinglib_dehydrate__hydratedTypeBit83 dehydrate_tArray_3_Array_8_Bit___inst1(.in_0(I_1_0), .in_1(I_1_1), .in_2(I_1_2), .out(dehydrate_tArray_3_Array_8_Bit___inst1_out));
assign out_0 = dehydrate_tArray_3_Array_8_Bit___inst0_out;
assign out_1 = dehydrate_tArray_3_Array_8_Bit___inst1_out;
endmodule

module NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit___ (input [7:0] I_0_0/*verilator public*/, input [7:0] I_1_0/*verilator public*/, output [7:0] out_0/*verilator public*/, output [7:0] out_1/*verilator public*/);
wire [7:0] dehydrate_tArray_1_Array_8_Out_Bit____inst0_out;
wire [7:0] dehydrate_tArray_1_Array_8_Out_Bit____inst1_out;
\aetherlinglib_dehydrate__hydratedTypeBit81 dehydrate_tArray_1_Array_8_Out_Bit____inst0(.in_0(I_0_0), .out(dehydrate_tArray_1_Array_8_Out_Bit____inst0_out));
\aetherlinglib_dehydrate__hydratedTypeBit81 dehydrate_tArray_1_Array_8_Out_Bit____inst1(.in_0(I_1_0), .out(dehydrate_tArray_1_Array_8_Out_Bit____inst1_out));
assign out_0 = dehydrate_tArray_1_Array_8_Out_Bit____inst0_out;
assign out_1 = dehydrate_tArray_1_Array_8_Out_Bit____inst1_out;
endmodule

module NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ (input [7:0] I0_0/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] sseqTupleCreator_tInt_inst0_O_0;
wire [7:0] sseqTupleCreator_tInt_inst0_O_1;
wire sseqTupleCreator_tInt_inst0_valid_down;
sseqTupleCreator_tInt sseqTupleCreator_tInt_inst0(.I0(I0_0), .I1(I1_0), .O_0(sseqTupleCreator_tInt_inst0_O_0), .O_1(sseqTupleCreator_tInt_inst0_O_1), .valid_down(sseqTupleCreator_tInt_inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = sseqTupleCreator_tInt_inst0_O_0;
assign O_0_1 = sseqTupleCreator_tInt_inst0_O_1;
assign valid_down = sseqTupleCreator_tInt_inst0_valid_down;
endmodule

module NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ (input [7:0] I0_0_0/*verilator public*/, input [7:0] I0_0_1/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] sseqTupleAppender_tInt_n2_inst0_O_0;
wire [7:0] sseqTupleAppender_tInt_n2_inst0_O_1;
wire [7:0] sseqTupleAppender_tInt_n2_inst0_O_2;
wire sseqTupleAppender_tInt_n2_inst0_valid_down;
sseqTupleAppender_tInt_n2 sseqTupleAppender_tInt_n2_inst0(.I0_0(I0_0_0), .I0_1(I0_0_1), .I1(I1_0), .O_0(sseqTupleAppender_tInt_n2_inst0_O_0), .O_1(sseqTupleAppender_tInt_n2_inst0_O_1), .O_2(sseqTupleAppender_tInt_n2_inst0_O_2), .valid_down(sseqTupleAppender_tInt_n2_inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = sseqTupleAppender_tInt_n2_inst0_O_0;
assign O_0_1 = sseqTupleAppender_tInt_n2_inst0_O_1;
assign O_0_2 = sseqTupleAppender_tInt_n2_inst0_O_2;
assign valid_down = sseqTupleAppender_tInt_n2_inst0_valid_down;
endmodule

module NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ (input [7:0] I0_0/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0__0/*verilator public*/, output [7:0] O_0__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I0_0), .I1(I1_0), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(valid_up));
assign O_0__0 = atomTupleCreator_t0Int_t1Int_inst0_O__0;
assign O_0__1 = atomTupleCreator_t0Int_t1Int_inst0_O__1;
assign valid_down = atomTupleCreator_t0Int_t1Int_inst0_valid_down;
endmodule

module NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit__ (input [7:0] I_0__0/*verilator public*/, input [7:0] I_0__1/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] RShift_Atom_inst0_O;
wire RShift_Atom_inst0_valid_down;
RShift_Atom RShift_Atom_inst0(.I__0(I_0__0), .I__1(I_0__1), .O(RShift_Atom_inst0_O), .valid_down(RShift_Atom_inst0_valid_down), .valid_up(valid_up));
assign O_0 = RShift_Atom_inst0_O;
assign valid_down = RShift_Atom_inst0_valid_down;
endmodule

module Mux_Array_3_Array_8_Bit__t_3n (input [7:0] data_0_0/*verilator public*/, input [7:0] data_0_1/*verilator public*/, input [7:0] data_0_2/*verilator public*/, input [7:0] data_1_0/*verilator public*/, input [7:0] data_1_1/*verilator public*/, input [7:0] data_1_2/*verilator public*/, input [7:0] data_2_0/*verilator public*/, input [7:0] data_2_1/*verilator public*/, input [7:0] data_2_2/*verilator public*/, output [7:0] out_0/*verilator public*/, output [7:0] out_1/*verilator public*/, output [7:0] out_2/*verilator public*/, input [1:0] sel/*verilator public*/);
wire [23:0] CommonlibMuxN_n3_w24_inst0_out;
wire [23:0] NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_0;
wire [23:0] NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_1;
wire [23:0] NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_2;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_0;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_1;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_2;
\commonlib_muxn__N3__width24 CommonlibMuxN_n3_w24_inst0(.in_data_0(NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_0), .in_data_1(NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_1), .in_data_2(NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_2), .in_sel(sel), .out(CommonlibMuxN_n3_w24_inst0_out));
NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit___ NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0(.I_0_0(data_0_0), .I_0_1(data_0_1), .I_0_2(data_0_2), .I_1_0(data_1_0), .I_1_1(data_1_1), .I_1_2(data_1_2), .I_2_0(data_2_0), .I_2_1(data_2_1), .I_2_2(data_2_2), .out_0(NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_0), .out_1(NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_1), .out_2(NativeMapParallel_n3_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_2));
\aetherlinglib_hydrate__hydratedTypeBit83 hydrate_tArray_3_Array_8_Bit___inst0(.in(CommonlibMuxN_n3_w24_inst0_out), .out_0(hydrate_tArray_3_Array_8_Bit___inst0_out_0), .out_1(hydrate_tArray_3_Array_8_Bit___inst0_out_1), .out_2(hydrate_tArray_3_Array_8_Bit___inst0_out_2));
assign out_0 = hydrate_tArray_3_Array_8_Bit___inst0_out_0;
assign out_1 = hydrate_tArray_3_Array_8_Bit___inst0_out_1;
assign out_2 = hydrate_tArray_3_Array_8_Bit___inst0_out_2;
endmodule

module Mux_Array_3_Array_8_Bit__t_2n (input [7:0] data_0_0/*verilator public*/, input [7:0] data_0_1/*verilator public*/, input [7:0] data_0_2/*verilator public*/, input [7:0] data_1_0/*verilator public*/, input [7:0] data_1_1/*verilator public*/, input [7:0] data_1_2/*verilator public*/, output [7:0] out_0/*verilator public*/, output [7:0] out_1/*verilator public*/, output [7:0] out_2/*verilator public*/, input [0:0] sel/*verilator public*/);
wire [23:0] CommonlibMuxN_n2_w24_inst0_out;
wire [23:0] NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_0;
wire [23:0] NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_1;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_0;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_1;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_2;
\commonlib_muxn__N2__width24 CommonlibMuxN_n2_w24_inst0(.in_data_0(NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_0), .in_data_1(NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_1), .in_sel(sel), .out(CommonlibMuxN_n2_w24_inst0_out));
NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit___ NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0(.I_0_0(data_0_0), .I_0_1(data_0_1), .I_0_2(data_0_2), .I_1_0(data_1_0), .I_1_1(data_1_1), .I_1_2(data_1_2), .out_0(NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_0), .out_1(NativeMapParallel_n2_opdehydrate_tArray_3_Array_8_Bit___I_Array_3_Array_8_In_Bit____out_Array_24_Out_Bit____inst0_out_1));
\aetherlinglib_hydrate__hydratedTypeBit83 hydrate_tArray_3_Array_8_Bit___inst0(.in(CommonlibMuxN_n2_w24_inst0_out), .out_0(hydrate_tArray_3_Array_8_Bit___inst0_out_0), .out_1(hydrate_tArray_3_Array_8_Bit___inst0_out_1), .out_2(hydrate_tArray_3_Array_8_Bit___inst0_out_2));
assign out_0 = hydrate_tArray_3_Array_8_Bit___inst0_out_0;
assign out_1 = hydrate_tArray_3_Array_8_Bit___inst0_out_1;
assign out_2 = hydrate_tArray_3_Array_8_Bit___inst0_out_2;
endmodule

module Mux_Array_1_Array_8_Out_Bit___t_2n (input [7:0] data_0_0/*verilator public*/, input [7:0] data_1_0/*verilator public*/, output [7:0] out_0/*verilator public*/, input [0:0] sel/*verilator public*/);
wire [7:0] CommonlibMuxN_n2_w8_inst0_out;
wire [7:0] NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_0;
wire [7:0] NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_1;
wire [7:0] hydrate_tArray_1_Array_8_Out_Bit____inst0_out_0;
\commonlib_muxn__N2__width8 CommonlibMuxN_n2_w8_inst0(.in_data_0(NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_0), .in_data_1(NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_1), .in_sel(sel), .out(CommonlibMuxN_n2_w8_inst0_out));
NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit___ NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0(.I_0_0(data_0_0), .I_1_0(data_1_0), .out_0(NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_0), .out_1(NativeMapParallel_n2_opdehydrate_tArray_1_Array_8_Out_Bit____I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_1));
\aetherlinglib_hydrate__hydratedTypeBit81 hydrate_tArray_1_Array_8_Out_Bit____inst0(.in(CommonlibMuxN_n2_w8_inst0_out), .out_0(hydrate_tArray_1_Array_8_Out_Bit____inst0_out_0));
assign out_0 = hydrate_tArray_1_Array_8_Out_Bit____inst0_out_0;
endmodule

module Mux_Array_1_Array_8_Bit__t_4n (input [7:0] data_0_0/*verilator public*/, input [7:0] data_1_0/*verilator public*/, input [7:0] data_2_0/*verilator public*/, input [7:0] data_3_0/*verilator public*/, output [7:0] out_0/*verilator public*/, input [1:0] sel/*verilator public*/);
wire [7:0] CommonlibMuxN_n4_w8_inst0_out;
wire [7:0] NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_0;
wire [7:0] NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_1;
wire [7:0] NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_2;
wire [7:0] NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_3;
wire [7:0] hydrate_tArray_1_Array_8_Bit___inst0_out_0;
\commonlib_muxn__N4__width8 CommonlibMuxN_n4_w8_inst0(.in_data_0(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_0), .in_data_1(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_1), .in_data_2(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_2), .in_data_3(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_3), .in_sel(sel), .out(CommonlibMuxN_n4_w8_inst0_out));
NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit___ NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0(.I_0_0(data_0_0), .I_1_0(data_1_0), .I_2_0(data_2_0), .I_3_0(data_3_0), .out_0(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_0), .out_1(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_1), .out_2(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_2), .out_3(NativeMapParallel_n4_opdehydrate_tArray_1_Array_8_Bit___I_Array_1_Array_8_In_Bit____out_Array_8_Out_Bit____inst0_out_3));
\aetherlinglib_hydrate__hydratedTypeBit81 hydrate_tArray_1_Array_8_Bit___inst0(.in(CommonlibMuxN_n4_w8_inst0_out), .out_0(hydrate_tArray_1_Array_8_Bit___inst0_out_0));
assign out_0 = hydrate_tArray_1_Array_8_Bit___inst0_out_0;
endmodule

module Mux_Array_1_Array_8_Bit__t_1n (input [7:0] data_0_0/*verilator public*/, output [7:0] out_0/*verilator public*/, input [0:0] sel/*verilator public*/);
Term_Bits_1_t Term_Bits_1_t_inst0(.I(sel));
assign out_0 = data_0_0;
endmodule

module Mux2xOutBits4 (input [3:0] I0/*verilator public*/, input [3:0] I1/*verilator public*/, output [3:0] O/*verilator public*/, input S/*verilator public*/);
wire [3:0] coreir_commonlib_mux2x4_inst0_out;
\commonlib_muxn__N2__width4 coreir_commonlib_mux2x4_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x4_inst0_out));
assign O = coreir_commonlib_mux2x4_inst0_out;
endmodule

module Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_4 (input CE/*verilator public*/, input CLK/*verilator public*/, input [3:0] I/*verilator public*/, output [3:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [3:0] Mux2xOutBits4_inst0_O;
wire [3:0] const_0_4_out;
wire [3:0] enable_mux_O;
wire [3:0] value_out;
Mux2xOutBits4 Mux2xOutBits4_inst0(.I0(enable_mux_O), .I1(const_0_4_out), .O(Mux2xOutBits4_inst0_O), .S(RESET));
coreir_const #(.value(4'h0), .width(4)) const_0_4(.out(const_0_4_out));
Mux2xOutBits4 enable_mux(.I0(value_out), .I1(I), .O(enable_mux_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(4'h0), .width(4)) value(.clk(CLK), .in(Mux2xOutBits4_inst0_O), .out(value_out));
assign O = value_out;
endmodule

module Mux2xOutBits3 (input [2:0] I0/*verilator public*/, input [2:0] I1/*verilator public*/, output [2:0] O/*verilator public*/, input S/*verilator public*/);
wire [2:0] coreir_commonlib_mux2x3_inst0_out;
\commonlib_muxn__N2__width3 coreir_commonlib_mux2x3_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x3_inst0_out));
assign O = coreir_commonlib_mux2x3_inst0_out;
endmodule

module Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3 (input CE/*verilator public*/, input CLK/*verilator public*/, input [2:0] I/*verilator public*/, output [2:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [2:0] Mux2xOutBits3_inst0_O;
wire [2:0] const_0_3_out;
wire [2:0] enable_mux_O;
wire [2:0] value_out;
Mux2xOutBits3 Mux2xOutBits3_inst0(.I0(enable_mux_O), .I1(const_0_3_out), .O(Mux2xOutBits3_inst0_O), .S(RESET));
coreir_const #(.value(3'h0), .width(3)) const_0_3(.out(const_0_3_out));
Mux2xOutBits3 enable_mux(.I0(value_out), .I1(I), .O(enable_mux_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(3'h0), .width(3)) value(.clk(CLK), .in(Mux2xOutBits3_inst0_O), .out(value_out));
assign O = value_out;
endmodule

module Mux2xOutBits2 (input [1:0] I0/*verilator public*/, input [1:0] I1/*verilator public*/, output [1:0] O/*verilator public*/, input S/*verilator public*/);
wire [1:0] coreir_commonlib_mux2x2_inst0_out;
\commonlib_muxn__N2__width2 coreir_commonlib_mux2x2_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x2_inst0_out));
assign O = coreir_commonlib_mux2x2_inst0_out;
endmodule

module Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2 (input CE/*verilator public*/, input CLK/*verilator public*/, input [1:0] I/*verilator public*/, output [1:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [1:0] Mux2xOutBits2_inst0_O;
wire [1:0] const_0_2_out;
wire [1:0] enable_mux_O;
wire [1:0] value_out;
Mux2xOutBits2 Mux2xOutBits2_inst0(.I0(enable_mux_O), .I1(const_0_2_out), .O(Mux2xOutBits2_inst0_O), .S(RESET));
coreir_const #(.value(2'h0), .width(2)) const_0_2(.out(const_0_2_out));
Mux2xOutBits2 enable_mux(.I0(value_out), .I1(I), .O(enable_mux_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(2'h0), .width(2)) value(.clk(CLK), .in(Mux2xOutBits2_inst0_O), .out(value_out));
assign O = value_out;
endmodule

module Mux2xNone (input I0/*verilator public*/, input I1/*verilator public*/, output O/*verilator public*/, input S/*verilator public*/);
wire [0:0] coreir_commonlib_mux2x1_inst0_out;
\commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x1_inst0_out));
assign O = coreir_commonlib_mux2x1_inst0_out[0];
endmodule

module Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I0_0/*verilator public*/, input [7:0] I0_1/*verilator public*/, input [7:0] I0_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0__0/*verilator public*/, output [7:0] O_0__1/*verilator public*/, output [7:0] O_1__0/*verilator public*/, output [7:0] O_1__1/*verilator public*/, output [7:0] O_2__0/*verilator public*/, output [7:0] O_2__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__0;
wire [7:0] NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__1;
wire [7:0] NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1__0;
wire [7:0] NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1__1;
wire [7:0] NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2__0;
wire [7:0] NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2__1;
wire NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0(.I0_0(I0_0), .I0_1(I0_1), .I0_2(I0_2), .I1_0(I1_0), .I1_1(I1_1), .I1_2(I1_2), .O_0__0(NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__0), .O_0__1(NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__1), .O_1__0(NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1__0), .O_1__1(NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1__1), .O_2__0(NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2__0), .O_2__1(NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2__1), .valid_down(NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0__0 = NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__0;
assign O_0__1 = NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__1;
assign O_1__0 = NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1__0;
assign O_1__1 = NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1__1;
assign O_2__0 = NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2__0;
assign O_2__1 = NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2__1;
assign valid_down = NativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I0_0/*verilator public*/, input [7:0] I0_1/*verilator public*/, input [7:0] I0_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output [7:0] O_1_0/*verilator public*/, output [7:0] O_1_1/*verilator public*/, output [7:0] O_1_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] sseqTupleCreator_tSSeq_3_Int__inst0_O_0_0;
wire [7:0] sseqTupleCreator_tSSeq_3_Int__inst0_O_0_1;
wire [7:0] sseqTupleCreator_tSSeq_3_Int__inst0_O_0_2;
wire [7:0] sseqTupleCreator_tSSeq_3_Int__inst0_O_1_0;
wire [7:0] sseqTupleCreator_tSSeq_3_Int__inst0_O_1_1;
wire [7:0] sseqTupleCreator_tSSeq_3_Int__inst0_O_1_2;
wire sseqTupleCreator_tSSeq_3_Int__inst0_valid_down;
sseqTupleCreator_tSSeq_3_Int_ sseqTupleCreator_tSSeq_3_Int__inst0(.I0_0(I0_0), .I0_1(I0_1), .I0_2(I0_2), .I1_0(I1_0), .I1_1(I1_1), .I1_2(I1_2), .O_0_0(sseqTupleCreator_tSSeq_3_Int__inst0_O_0_0), .O_0_1(sseqTupleCreator_tSSeq_3_Int__inst0_O_0_1), .O_0_2(sseqTupleCreator_tSSeq_3_Int__inst0_O_0_2), .O_1_0(sseqTupleCreator_tSSeq_3_Int__inst0_O_1_0), .O_1_1(sseqTupleCreator_tSSeq_3_Int__inst0_O_1_1), .O_1_2(sseqTupleCreator_tSSeq_3_Int__inst0_O_1_2), .valid_down(sseqTupleCreator_tSSeq_3_Int__inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = sseqTupleCreator_tSSeq_3_Int__inst0_O_0_0;
assign O_0_1 = sseqTupleCreator_tSSeq_3_Int__inst0_O_0_1;
assign O_0_2 = sseqTupleCreator_tSSeq_3_Int__inst0_O_0_2;
assign O_1_0 = sseqTupleCreator_tSSeq_3_Int__inst0_O_1_0;
assign O_1_1 = sseqTupleCreator_tSSeq_3_Int__inst0_O_1_1;
assign O_1_2 = sseqTupleCreator_tSSeq_3_Int__inst0_O_1_2;
assign valid_down = sseqTupleCreator_tSSeq_3_Int__inst0_valid_down;
endmodule

module Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I0_0_0/*verilator public*/, input [7:0] I0_0_1/*verilator public*/, input [7:0] I0_0_2/*verilator public*/, input [7:0] I0_1_0/*verilator public*/, input [7:0] I0_1_1/*verilator public*/, input [7:0] I0_1_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output [7:0] O_1_0/*verilator public*/, output [7:0] O_1_1/*verilator public*/, output [7:0] O_1_2/*verilator public*/, output [7:0] O_2_0/*verilator public*/, output [7:0] O_2_1/*verilator public*/, output [7:0] O_2_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_0;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_1;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_2;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_0;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_1;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_2;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_0;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_1;
wire [7:0] sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_2;
wire sseqTupleAppender_tSSeq_3_Int__n2_inst0_valid_down;
sseqTupleAppender_tSSeq_3_Int__n2 sseqTupleAppender_tSSeq_3_Int__n2_inst0(.I0_0_0(I0_0_0), .I0_0_1(I0_0_1), .I0_0_2(I0_0_2), .I0_1_0(I0_1_0), .I0_1_1(I0_1_1), .I0_1_2(I0_1_2), .I1_0(I1_0), .I1_1(I1_1), .I1_2(I1_2), .O_0_0(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_0), .O_0_1(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_1), .O_0_2(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_2), .O_1_0(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_0), .O_1_1(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_1), .O_1_2(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_2), .O_2_0(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_0), .O_2_1(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_1), .O_2_2(sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_2), .valid_down(sseqTupleAppender_tSSeq_3_Int__n2_inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_0;
assign O_0_1 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_1;
assign O_0_2 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_0_2;
assign O_1_0 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_0;
assign O_1_1 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_1;
assign O_1_2 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_1_2;
assign O_2_0 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_0;
assign O_2_1 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_1;
assign O_2_2 = sseqTupleAppender_tSSeq_3_Int__n2_inst0_O_2_2;
assign valid_down = sseqTupleAppender_tSSeq_3_Int__n2_inst0_valid_down;
endmodule

module Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I_0_0/*verilator public*/, input [7:0] I_0_1/*verilator public*/, input [7:0] I_0_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0(.I_0_0(I_0_0), .I_0_1(I_0_1), .I_0_2(I_0_2), .O_0(Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_2(Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .valid_down(Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0 = Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
assign O_1 = Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
assign O_2 = Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
assign valid_down = Remove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit____O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I0_0/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_0;
wire [7:0] NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_1;
wire NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0(.I0_0(I0_0), .I1_0(I1_0), .O_0_0(NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_0), .O_0_1(NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_1), .valid_down(NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_0;
assign O_0_1 = NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_1;
assign valid_down = NativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Array_2_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I0_0_0/*verilator public*/, input [7:0] I0_0_1/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_0;
wire [7:0] NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_1;
wire [7:0] NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_2;
wire NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0(.I0_0_0(I0_0_0), .I0_0_1(I0_0_1), .I1_0(I1_0), .O_0_0(NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_0), .O_0_1(NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_1), .O_0_2(NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_2), .valid_down(NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_0;
assign O_0_1 = NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_1;
assign O_0_2 = NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0_2;
assign valid_down = NativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit____I1_Array_8_In_Bit___O_Array_3_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I0_0/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0__0/*verilator public*/, output [7:0] O_0__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__0;
wire [7:0] NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__1;
wire NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0(.I0_0(I0_0), .I1_0(I1_0), .O_0__0(NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__0), .O_0__1(NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__1), .valid_down(NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0__0 = NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__0;
assign O_0__1 = NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0__1;
assign valid_down = NativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit___I1_Array_8_In_Bit___O_Tuple_0_Array_8_Out_Bit___1_Array_8_Out_Bit____valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I_0__0/*verilator public*/, input [7:0] I_0__1/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0(.I_0__0(I_0__0), .I_0__1(I_0__1), .O_0(NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .valid_down(NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0 = NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
assign valid_down = NativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ (input CLK/*verilator public*/, input [7:0] I0_0/*verilator public*/, input [7:0] I0_1/*verilator public*/, input [7:0] I0_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output [7:0] O_1_0/*verilator public*/, output [7:0] O_1_1/*verilator public*/, output [7:0] O_1_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
wire [7:0] Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
wire [7:0] Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2;
wire [7:0] Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_0;
wire [7:0] Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_1;
wire [7:0] Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_2;
wire Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0(I0_0), .I0_1(I0_1), .I0_2(I0_2), .I1_0(I1_0), .I1_1(I1_1), .I1_2(I1_2), .O_0_0(Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0), .O_0_1(Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1), .O_0_2(Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2), .O_1_0(Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_0), .O_1_1(Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_1), .O_1_2(Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_2), .valid_down(Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
assign O_0_1 = Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
assign O_0_2 = Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2;
assign O_1_0 = Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_0;
assign O_1_1 = Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_1;
assign O_1_2 = Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_2;
assign valid_down = Map_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
endmodule

module Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ (input CLK/*verilator public*/, input [7:0] I0_0_0/*verilator public*/, input [7:0] I0_0_1/*verilator public*/, input [7:0] I0_0_2/*verilator public*/, input [7:0] I0_1_0/*verilator public*/, input [7:0] I0_1_1/*verilator public*/, input [7:0] I0_1_2/*verilator public*/, input [7:0] I1_0/*verilator public*/, input [7:0] I1_1/*verilator public*/, input [7:0] I1_2/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output [7:0] O_1_0/*verilator public*/, output [7:0] O_1_1/*verilator public*/, output [7:0] O_1_2/*verilator public*/, output [7:0] O_2_0/*verilator public*/, output [7:0] O_2_1/*verilator public*/, output [7:0] O_2_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_0;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_1;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_2;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_0;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_1;
wire [7:0] Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_2;
wire Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0_0(I0_0_0), .I0_0_1(I0_0_1), .I0_0_2(I0_0_2), .I0_1_0(I0_1_0), .I0_1_1(I0_1_1), .I0_1_2(I0_1_2), .I1_0(I1_0), .I1_1(I1_1), .I1_2(I1_2), .O_0_0(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0), .O_0_1(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1), .O_0_2(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2), .O_1_0(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_0), .O_1_1(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_1), .O_1_2(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_2), .O_2_0(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_0), .O_2_1(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_1), .O_2_2(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_2), .valid_down(Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
assign O_0_1 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
assign O_0_2 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2;
assign O_1_0 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_0;
assign O_1_1 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_1;
assign O_1_2 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1_2;
assign O_2_0 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_0;
assign O_2_1 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_1;
assign O_2_2 = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2_2;
assign valid_down = Map_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
endmodule

module Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ (input CLK/*verilator public*/, input [7:0] I_0_0/*verilator public*/, input [7:0] I_0_1/*verilator public*/, input [7:0] I_0_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire [7:0] Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1;
wire [7:0] Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2;
wire Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0_0(I_0_0), .I_0_1(I_0_1), .I_0_2(I_0_2), .O_0(Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_1(Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1), .O_2(Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2), .valid_down(Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(valid_up));
assign O_0 = Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
assign O_1 = Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1;
assign O_2 = Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2;
assign valid_down = Map_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
endmodule

module Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ (input CLK/*verilator public*/, input [7:0] I0_0/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
wire Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0(I0_0), .I1_0(I1_0), .O_0_0(Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0), .O_0_1(Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1), .valid_down(Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
assign O_0_1 = Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
assign valid_down = Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
endmodule

module Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ (input CLK/*verilator public*/, input [7:0] I0_0_0/*verilator public*/, input [7:0] I0_0_1/*verilator public*/, input [7:0] I1_0/*verilator public*/, output [7:0] O_0_0/*verilator public*/, output [7:0] O_0_1/*verilator public*/, output [7:0] O_0_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2;
wire Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0_0(I0_0_0), .I0_0_1(I0_0_1), .I1_0(I1_0), .O_0_0(Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0), .O_0_1(Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1), .O_0_2(Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2), .valid_down(Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_0;
assign O_0_1 = Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_1;
assign O_0_2 = Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0_2;
assign valid_down = Map_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
endmodule

module LUT4_5 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, input I3/*verilator public*/, output O/*verilator public*/);
wire coreir_lut4_inst0_out;
lutN #(.init(16'h0005), .N(4)) coreir_lut4_inst0(.in({I3,I2,I1,I0}), .out(coreir_lut4_inst0_out));
assign O = coreir_lut4_inst0_out;
endmodule

module LUT4_256 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, input I3/*verilator public*/, output O/*verilator public*/);
wire coreir_lut4_inst0_out;
lutN #(.init(16'h0100), .N(4)) coreir_lut4_inst0(.in({I3,I2,I1,I0}), .out(coreir_lut4_inst0_out));
assign O = coreir_lut4_inst0_out;
endmodule

module LUT4_2048 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, input I3/*verilator public*/, output O/*verilator public*/);
wire coreir_lut4_inst0_out;
lutN #(.init(16'h0800), .N(4)) coreir_lut4_inst0(.in({I3,I2,I1,I0}), .out(coreir_lut4_inst0_out));
assign O = coreir_lut4_inst0_out;
endmodule

module LUT4_2 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, input I3/*verilator public*/, output O/*verilator public*/);
wire coreir_lut4_inst0_out;
lutN #(.init(16'h0002), .N(4)) coreir_lut4_inst0(.in({I3,I2,I1,I0}), .out(coreir_lut4_inst0_out));
assign O = coreir_lut4_inst0_out;
endmodule

module LUT4_1 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, input I3/*verilator public*/, output O/*verilator public*/);
wire coreir_lut4_inst0_out;
lutN #(.init(16'h0001), .N(4)) coreir_lut4_inst0(.in({I3,I2,I1,I0}), .out(coreir_lut4_inst0_out));
assign O = coreir_lut4_inst0_out;
endmodule

module LUT4_0 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, input I3/*verilator public*/, output O/*verilator public*/);
wire coreir_lut4_inst0_out;
lutN #(.init(16'h0000), .N(4)) coreir_lut4_inst0(.in({I3,I2,I1,I0}), .out(coreir_lut4_inst0_out));
assign O = coreir_lut4_inst0_out;
endmodule

module LUT_Array_3_Array_8_Bit__t_9n (input CLK/*verilator public*/, input [3:0] addr/*verilator public*/, output [7:0] data_0/*verilator public*/, output [7:0] data_1/*verilator public*/, output [7:0] data_2/*verilator public*/);
wire LUT4_0_inst0_O;
wire LUT4_0_inst1_O;
wire LUT4_0_inst10_O;
wire LUT4_0_inst11_O;
wire LUT4_0_inst12_O;
wire LUT4_0_inst13_O;
wire LUT4_0_inst14_O;
wire LUT4_0_inst15_O;
wire LUT4_0_inst16_O;
wire LUT4_0_inst17_O;
wire LUT4_0_inst18_O;
wire LUT4_0_inst19_O;
wire LUT4_0_inst2_O;
wire LUT4_0_inst3_O;
wire LUT4_0_inst4_O;
wire LUT4_0_inst5_O;
wire LUT4_0_inst6_O;
wire LUT4_0_inst7_O;
wire LUT4_0_inst8_O;
wire LUT4_0_inst9_O;
wire LUT4_2_inst0_O;
wire LUT4_2_inst1_O;
wire LUT4_2_inst2_O;
wire LUT4_5_inst0_O;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_0;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_1;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_2;
LUT4_0 LUT4_0_inst0(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst0_O));
LUT4_0 LUT4_0_inst1(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst1_O));
LUT4_0 LUT4_0_inst10(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst10_O));
LUT4_0 LUT4_0_inst11(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst11_O));
LUT4_0 LUT4_0_inst12(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst12_O));
LUT4_0 LUT4_0_inst13(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst13_O));
LUT4_0 LUT4_0_inst14(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst14_O));
LUT4_0 LUT4_0_inst15(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst15_O));
LUT4_0 LUT4_0_inst16(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst16_O));
LUT4_0 LUT4_0_inst17(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst17_O));
LUT4_0 LUT4_0_inst18(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst18_O));
LUT4_0 LUT4_0_inst19(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst19_O));
LUT4_0 LUT4_0_inst2(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst2_O));
LUT4_0 LUT4_0_inst3(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst3_O));
LUT4_0 LUT4_0_inst4(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst4_O));
LUT4_0 LUT4_0_inst5(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst5_O));
LUT4_0 LUT4_0_inst6(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst6_O));
LUT4_0 LUT4_0_inst7(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst7_O));
LUT4_0 LUT4_0_inst8(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst8_O));
LUT4_0 LUT4_0_inst9(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst9_O));
LUT4_2 LUT4_2_inst0(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_2_inst0_O));
LUT4_2 LUT4_2_inst1(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_2_inst1_O));
LUT4_2 LUT4_2_inst2(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_2_inst2_O));
LUT4_5 LUT4_5_inst0(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_5_inst0_O));
\aetherlinglib_hydrate__hydratedTypeBit83 hydrate_tArray_3_Array_8_Bit___inst0(.in({LUT4_0_inst19_O,LUT4_0_inst18_O,LUT4_0_inst17_O,LUT4_0_inst16_O,LUT4_0_inst15_O,LUT4_0_inst14_O,LUT4_0_inst13_O,LUT4_2_inst2_O,LUT4_0_inst12_O,LUT4_0_inst11_O,LUT4_0_inst10_O,LUT4_0_inst9_O,LUT4_0_inst8_O,LUT4_0_inst7_O,LUT4_2_inst1_O,LUT4_5_inst0_O,LUT4_0_inst6_O,LUT4_0_inst5_O,LUT4_0_inst4_O,LUT4_0_inst3_O,LUT4_0_inst2_O,LUT4_0_inst1_O,LUT4_0_inst0_O,LUT4_2_inst0_O}), .out_0(hydrate_tArray_3_Array_8_Bit___inst0_out_0), .out_1(hydrate_tArray_3_Array_8_Bit___inst0_out_1), .out_2(hydrate_tArray_3_Array_8_Bit___inst0_out_2));
assign data_0 = hydrate_tArray_3_Array_8_Bit___inst0_out_0;
assign data_1 = hydrate_tArray_3_Array_8_Bit___inst0_out_1;
assign data_2 = hydrate_tArray_3_Array_8_Bit___inst0_out_2;
endmodule

module LUT_Array_1_Array_8_Bit__t_9n (input CLK/*verilator public*/, input [3:0] addr/*verilator public*/, output [7:0] data_0/*verilator public*/);
wire LUT4_0_inst0_O;
wire LUT4_0_inst1_O;
wire LUT4_0_inst2_O;
wire LUT4_0_inst3_O;
wire LUT4_0_inst4_O;
wire LUT4_0_inst5_O;
wire LUT4_0_inst6_O;
wire LUT4_1_inst0_O;
wire [7:0] hydrate_tArray_1_Array_8_Bit___inst0_out_0;
LUT4_0 LUT4_0_inst0(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst0_O));
LUT4_0 LUT4_0_inst1(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst1_O));
LUT4_0 LUT4_0_inst2(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst2_O));
LUT4_0 LUT4_0_inst3(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst3_O));
LUT4_0 LUT4_0_inst4(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst4_O));
LUT4_0 LUT4_0_inst5(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst5_O));
LUT4_0 LUT4_0_inst6(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_0_inst6_O));
LUT4_1 LUT4_1_inst0(.I0(addr[0]), .I1(addr[1]), .I2(addr[2]), .I3(addr[3]), .O(LUT4_1_inst0_O));
\aetherlinglib_hydrate__hydratedTypeBit81 hydrate_tArray_1_Array_8_Bit___inst0(.in({LUT4_0_inst6_O,LUT4_0_inst5_O,LUT4_0_inst4_O,LUT4_0_inst3_O,LUT4_0_inst2_O,LUT4_1_inst0_O,LUT4_0_inst1_O,LUT4_0_inst0_O}), .out_0(hydrate_tArray_1_Array_8_Bit___inst0_out_0));
assign data_0 = hydrate_tArray_1_Array_8_Bit___inst0_out_0;
endmodule

module LUT3_64 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, output O/*verilator public*/);
wire coreir_lut3_inst0_out;
lutN #(.init(8'h40), .N(3)) coreir_lut3_inst0(.in({I2,I1,I0}), .out(coreir_lut3_inst0_out));
assign O = coreir_lut3_inst0_out;
endmodule

module LUT3_128 (input I0/*verilator public*/, input I1/*verilator public*/, input I2/*verilator public*/, output O/*verilator public*/);
wire coreir_lut3_inst0_out;
lutN #(.init(8'h80), .N(3)) coreir_lut3_inst0(.in({I2,I1,I0}), .out(coreir_lut3_inst0_out));
assign O = coreir_lut3_inst0_out;
endmodule

module LUT2_8 (input I0/*verilator public*/, input I1/*verilator public*/, output O/*verilator public*/);
wire coreir_lut2_inst0_out;
lutN #(.init(4'h8), .N(2)) coreir_lut2_inst0(.in({I1,I0}), .out(coreir_lut2_inst0_out));
assign O = coreir_lut2_inst0_out;
endmodule

module LUT2_4 (input I0/*verilator public*/, input I1/*verilator public*/, output O/*verilator public*/);
wire coreir_lut2_inst0_out;
lutN #(.init(4'h4), .N(2)) coreir_lut2_inst0(.in({I1,I0}), .out(coreir_lut2_inst0_out));
assign O = coreir_lut2_inst0_out;
endmodule

module LUT2_2 (input I0/*verilator public*/, input I1/*verilator public*/, output O/*verilator public*/);
wire coreir_lut2_inst0_out;
lutN #(.init(4'h2), .N(2)) coreir_lut2_inst0(.in({I1,I0}), .out(coreir_lut2_inst0_out));
assign O = coreir_lut2_inst0_out;
endmodule

module LUT2_1 (input I0/*verilator public*/, input I1/*verilator public*/, output O/*verilator public*/);
wire coreir_lut2_inst0_out;
lutN #(.init(4'h1), .N(2)) coreir_lut2_inst0(.in({I1,I0}), .out(coreir_lut2_inst0_out));
assign O = coreir_lut2_inst0_out;
endmodule

module LUT1_1 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h1), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LShift_Atom (input [7:0] I__0/*verilator public*/, input [7:0] I__1/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] shl8_inst0_out;
coreir_shl #(.width(8)) shl8_inst0(.in0(I__0), .in1(I__1), .out(shl8_inst0_out));
assign O = shl8_inst0_out;
assign valid_down = valid_up;
endmodule

module NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit__ (input [7:0] I_0__0/*verilator public*/, input [7:0] I_0__1/*verilator public*/, input [7:0] I_1__0/*verilator public*/, input [7:0] I_1__1/*verilator public*/, input [7:0] I_2__0/*verilator public*/, input [7:0] I_2__1/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] LShift_Atom_inst0_O;
wire LShift_Atom_inst0_valid_down;
wire [7:0] LShift_Atom_inst1_O;
wire LShift_Atom_inst1_valid_down;
wire [7:0] LShift_Atom_inst2_O;
wire LShift_Atom_inst2_valid_down;
wire and_inst0_out;
wire and_inst1_out;
LShift_Atom LShift_Atom_inst0(.I__0(I_0__0), .I__1(I_0__1), .O(LShift_Atom_inst0_O), .valid_down(LShift_Atom_inst0_valid_down), .valid_up(valid_up));
LShift_Atom LShift_Atom_inst1(.I__0(I_1__0), .I__1(I_1__1), .O(LShift_Atom_inst1_O), .valid_down(LShift_Atom_inst1_valid_down), .valid_up(valid_up));
LShift_Atom LShift_Atom_inst2(.I__0(I_2__0), .I__1(I_2__1), .O(LShift_Atom_inst2_O), .valid_down(LShift_Atom_inst2_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(LShift_Atom_inst0_valid_down), .in1(LShift_Atom_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(LShift_Atom_inst2_valid_down), .out(and_inst1_out));
assign O_0 = LShift_Atom_inst0_O;
assign O_1 = LShift_Atom_inst1_O;
assign O_2 = LShift_Atom_inst2_O;
assign valid_down = and_inst1_out;
endmodule

module Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I_0__0/*verilator public*/, input [7:0] I_0__1/*verilator public*/, input [7:0] I_1__0/*verilator public*/, input [7:0] I_1__1/*verilator public*/, input [7:0] I_2__0/*verilator public*/, input [7:0] I_2__1/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0(.I_0__0(I_0__0), .I_0__1(I_0__1), .I_1__0(I_1__0), .I_1__1(I_1__1), .I_2__0(I_2__0), .I_2__1(I_2__1), .O_0(NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_2(NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .valid_down(NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0 = NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
assign O_1 = NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
assign O_2 = NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
assign valid_down = NativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire Mux2xNone_inst0_O;
wire [0:0] reg_P_inst0_out;
Mux2xNone Mux2xNone_inst0(.I0(reg_P_inst0_out[0]), .I1(I), .O(Mux2xNone_inst0_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(Mux2xNone_inst0_O), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Register8CE (input CE/*verilator public*/, input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7_O;
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0(.CE(CE), .CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1(.CE(CE), .CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2(.CE(CE), .CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3(.CE(CE), .CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4(.CE(CE), .CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5(.CE(CE), .CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6(.CE(CE), .CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7(.CE(CE), .CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7_O));
assign O = {DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_8_Out_Bit__t_0init_TrueCE_FalseRESET (input CE/*verilator public*/, input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] Register8CE_inst0_O;
Register8CE Register8CE_inst0(.CE(CE), .CLK(CLK), .I(I), .O(Register8CE_inst0_O));
assign O = Register8CE_inst0_O;
endmodule

module Register_Array_1_Array_8_Out_Bit___t_0init_TrueCE_FalseRESET (input CE/*verilator public*/, input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] O_0/*verilator public*/);
wire [7:0] Register_Array_8_Out_Bit__t_0init_TrueCE_FalseRESET_inst0_O;
Register_Array_8_Out_Bit__t_0init_TrueCE_FalseRESET Register_Array_8_Out_Bit__t_0init_TrueCE_FalseRESET_inst0(.CE(CE), .CLK(CLK), .I(I_0), .O(Register_Array_8_Out_Bit__t_0init_TrueCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_8_Out_Bit__t_0init_TrueCE_FalseRESET_inst0_O;
endmodule

module Register_Array_8_Bit_t_0init_TrueCE_FalseRESET (input CE/*verilator public*/, input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] Register8CE_inst0_O;
Register8CE Register8CE_inst0(.CE(CE), .CLK(CLK), .I(I), .O(Register8CE_inst0_O));
assign O = Register8CE_inst0_O;
endmodule

module Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET (input CE/*verilator public*/, input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/);
wire [7:0] Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0_O;
wire [7:0] Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst1_O;
wire [7:0] Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst2_O;
Register_Array_8_Bit_t_0init_TrueCE_FalseRESET Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0(.CE(CE), .CLK(CLK), .I(I_0), .O(Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0_O));
Register_Array_8_Bit_t_0init_TrueCE_FalseRESET Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst1(.CE(CE), .CLK(CLK), .I(I_1), .O(Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst1_O));
Register_Array_8_Bit_t_0init_TrueCE_FalseRESET Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst2(.CE(CE), .CLK(CLK), .I(I_2), .O(Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst2_O));
assign O_0 = Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0_O;
assign O_1 = Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst1_O;
assign O_2 = Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst2_O;
endmodule

module DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Register8 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_8_Bit_t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] Register8_inst0_O;
Register8 Register8_inst0(.CLK(CLK), .I(I), .O(Register8_inst0_O));
assign O = Register8_inst0_O;
endmodule

module Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/);
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O;
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(I_0), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1(.CLK(CLK), .I(I_1), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2(.CLK(CLK), .I(I_2), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O));
assign O_0 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
assign O_1 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O;
assign O_2 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O;
endmodule

module Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] O_0/*verilator public*/);
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(I_0), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Register1 (input CLK/*verilator public*/, input [0:0] I/*verilator public*/, output [0:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
assign O = DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
endmodule

module Register_Bitt_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] Register1_inst0_O;
Register1 Register1_inst0(.CLK(CLK), .I(I), .O(Register1_inst0_O));
assign O = Register1_inst0_O[0];
endmodule

module FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(I_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Counter4CER (input CE/*verilator public*/, input CLK/*verilator public*/, output [3:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [3:0] Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_4_inst0_O;
wire [3:0] const_1_4_out;
wire [3:0] coreir_add4_inst0_out;
Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_4 Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_4_inst0(.CE(CE), .CLK(CLK), .I(coreir_add4_inst0_out), .O(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_4_inst0_O), .RESET(RESET));
coreir_const #(.value(4'h1), .width(4)) const_1_4(.out(const_1_4_out));
coreir_add #(.width(4)) coreir_add4_inst0(.in0(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_4_inst0_O), .in1(const_1_4_out), .out(coreir_add4_inst0_out));
assign O = Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_4_inst0_O;
endmodule

module Counter4_Mod9CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [3:0] O/*verilator public*/);
wire [3:0] Counter4CER_inst0_O;
wire LUT4_256_inst0_O;
wire and_inst0_out;
Counter4CER Counter4CER_inst0(.CE(CE), .CLK(CLK), .O(Counter4CER_inst0_O), .RESET(and_inst0_out));
LUT4_256 LUT4_256_inst0(.I0(Counter4CER_inst0_O[0]), .I1(Counter4CER_inst0_O[1]), .I2(Counter4CER_inst0_O[2]), .I3(Counter4CER_inst0_O[3]), .O(LUT4_256_inst0_O));
corebit_and and_inst0(.in0(LUT4_256_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter4CER_inst0_O;
endmodule

module serialize_tSSeq_3_Int__n3_i6_hasRESETFalse (input CLK/*verilator public*/, input [7:0] I_0_0/*verilator public*/, input [7:0] I_0_1/*verilator public*/, input [7:0] I_0_2/*verilator public*/, input [7:0] I_1_0/*verilator public*/, input [7:0] I_1_1/*verilator public*/, input [7:0] I_1_2/*verilator public*/, input [7:0] I_2_0/*verilator public*/, input [7:0] I_2_1/*verilator public*/, input [7:0] I_2_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire LUT2_1_inst0_O;
wire [7:0] Mux_Array_3_Array_8_Bit__t_2n_inst0_out_0;
wire [7:0] Mux_Array_3_Array_8_Bit__t_2n_inst0_out_1;
wire [7:0] Mux_Array_3_Array_8_Bit__t_2n_inst0_out_2;
wire [7:0] Mux_Array_3_Array_8_Bit__t_3n_inst0_out_0;
wire [7:0] Mux_Array_3_Array_8_Bit__t_3n_inst0_out_1;
wire [7:0] Mux_Array_3_Array_8_Bit__t_3n_inst0_out_2;
wire [0:0] Register1_inst0_O;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_1;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_2;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_0;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_1;
wire [7:0] Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_2;
wire and_inst0_out;
wire and_inst1_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(valid_up), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
LUT2_1 LUT2_1_inst0(.I0(Counter4_Mod9CE_inst0_O[0]), .I1(Counter4_Mod9CE_inst0_O[1]), .O(LUT2_1_inst0_O));
Mux_Array_3_Array_8_Bit__t_2n Mux_Array_3_Array_8_Bit__t_2n_inst0(.data_0_0(Mux_Array_3_Array_8_Bit__t_3n_inst0_out_0), .data_0_1(Mux_Array_3_Array_8_Bit__t_3n_inst0_out_1), .data_0_2(Mux_Array_3_Array_8_Bit__t_3n_inst0_out_2), .data_1_0(I_0_0), .data_1_1(I_0_1), .data_1_2(I_0_2), .out_0(Mux_Array_3_Array_8_Bit__t_2n_inst0_out_0), .out_1(Mux_Array_3_Array_8_Bit__t_2n_inst0_out_1), .out_2(Mux_Array_3_Array_8_Bit__t_2n_inst0_out_2), .sel(LUT2_1_inst0_O));
Mux_Array_3_Array_8_Bit__t_3n Mux_Array_3_Array_8_Bit__t_3n_inst0(.data_0_0(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_0), .data_0_1(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_1), .data_0_2(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_2), .data_1_0(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_0), .data_1_1(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_1), .data_1_2(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_2), .data_2_0(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_0), .data_2_1(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_1), .data_2_2(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_2), .out_0(Mux_Array_3_Array_8_Bit__t_3n_inst0_out_0), .out_1(Mux_Array_3_Array_8_Bit__t_3n_inst0_out_1), .out_2(Mux_Array_3_Array_8_Bit__t_3n_inst0_out_2), .sel({Counter4_Mod9CE_inst0_O[1],Counter4_Mod9CE_inst0_O[0]}));
Register1 Register1_inst0(.CLK(CLK), .I(valid_up), .O(Register1_inst0_O));
Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(Mux_Array_3_Array_8_Bit__t_2n_inst0_out_0), .I_1(Mux_Array_3_Array_8_Bit__t_2n_inst0_out_1), .I_2(Mux_Array_3_Array_8_Bit__t_2n_inst0_out_2), .O_0(Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0), .O_1(Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1), .O_2(Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2));
Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0(.CE(and_inst0_out), .CLK(CLK), .I_0(I_1_0), .I_1(I_1_1), .I_2(I_1_2), .O_0(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_0), .O_1(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_1), .O_2(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst0_O_2));
Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1(.CE(and_inst1_out), .CLK(CLK), .I_0(I_2_0), .I_1(I_2_1), .I_2(I_2_2), .O_0(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_0), .O_1(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_1), .O_2(Register_Array_3_Array_8_Bit__t_0init_TrueCE_FalseRESET_inst1_O_2));
Term_Array_2_Bit_t Term_Array_2_Bit_t_inst0(.I({Counter4_Mod9CE_inst0_O[3],Counter4_Mod9CE_inst0_O[2]}));
corebit_and and_inst0(.in0(LUT2_1_inst0_O), .in1(valid_up), .out(and_inst0_out));
corebit_and and_inst1(.in0(LUT2_1_inst0_O), .in1(valid_up), .out(and_inst1_out));
assign O_0 = Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign O_1 = Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
assign O_2 = Register_Array_3_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
assign valid_down = Register1_inst0_O[0];
endmodule

module Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I_0_0/*verilator public*/, input [7:0] I_0_1/*verilator public*/, input [7:0] I_0_2/*verilator public*/, input [7:0] I_1_0/*verilator public*/, input [7:0] I_1_1/*verilator public*/, input [7:0] I_1_2/*verilator public*/, input [7:0] I_2_0/*verilator public*/, input [7:0] I_2_1/*verilator public*/, input [7:0] I_2_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_0;
wire [7:0] serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_1;
wire [7:0] serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_2;
wire serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_valid_down;
serialize_tSSeq_3_Int__n3_i6_hasRESETFalse serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0(.CLK(CLK), .I_0_0(I_0_0), .I_0_1(I_0_1), .I_0_2(I_0_2), .I_1_0(I_1_0), .I_1_1(I_1_1), .I_1_2(I_1_2), .I_2_0(I_2_0), .I_2_1(I_2_1), .I_2_2(I_2_2), .O_0(serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_0), .O_1(serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_1), .O_2(serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_2), .valid_down(serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_valid_down), .valid_up(valid_up));
assign O_0 = serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_0;
assign O_1 = serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_1;
assign O_2 = serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_O_2;
assign valid_down = serialize_tSSeq_3_Int__n3_i6_hasRESETFalse_inst0_valid_down;
endmodule

module NestedCounters_TSeq_3_6_SSeq_1_Int___hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid;
wire and_inst0_out;
wire and_inst1_out;
wire [3:0] coreir_const43_inst0_out;
wire coreir_ult4_inst0_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(and_inst1_out), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0(.CE(CE), .CLK(CLK), .last(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid));
corebit_and and_inst0(.in0(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid), .in1(coreir_ult4_inst0_out), .out(and_inst0_out));
corebit_and and_inst1(.in0(CE), .in1(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .out(and_inst1_out));
coreir_const #(.value(4'h3), .width(4)) coreir_const43_inst0(.out(coreir_const43_inst0_out));
coreir_ult #(.width(4)) coreir_ult4_inst0(.in0(Counter4_Mod9CE_inst0_O), .in1(coreir_const43_inst0_out), .out(coreir_ult4_inst0_out));
assign valid = and_inst0_out;
endmodule

module NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_unq1 (input CE/*verilator public*/, input CLK/*verilator public*/, output last/*verilator public*/, output valid/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire LUT4_256_inst0_O;
wire NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire [3:0] coreir_const41_inst0_out;
wire coreir_ult4_inst0_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(and_inst2_out), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
LUT4_256 LUT4_256_inst0(.I0(Counter4_Mod9CE_inst0_O[0]), .I1(Counter4_Mod9CE_inst0_O[1]), .I2(Counter4_Mod9CE_inst0_O[2]), .I3(Counter4_Mod9CE_inst0_O[3]), .O(LUT4_256_inst0_O));
NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0(.CE(CE), .CLK(CLK), .last(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid));
corebit_and and_inst0(.in0(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid), .in1(coreir_ult4_inst0_out), .out(and_inst0_out));
corebit_and and_inst1(.in0(LUT4_256_inst0_O), .in1(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .out(and_inst1_out));
corebit_and and_inst2(.in0(CE), .in1(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .out(and_inst2_out));
coreir_const #(.value(4'h1), .width(4)) coreir_const41_inst0(.out(coreir_const41_inst0_out));
coreir_ult #(.width(4)) coreir_ult4_inst0(.in0(Counter4_Mod9CE_inst0_O), .in1(coreir_const41_inst0_out), .out(coreir_ult4_inst0_out));
assign last = and_inst1_out;
assign valid = and_inst0_out;
endmodule

module NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] cur_valid/*verilator public*/, output last/*verilator public*/, output valid/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire LUT4_256_inst0_O;
wire NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire [3:0] coreir_const41_inst0_out;
wire coreir_ult4_inst0_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(and_inst2_out), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
LUT4_256 LUT4_256_inst0(.I0(Counter4_Mod9CE_inst0_O[0]), .I1(Counter4_Mod9CE_inst0_O[1]), .I2(Counter4_Mod9CE_inst0_O[2]), .I3(Counter4_Mod9CE_inst0_O[3]), .O(LUT4_256_inst0_O));
NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0(.CE(CE), .CLK(CLK), .last(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(and_inst4_out), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
corebit_and and_inst0(.in0(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid), .in1(coreir_ult4_inst0_out), .out(and_inst0_out));
corebit_and and_inst1(.in0(LUT4_256_inst0_O), .in1(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .out(and_inst1_out));
corebit_and and_inst2(.in0(CE), .in1(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_last), .out(and_inst2_out));
corebit_and and_inst3(.in0(CE), .in1(NestedCounters_SSeq_1_Int__hasCETrue_hasResetFalse_inst0_valid), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(coreir_ult4_inst0_out), .out(and_inst4_out));
coreir_const #(.value(4'h1), .width(4)) coreir_const41_inst0(.out(coreir_const41_inst0_out));
coreir_ult #(.width(4)) coreir_ult4_inst0(.in0(Counter4_Mod9CE_inst0_O), .in1(coreir_const41_inst0_out), .out(coreir_ult4_inst0_out));
assign cur_valid = SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
assign last = and_inst1_out;
assign valid = and_inst0_out;
endmodule

module RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_unq1 (input CLK/*verilator public*/, input [0:0] RADDR/*verilator public*/, output [7:0] RDATA_0/*verilator public*/, input RE/*verilator public*/, input [0:0] WADDR/*verilator public*/, input [7:0] WDATA_0/*verilator public*/, input WE/*verilator public*/);
wire LUT1_1_inst0_O;
wire [7:0] Mux_Array_1_Array_8_Bit__t_1n_inst0_out_0;
wire [0:0] NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid;
wire [0:0] NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_last;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid;
wire [7:0] RAM_Array_1_Array_8_Bit__t_1n_inst0_RDATA_0;
wire and_inst0_out;
LUT1_1 LUT1_1_inst0(.I0(WADDR[0]), .O(LUT1_1_inst0_O));
Mux_Array_1_Array_8_Bit__t_1n Mux_Array_1_Array_8_Bit__t_1n_inst0(.data_0_0(RAM_Array_1_Array_8_Bit__t_1n_inst0_RDATA_0), .out_0(Mux_Array_1_Array_8_Bit__t_1n_inst0_out_0), .sel(RADDR));
NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0(.CE(RE), .CLK(CLK), .cur_valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid), .last(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1(.CE(WE), .CLK(CLK), .cur_valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid), .last(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_last), .valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid));
RAM_Array_1_Array_8_Bit__t_1n RAM_Array_1_Array_8_Bit__t_1n_inst0(.CLK(CLK), .RADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid), .RDATA_0(RAM_Array_1_Array_8_Bit__t_1n_inst0_RDATA_0), .WADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid), .WDATA_0(WDATA_0), .WE(and_inst0_out));
Term_Bitt Term_Bitt_inst0(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
Term_Bitt Term_Bitt_inst1(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last));
Term_Bitt Term_Bitt_inst2(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid));
Term_Bitt Term_Bitt_inst3(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_last));
corebit_and and_inst0(.in0(LUT1_1_inst0_O), .in1(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid), .out(and_inst0_out));
assign RDATA_0 = Mux_Array_1_Array_8_Bit__t_1n_inst0_out_0;
endmodule

module Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid;
wire [7:0] RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0_RDATA_0;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire and_inst0_out;
wire and_inst1_out;
wire [0:0] coreir_const11_inst0_out;
NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_unq1 NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0(.CE(and_inst0_out), .CLK(CLK), .last(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_unq1 RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0(.CLK(CLK), .RADDR(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .RDATA_0(RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0_RDATA_0), .RE(and_inst0_out), .WADDR(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .WDATA_0(I_0), .WE(and_inst0_out));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(and_inst1_out), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
corebit_and and_inst0(.in0(valid_up), .in1(coreir_const11_inst0_out[0]), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last), .out(and_inst1_out));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0_RDATA_0;
assign valid_down = valid_up;
endmodule

module RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse (input CLK/*verilator public*/, input [1:0] RADDR/*verilator public*/, output [7:0] RDATA_0/*verilator public*/, input RE/*verilator public*/, input [1:0] WADDR/*verilator public*/, input [7:0] WDATA_0/*verilator public*/, input WE/*verilator public*/);
wire LUT2_1_inst0_O;
wire LUT2_2_inst0_O;
wire LUT2_4_inst0_O;
wire LUT2_8_inst0_O;
wire [7:0] Mux_Array_1_Array_8_Bit__t_4n_inst0_out_0;
wire [0:0] NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid;
wire [0:0] NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_last;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid;
wire [7:0] RAM_Array_1_Array_8_Bit__t_1n_inst0_RDATA_0;
wire [7:0] RAM_Array_1_Array_8_Bit__t_1n_inst1_RDATA_0;
wire [7:0] RAM_Array_1_Array_8_Bit__t_1n_inst2_RDATA_0;
wire [7:0] RAM_Array_1_Array_8_Bit__t_1n_inst3_RDATA_0;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
LUT2_1 LUT2_1_inst0(.I0(WADDR[0]), .I1(WADDR[1]), .O(LUT2_1_inst0_O));
LUT2_2 LUT2_2_inst0(.I0(WADDR[0]), .I1(WADDR[1]), .O(LUT2_2_inst0_O));
LUT2_4 LUT2_4_inst0(.I0(WADDR[0]), .I1(WADDR[1]), .O(LUT2_4_inst0_O));
LUT2_8 LUT2_8_inst0(.I0(WADDR[0]), .I1(WADDR[1]), .O(LUT2_8_inst0_O));
Mux_Array_1_Array_8_Bit__t_4n Mux_Array_1_Array_8_Bit__t_4n_inst0(.data_0_0(RAM_Array_1_Array_8_Bit__t_1n_inst0_RDATA_0), .data_1_0(RAM_Array_1_Array_8_Bit__t_1n_inst1_RDATA_0), .data_2_0(RAM_Array_1_Array_8_Bit__t_1n_inst2_RDATA_0), .data_3_0(RAM_Array_1_Array_8_Bit__t_1n_inst3_RDATA_0), .out_0(Mux_Array_1_Array_8_Bit__t_4n_inst0_out_0), .sel(RADDR));
NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0(.CE(RE), .CLK(CLK), .cur_valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid), .last(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1(.CE(WE), .CLK(CLK), .cur_valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid), .last(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_last), .valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid));
RAM_Array_1_Array_8_Bit__t_1n RAM_Array_1_Array_8_Bit__t_1n_inst0(.CLK(CLK), .RADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid), .RDATA_0(RAM_Array_1_Array_8_Bit__t_1n_inst0_RDATA_0), .WADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid), .WDATA_0(WDATA_0), .WE(and_inst0_out));
RAM_Array_1_Array_8_Bit__t_1n RAM_Array_1_Array_8_Bit__t_1n_inst1(.CLK(CLK), .RADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid), .RDATA_0(RAM_Array_1_Array_8_Bit__t_1n_inst1_RDATA_0), .WADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid), .WDATA_0(WDATA_0), .WE(and_inst1_out));
RAM_Array_1_Array_8_Bit__t_1n RAM_Array_1_Array_8_Bit__t_1n_inst2(.CLK(CLK), .RADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid), .RDATA_0(RAM_Array_1_Array_8_Bit__t_1n_inst2_RDATA_0), .WADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid), .WDATA_0(WDATA_0), .WE(and_inst2_out));
RAM_Array_1_Array_8_Bit__t_1n RAM_Array_1_Array_8_Bit__t_1n_inst3(.CLK(CLK), .RADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_cur_valid), .RDATA_0(RAM_Array_1_Array_8_Bit__t_1n_inst3_RDATA_0), .WADDR(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_cur_valid), .WDATA_0(WDATA_0), .WE(and_inst3_out));
Term_Bitt Term_Bitt_inst0(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
Term_Bitt Term_Bitt_inst1(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last));
Term_Bitt Term_Bitt_inst2(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid));
Term_Bitt Term_Bitt_inst3(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_last));
corebit_and and_inst0(.in0(LUT2_1_inst0_O), .in1(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid), .out(and_inst0_out));
corebit_and and_inst1(.in0(LUT2_2_inst0_O), .in1(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid), .out(and_inst1_out));
corebit_and and_inst2(.in0(LUT2_4_inst0_O), .in1(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid), .out(and_inst2_out));
corebit_and and_inst3(.in0(LUT2_8_inst0_O), .in1(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst1_valid), .out(and_inst3_out));
assign RDATA_0 = Mux_Array_1_Array_8_Bit__t_4n_inst0_out_0;
endmodule

module Counter4_Mod12CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [3:0] O/*verilator public*/);
wire [3:0] Counter4CER_inst0_O;
wire LUT4_2048_inst0_O;
wire and_inst0_out;
Counter4CER Counter4CER_inst0(.CE(CE), .CLK(CLK), .O(Counter4CER_inst0_O), .RESET(and_inst0_out));
LUT4_2048 LUT4_2048_inst0(.I0(Counter4CER_inst0_O[0]), .I1(Counter4CER_inst0_O[1]), .I2(Counter4CER_inst0_O[2]), .I3(Counter4CER_inst0_O[3]), .O(LUT4_2048_inst0_O));
corebit_and and_inst0(.in0(LUT4_2048_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter4CER_inst0_O;
endmodule

module InitialDelayCounter_11 (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [3:0] Counter4_Mod12CE_inst0_O;
wire and_inst0_out;
wire [3:0] coreir_const411_inst0_out;
wire coreir_eq_4_inst0_out;
wire coreir_ult4_inst0_out;
Counter4_Mod12CE Counter4_Mod12CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter4_Mod12CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult4_inst0_out), .out(and_inst0_out));
coreir_const #(.value(4'hb), .width(4)) coreir_const411_inst0(.out(coreir_const411_inst0_out));
coreir_eq #(.width(4)) coreir_eq_4_inst0(.in0(Counter4_Mod12CE_inst0_O), .in1(coreir_const411_inst0_out), .out(coreir_eq_4_inst0_out));
coreir_ult #(.width(4)) coreir_ult4_inst0(.in0(Counter4_Mod12CE_inst0_O), .in1(coreir_const411_inst0_out), .out(coreir_ult4_inst0_out));
assign valid = coreir_eq_4_inst0_out;
endmodule

module Counter3CER (input CE/*verilator public*/, input CLK/*verilator public*/, output [2:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [2:0] Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0_O;
wire [2:0] const_1_3_out;
wire [2:0] coreir_add3_inst0_out;
Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3 Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0(.CE(CE), .CLK(CLK), .I(coreir_add3_inst0_out), .O(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0_O), .RESET(RESET));
coreir_const #(.value(3'h1), .width(3)) const_1_3(.out(const_1_3_out));
coreir_add #(.width(3)) coreir_add3_inst0(.in0(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0_O), .in1(const_1_3_out), .out(coreir_add3_inst0_out));
assign O = Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0_O;
endmodule

module Counter3_Mod8CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [2:0] O/*verilator public*/);
wire [2:0] Counter3CER_inst0_O;
wire LUT3_128_inst0_O;
wire and_inst0_out;
Counter3CER Counter3CER_inst0(.CE(CE), .CLK(CLK), .O(Counter3CER_inst0_O), .RESET(and_inst0_out));
LUT3_128 LUT3_128_inst0(.I0(Counter3CER_inst0_O[0]), .I1(Counter3CER_inst0_O[1]), .I2(Counter3CER_inst0_O[2]), .O(LUT3_128_inst0_O));
corebit_and and_inst0(.in0(LUT3_128_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter3CER_inst0_O;
endmodule

module InitialDelayCounter_7 (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [2:0] Counter3_Mod8CE_inst0_O;
wire and_inst0_out;
wire [2:0] coreir_const37_inst0_out;
wire coreir_eq_3_inst0_out;
wire coreir_ult3_inst0_out;
Counter3_Mod8CE Counter3_Mod8CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter3_Mod8CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult3_inst0_out), .out(and_inst0_out));
coreir_const #(.value(3'h7), .width(3)) coreir_const37_inst0(.out(coreir_const37_inst0_out));
coreir_eq #(.width(3)) coreir_eq_3_inst0(.in0(Counter3_Mod8CE_inst0_O), .in1(coreir_const37_inst0_out), .out(coreir_eq_3_inst0_out));
coreir_ult #(.width(3)) coreir_ult3_inst0(.in0(Counter3_Mod8CE_inst0_O), .in1(coreir_const37_inst0_out), .out(coreir_ult3_inst0_out));
assign valid = coreir_eq_3_inst0_out;
endmodule

module Counter3_Mod7CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [2:0] O/*verilator public*/);
wire [2:0] Counter3CER_inst0_O;
wire LUT3_64_inst0_O;
wire and_inst0_out;
Counter3CER Counter3CER_inst0(.CE(CE), .CLK(CLK), .O(Counter3CER_inst0_O), .RESET(and_inst0_out));
LUT3_64 LUT3_64_inst0(.I0(Counter3CER_inst0_O[0]), .I1(Counter3CER_inst0_O[1]), .I2(Counter3CER_inst0_O[2]), .O(LUT3_64_inst0_O));
corebit_and and_inst0(.in0(LUT3_64_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter3CER_inst0_O;
endmodule

module InitialDelayCounter_6 (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [2:0] Counter3_Mod7CE_inst0_O;
wire and_inst0_out;
wire [2:0] coreir_const36_inst0_out;
wire coreir_eq_3_inst0_out;
wire coreir_ult3_inst0_out;
Counter3_Mod7CE Counter3_Mod7CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter3_Mod7CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult3_inst0_out), .out(and_inst0_out));
coreir_const #(.value(3'h6), .width(3)) coreir_const36_inst0(.out(coreir_const36_inst0_out));
coreir_eq #(.width(3)) coreir_eq_3_inst0(.in0(Counter3_Mod7CE_inst0_O), .in1(coreir_const36_inst0_out), .out(coreir_eq_3_inst0_out));
coreir_ult #(.width(3)) coreir_ult3_inst0(.in0(Counter3_Mod7CE_inst0_O), .in1(coreir_const36_inst0_out), .out(coreir_ult3_inst0_out));
assign valid = coreir_eq_3_inst0_out;
endmodule

module Counter2CER (input CE/*verilator public*/, input CLK/*verilator public*/, output [1:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [1:0] Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O;
wire [1:0] const_1_2_out;
wire [1:0] coreir_add2_inst0_out;
Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2 Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0(.CE(CE), .CLK(CLK), .I(coreir_add2_inst0_out), .O(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O), .RESET(RESET));
coreir_const #(.value(2'h1), .width(2)) const_1_2(.out(const_1_2_out));
coreir_add #(.width(2)) coreir_add2_inst0(.in0(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O), .in1(const_1_2_out), .out(coreir_add2_inst0_out));
assign O = Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O;
endmodule

module Counter2_Mod4CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [1:0] O/*verilator public*/);
wire [1:0] Counter2CER_inst0_O;
wire LUT2_8_inst0_O;
wire and_inst0_out;
Counter2CER Counter2CER_inst0(.CE(CE), .CLK(CLK), .O(Counter2CER_inst0_O), .RESET(and_inst0_out));
LUT2_8 LUT2_8_inst0(.I0(Counter2CER_inst0_O[0]), .I1(Counter2CER_inst0_O[1]), .O(LUT2_8_inst0_O));
corebit_and and_inst0(.in0(LUT2_8_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter2CER_inst0_O;
endmodule

module Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [1:0] Counter2_Mod4CE_inst0_O;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last;
wire NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid;
wire [7:0] RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0_RDATA_0;
wire and_inst0_out;
wire and_inst1_out;
wire [0:0] coreir_const11_inst0_out;
Counter2_Mod4CE Counter2_Mod4CE_inst0(.CE(and_inst1_out), .CLK(CLK), .O(Counter2_Mod4CE_inst0_O));
NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_unq1 NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0(.CE(and_inst0_out), .CLK(CLK), .last(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last), .valid(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0(.CLK(CLK), .RADDR(Counter2_Mod4CE_inst0_O), .RDATA_0(RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0_RDATA_0), .RE(and_inst0_out), .WADDR(Counter2_Mod4CE_inst0_O), .WDATA_0(I_0), .WE(and_inst0_out));
Term_Bitt Term_Bitt_inst0(.I(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
corebit_and and_inst0(.in0(valid_up), .in1(coreir_const11_inst0_out[0]), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(NestedCounters_TSeq_1_8_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_last), .out(and_inst1_out));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = RAM_ST_TSeq_1_8_SSeq_1_Int___hasResetFalse_inst0_RDATA_0;
assign valid_down = valid_up;
endmodule

module InitialDelayCounter_3 (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [1:0] Counter2_Mod4CE_inst0_O;
wire and_inst0_out;
wire [1:0] coreir_const23_inst0_out;
wire coreir_eq_2_inst0_out;
wire coreir_ult2_inst0_out;
Counter2_Mod4CE Counter2_Mod4CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter2_Mod4CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult2_inst0_out), .out(and_inst0_out));
coreir_const #(.value(2'h3), .width(2)) coreir_const23_inst0(.out(coreir_const23_inst0_out));
coreir_eq #(.width(2)) coreir_eq_2_inst0(.in0(Counter2_Mod4CE_inst0_O), .in1(coreir_const23_inst0_out), .out(coreir_eq_2_inst0_out));
coreir_ult #(.width(2)) coreir_ult2_inst0(.in0(Counter2_Mod4CE_inst0_O), .in1(coreir_const23_inst0_out), .out(coreir_ult2_inst0_out));
assign valid = coreir_eq_2_inst0_out;
endmodule

module Counter2_Mod3CE_COUT (input CE/*verilator public*/, input CLK/*verilator public*/, output COUT/*verilator public*/, output [1:0] O/*verilator public*/);
wire [1:0] Counter2CER_inst0_O;
wire LUT2_4_inst0_O;
wire and_inst0_out;
Counter2CER Counter2CER_inst0(.CE(CE), .CLK(CLK), .O(Counter2CER_inst0_O), .RESET(and_inst0_out));
LUT2_4 LUT2_4_inst0(.I0(Counter2CER_inst0_O[0]), .I1(Counter2CER_inst0_O[1]), .O(LUT2_4_inst0_O));
corebit_and and_inst0(.in0(LUT2_4_inst0_O), .in1(CE), .out(and_inst0_out));
assign COUT = and_inst0_out;
assign O = Counter2CER_inst0_O;
endmodule

module Counter2_Mod3CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [1:0] O/*verilator public*/);
wire [1:0] Counter2CER_inst0_O;
wire LUT2_4_inst0_O;
wire and_inst0_out;
Counter2CER Counter2CER_inst0(.CE(CE), .CLK(CLK), .O(Counter2CER_inst0_O), .RESET(and_inst0_out));
LUT2_4 LUT2_4_inst0(.I0(Counter2CER_inst0_O[0]), .I1(Counter2CER_inst0_O[1]), .O(LUT2_4_inst0_O));
corebit_and and_inst0(.in0(LUT2_4_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter2CER_inst0_O;
endmodule

module InitialDelayCounter_2 (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [1:0] Counter2_Mod3CE_inst0_O;
wire and_inst0_out;
wire [1:0] coreir_const22_inst0_out;
wire coreir_eq_2_inst0_out;
wire coreir_ult2_inst0_out;
Counter2_Mod3CE Counter2_Mod3CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter2_Mod3CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult2_inst0_out), .out(and_inst0_out));
coreir_const #(.value(2'h2), .width(2)) coreir_const22_inst0(.out(coreir_const22_inst0_out));
coreir_eq #(.width(2)) coreir_eq_2_inst0(.in0(Counter2_Mod3CE_inst0_O), .in1(coreir_const22_inst0_out), .out(coreir_eq_2_inst0_out));
coreir_ult #(.width(2)) coreir_ult2_inst0(.in0(Counter2_Mod3CE_inst0_O), .in1(coreir_const22_inst0_out), .out(coreir_ult2_inst0_out));
assign valid = coreir_eq_2_inst0_out;
endmodule

module Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_unq1 (input CLK/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire InitialDelayCounter_7_inst0_valid;
wire [7:0] LUT_Array_3_Array_8_Bit__t_9n_inst0_data_0;
wire [7:0] LUT_Array_3_Array_8_Bit__t_9n_inst0_data_1;
wire [7:0] LUT_Array_3_Array_8_Bit__t_9n_inst0_data_2;
wire [0:0] coreir_const11_inst0_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(InitialDelayCounter_7_inst0_valid), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
InitialDelayCounter_7 InitialDelayCounter_7_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_7_inst0_valid));
LUT_Array_3_Array_8_Bit__t_9n LUT_Array_3_Array_8_Bit__t_9n_inst0(.CLK(CLK), .addr(Counter4_Mod9CE_inst0_O), .data_0(LUT_Array_3_Array_8_Bit__t_9n_inst0_data_0), .data_1(LUT_Array_3_Array_8_Bit__t_9n_inst0_data_1), .data_2(LUT_Array_3_Array_8_Bit__t_9n_inst0_data_2));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_3_Array_8_Bit__t_9n_inst0_data_0;
assign O_1 = LUT_Array_3_Array_8_Bit__t_9n_inst0_data_1;
assign O_2 = LUT_Array_3_Array_8_Bit__t_9n_inst0_data_2;
assign valid_down = InitialDelayCounter_7_inst0_valid;
endmodule

module Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire InitialDelayCounter_2_inst0_valid;
wire [7:0] LUT_Array_3_Array_8_Bit__t_9n_inst0_data_0;
wire [7:0] LUT_Array_3_Array_8_Bit__t_9n_inst0_data_1;
wire [7:0] LUT_Array_3_Array_8_Bit__t_9n_inst0_data_2;
wire [0:0] coreir_const11_inst0_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(InitialDelayCounter_2_inst0_valid), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
InitialDelayCounter_2 InitialDelayCounter_2_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_2_inst0_valid));
LUT_Array_3_Array_8_Bit__t_9n LUT_Array_3_Array_8_Bit__t_9n_inst0(.CLK(CLK), .addr(Counter4_Mod9CE_inst0_O), .data_0(LUT_Array_3_Array_8_Bit__t_9n_inst0_data_0), .data_1(LUT_Array_3_Array_8_Bit__t_9n_inst0_data_1), .data_2(LUT_Array_3_Array_8_Bit__t_9n_inst0_data_2));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_3_Array_8_Bit__t_9n_inst0_data_0;
assign O_1 = LUT_Array_3_Array_8_Bit__t_9n_inst0_data_1;
assign O_2 = LUT_Array_3_Array_8_Bit__t_9n_inst0_data_2;
assign valid_down = InitialDelayCounter_2_inst0_valid;
endmodule

module Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_unq1 (input CLK/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire InitialDelayCounter_11_inst0_valid;
wire [7:0] LUT_Array_1_Array_8_Bit__t_9n_inst0_data_0;
wire [0:0] coreir_const11_inst0_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(InitialDelayCounter_11_inst0_valid), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
InitialDelayCounter_11 InitialDelayCounter_11_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_11_inst0_valid));
LUT_Array_1_Array_8_Bit__t_9n LUT_Array_1_Array_8_Bit__t_9n_inst0(.CLK(CLK), .addr(Counter4_Mod9CE_inst0_O), .data_0(LUT_Array_1_Array_8_Bit__t_9n_inst0_data_0));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_1_Array_8_Bit__t_9n_inst0_data_0;
assign valid_down = InitialDelayCounter_11_inst0_valid;
endmodule

module Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [3:0] Counter4_Mod9CE_inst0_O;
wire InitialDelayCounter_6_inst0_valid;
wire [7:0] LUT_Array_1_Array_8_Bit__t_9n_inst0_data_0;
wire [0:0] coreir_const11_inst0_out;
Counter4_Mod9CE Counter4_Mod9CE_inst0(.CE(InitialDelayCounter_6_inst0_valid), .CLK(CLK), .O(Counter4_Mod9CE_inst0_O));
InitialDelayCounter_6 InitialDelayCounter_6_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_6_inst0_valid));
LUT_Array_1_Array_8_Bit__t_9n LUT_Array_1_Array_8_Bit__t_9n_inst0(.CLK(CLK), .addr(Counter4_Mod9CE_inst0_O), .data_0(LUT_Array_1_Array_8_Bit__t_9n_inst0_data_0));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_1_Array_8_Bit__t_9n_inst0_data_0;
assign valid_down = InitialDelayCounter_6_inst0_valid;
endmodule

module Add_Atom (input [7:0] I__0/*verilator public*/, input [7:0] I__1/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] coreir_add8_inst0_out;
coreir_add #(.width(8)) coreir_add8_inst0(.in0(I__0), .in1(I__1), .out(coreir_add8_inst0_out));
assign O = coreir_add8_inst0_out;
endmodule

module renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___ (input [7:0] in0/*verilator public*/, input [7:0] in1/*verilator public*/, output [7:0] out/*verilator public*/);
wire [7:0] Add_Atom_inst0_O;
Add_Atom Add_Atom_inst0(.I__0(in0), .I__1(in1), .O(Add_Atom_inst0_O));
assign out = Add_Atom_inst0_O;
endmodule

module ReduceParallel_n3_oprenamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____in0_Array_8_In_Bit___in1_Array_8_In_Bit___out_Array_8_Out_Bit___ (input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_out;
wire [7:0] renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst1_out;
renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___ renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0(.in0(I_0), .in1(renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst1_out), .out(renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_out));
renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___ renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst1(.in0(I_1), .in1(I_2), .out(renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst1_out));
assign O = renamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_out;
endmodule

module Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] ReduceParallel_n3_oprenamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____in0_Array_8_In_Bit___in1_Array_8_In_Bit___out_Array_8_Out_Bit____inst0_O;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [0:0] reg_P_inst0_out;
ReduceParallel_n3_oprenamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____in0_Array_8_In_Bit___in1_Array_8_In_Bit___out_Array_8_Out_Bit___ ReduceParallel_n3_oprenamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____in0_Array_8_In_Bit___in1_Array_8_In_Bit___out_Array_8_Out_Bit____inst0(.I_0(I_0), .I_1(I_1), .I_2(I_2), .O(ReduceParallel_n3_oprenamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____in0_Array_8_In_Bit___in1_Array_8_In_Bit___out_Array_8_Out_Bit____inst0_O));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(ReduceParallel_n3_oprenamedForReduce_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____in0_Array_8_In_Bit___in1_Array_8_In_Bit___out_Array_8_Out_Bit____inst0_O), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(valid_up), .out(reg_P_inst0_out));
assign O_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign valid_down = reg_P_inst0_out[0];
endmodule

module Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_O_0;
wire Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_valid_down;
Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___ Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_2(I_2), .O_0(Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_O_0), .valid_down(Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_valid_down), .valid_up(valid_up));
assign O_0 = Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_O_0;
assign valid_down = Reduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_valid_down;
endmodule

module NativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___ (input [7:0] I_0__0/*verilator public*/, input [7:0] I_0__1/*verilator public*/, output [7:0] O_0/*verilator public*/);
wire [7:0] Add_Atom_inst0_O;
Add_Atom Add_Atom_inst0(.I__0(I_0__0), .I__1(I_0__1), .O(Add_Atom_inst0_O));
assign O_0 = Add_Atom_inst0_O;
endmodule

module renamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit____ (input [7:0] in0_0/*verilator public*/, input [7:0] in1_0/*verilator public*/, output [7:0] out_0/*verilator public*/);
wire [7:0] NativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_O_0;
NativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit___ NativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0(.I_0__0(in0_0), .I_0__1(in1_0), .O_0(NativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_O_0));
assign out_0 = NativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____inst0_O_0;
endmodule

module ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue (input CE/*verilator public*/, input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] out_0/*verilator public*/, output ready/*verilator public*/, output valid/*verilator public*/);
wire Counter2_Mod3CE_COUT_inst0_COUT;
wire [1:0] Counter2_Mod3CE_COUT_inst0_O;
wire [7:0] Mux_Array_1_Array_8_Out_Bit___t_2n_inst0_out_0;
wire [7:0] Register_Array_1_Array_8_Out_Bit___t_0init_TrueCE_FalseRESET_inst0_O_0;
wire bit_const_1_None_out;
wire [1:0] const_0_2_out;
wire corebit_eq_inst0_O;
wire coreir_eq_2_inst0_out;
wire [7:0] renamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_out_0;
Counter2_Mod3CE_COUT Counter2_Mod3CE_COUT_inst0(.CE(CE), .CLK(CLK), .COUT(Counter2_Mod3CE_COUT_inst0_COUT), .O(Counter2_Mod3CE_COUT_inst0_O));
Mux_Array_1_Array_8_Out_Bit___t_2n Mux_Array_1_Array_8_Out_Bit___t_2n_inst0(.data_0_0(renamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_out_0), .data_1_0(I_0), .out_0(Mux_Array_1_Array_8_Out_Bit___t_2n_inst0_out_0), .sel(coreir_eq_2_inst0_out));
Register_Array_1_Array_8_Out_Bit___t_0init_TrueCE_FalseRESET Register_Array_1_Array_8_Out_Bit___t_0init_TrueCE_FalseRESET_inst0(.CE(CE), .CLK(CLK), .I_0(Mux_Array_1_Array_8_Out_Bit___t_2n_inst0_out_0), .O_0(Register_Array_1_Array_8_Out_Bit___t_0init_TrueCE_FalseRESET_inst0_O_0));
corebit_const #(.value(1)) bit_const_1_None(.out(bit_const_1_None_out));
coreir_const #(.value(2'h0), .width(2)) const_0_2(.out(const_0_2_out));
corebit_eq corebit_eq_inst0(.I0(Counter2_Mod3CE_COUT_inst0_COUT), .I1(bit_const_1_None_out), .O(corebit_eq_inst0_O));
coreir_eq #(.width(2)) coreir_eq_2_inst0(.in0(Counter2_Mod3CE_COUT_inst0_O), .in1(const_0_2_out), .out(coreir_eq_2_inst0_out));
renamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit____ renamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0(.in0_0(I_0), .in1_0(Register_Array_1_Array_8_Out_Bit___t_0init_TrueCE_FalseRESET_inst0_O_0), .out_0(renamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_out_0));
assign out_0 = renamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_out_0;
assign ready = bit_const_1_None_out;
assign valid = corebit_eq_inst0_O;
endmodule

module Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit____ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire InitialDelayCounter_3_inst0_valid;
wire NestedCounters_TSeq_3_6_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid;
wire [7:0] ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_out_0;
wire ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_ready;
wire ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_valid;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
InitialDelayCounter_3 InitialDelayCounter_3_inst0(.CE(valid_up), .CLK(CLK), .valid(InitialDelayCounter_3_inst0_valid));
NestedCounters_TSeq_3_6_SSeq_1_Int___hasCETrue_hasResetFalse NestedCounters_TSeq_3_6_SSeq_1_Int___hasCETrue_hasResetFalse_inst0(.CE(valid_up), .CLK(CLK), .valid(NestedCounters_TSeq_3_6_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid));
ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0(.CE(NestedCounters_TSeq_3_6_SSeq_1_Int___hasCETrue_hasResetFalse_inst0_valid), .CLK(CLK), .I_0(I_0), .out_0(ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_out_0), .ready(ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_ready), .valid(ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_valid));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_out_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0));
Term_Bitt Term_Bitt_inst0(.I(ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_valid));
Term_Bitt Term_Bitt_inst1(.I(ReduceSequential_n3_oprenamedForReduce_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____in0_Array_1_Array_8_In_Bit____in1_Array_1_Array_8_In_Bit____out_Array_1_Array_8_Out_Bit_____ceTrue_inst0_ready));
assign O_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign valid_down = InitialDelayCounter_3_inst0_valid;
endmodule

module Module_1 (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1;
wire Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2;
wire Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__1;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__1;
wire Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_O_0;
wire Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_valid_down;
wire and_inst0_out;
wire and_inst1_out;
Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_unq1 Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .valid_down(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_unq1 Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_2(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .valid_down(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0__0(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .I_0__1(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .O_0(Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .valid_down(Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_O_0), .I1_0(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0__0(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .O_0__1(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .valid_down(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(and_inst1_out));
Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .I_0__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .I_1__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__0), .I_1__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__1), .I_2__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__0), .I_2__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__1), .O_0(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_1(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1), .O_2(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2), .valid_down(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0(I_0), .I0_1(I_1), .I0_2(I_2), .I1_0(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I1_1(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I1_2(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_0__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .O_0__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .O_1__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__0), .O_1__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__1), .O_2__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__0), .O_2__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__1), .valid_down(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(and_inst0_out));
Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .I_1(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1), .I_2(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2), .O_0(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .valid_down(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit____ Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0(.CLK(CLK), .I_0(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_0(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_O_0), .valid_down(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_valid_down), .valid_up(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
corebit_and and_inst0(.in0(valid_up), .in1(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_valid_down), .in1(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst1_out));
assign O_0 = Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
assign valid_down = Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
endmodule

module Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Module_1_inst0_O_0;
wire Module_1_inst0_valid_down;
Module_1 Module_1_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_2(I_2), .O_0(Module_1_inst0_O_0), .valid_down(Module_1_inst0_valid_down), .valid_up(valid_up));
assign O_0 = Module_1_inst0_O_0;
assign valid_down = Module_1_inst0_valid_down;
endmodule

module Module_0 (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0;
wire [7:0] Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1;
wire Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2;
wire Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__1;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__0;
wire [7:0] Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__1;
wire Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_O_0;
wire Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_valid_down;
wire and_inst0_out;
wire and_inst1_out;
Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .valid_down(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_2(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .valid_down(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0__0(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .I_0__1(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .O_0(Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .valid_down(Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_O_0), .I1_0(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0__0(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .O_0__1(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .valid_down(Map_T_n1_i8_opNativeMapParallel_n1_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(and_inst1_out));
Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .I_0__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .I_1__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__0), .I_1__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__1), .I_2__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__0), .I_2__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__1), .O_0(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_1(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1), .O_2(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2), .valid_down(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I0_0(I_0), .I0_1(I_1), .I0_2(I_2), .I1_0(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I1_1(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I1_2(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_0__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__0), .O_0__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0__1), .O_1__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__0), .O_1__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1__1), .O_2__0(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__0), .O_2__1(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2__1), .valid_down(Map_T_n3_i6_opNativeMapParallel_n3_opatomTupleCreator_t0Int_t1Int_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Tuple_0_Array_8_Out_Bit_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(and_inst0_out));
Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .I_1(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1), .I_2(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2), .O_0(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .valid_down(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n3_i6_opNativeMapParallel_n3_opLShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_3_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit____ Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0(.CLK(CLK), .I_0(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_0(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_O_0), .valid_down(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_valid_down), .valid_up(Map_T_n3_i6_opReduce_S_n3_opAdd_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
corebit_and and_inst0(.in0(valid_up), .in1(Const_tTSeq_3_6_SSeq_3_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(Reduce_T_n3_i6_opNativeMapParallel_n1_opAdd_Atom_I_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit____O_Array_8_Out_Bit____I_Array_1_Tuple_0_Array_8_In_Bit___1_Array_8_In_Bit_____O_Array_1_Array_8_Out_Bit_____inst0_valid_down), .in1(Const_tTSeq_1_8_SSeq_1_Int___hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst1_out));
assign O_0 = Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
assign valid_down = Map_T_n1_i8_opNativeMapParallel_n1_opRShift_Atom_I_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Tuple_0_Array_8_In_Bit_1_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
endmodule

module Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_2/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Module_0_inst0_O_0;
wire Module_0_inst0_valid_down;
Module_0 Module_0_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_2(I_2), .O_0(Module_0_inst0_O_0), .valid_down(Module_0_inst0_valid_down), .valid_up(valid_up));
assign O_0 = Module_0_inst0_O_0;
assign valid_down = Module_0_inst0_valid_down;
endmodule

module top (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, output [7:0] O_0/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0;
wire FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
wire FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_1;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_1;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_1;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_1;
wire Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_2;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_2;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_0;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_1;
wire [7:0] Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_2;
wire Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down;
wire [7:0] Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0;
wire [7:0] Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1;
wire [7:0] Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2;
wire Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down;
wire [7:0] Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_0;
wire [7:0] Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_1;
wire [7:0] Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_2;
wire Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst11_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst11_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst5_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst7_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst7_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_valid_down;
wire [7:0] Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst9_O_0;
wire Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst9_valid_down;
wire [7:0] Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0;
wire Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
wire Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0;
wire Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst11_out;
wire and_inst12_out;
wire and_inst13_out;
wire and_inst14_out;
wire and_inst15_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
wire and_inst8_out;
wire and_inst9_out;
FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0(I_0), .O_0(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .valid_down(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0(Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_0(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .valid_down(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .O_0(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .valid_down(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .I1_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .valid_up(and_inst1_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .I1_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .valid_up(and_inst3_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_1), .I1_0(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down), .valid_up(and_inst6_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_1), .I1_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down), .valid_up(and_inst9_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_1), .I1_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down), .valid_up(and_inst11_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_1), .I1_0(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down), .valid_up(and_inst14_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0(.CLK(CLK), .I0_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .I1_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .valid_up(and_inst0_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1(.CLK(CLK), .I0_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .I1_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .valid_up(and_inst2_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2(.CLK(CLK), .I0_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_0), .I1_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_1), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down), .valid_up(and_inst5_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3(.CLK(CLK), .I0_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst7_O_0), .I1_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_1), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down), .valid_up(and_inst8_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4(.CLK(CLK), .I0_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst9_O_0), .I1_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_1), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down), .valid_up(and_inst10_out));
Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5(.CLK(CLK), .I0_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst11_O_0), .I1_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_O_0), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_1), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down), .valid_up(and_inst13_out));
Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2), .O_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0), .O_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1), .O_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down));
Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2), .O_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0), .O_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1), .O_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down));
Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0_2), .O_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0), .O_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_1), .O_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down));
Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0_2), .O_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0), .O_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_1), .O_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down));
Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0_2), .O_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0), .O_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_1), .O_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down));
Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0_2), .O_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0), .O_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_1), .O_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleAppender_tInt_n2_I0_Array_2_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_2_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down));
Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .I0_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2), .I0_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_0), .I0_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_1), .I0_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_2), .I1_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_0), .I1_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_1), .I1_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_O_2), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2), .O_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_0), .O_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_1), .O_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_2), .O_2_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_0), .O_2_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_1), .O_2_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .valid_up(and_inst7_out));
Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1(.CLK(CLK), .I0_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .I0_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .I0_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2), .I0_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_0), .I0_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_1), .I0_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_2), .I1_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_0), .I1_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_1), .I1_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_O_2), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2), .O_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_0), .O_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_1), .O_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_2), .O_2_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_0), .O_2_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_1), .O_2_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .valid_up(and_inst15_out));
Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0(.CLK(CLK), .I0_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0), .I0_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1), .I0_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2), .I1_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0), .I1_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1), .I1_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2), .O_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_0), .O_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_1), .O_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .valid_up(and_inst4_out));
Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock_ Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1(.CLK(CLK), .I0_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_0), .I0_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_1), .I0_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_O_2), .I1_0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_0), .I1_1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_1), .I1_2(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_O_2), .O_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .O_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .O_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2), .O_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_0), .O_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_1), .O_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_2), .valid_down(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .valid_up(and_inst12_out));
Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .I_1(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1), .I_2(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2), .O_0(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .valid_down(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_0), .I_1(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_1), .I_2(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_2), .O_0(Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .valid_down(Map_T_n16_i0_opModule_1_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_valid_down));
Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_0_2), .I_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_0), .I_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_1), .I_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_1_2), .I_2_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_0), .I_2_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_1), .I_2_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_O_2_2), .O_0(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_1(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_1), .O_2(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_2), .valid_down(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down));
Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit_ Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1(.CLK(CLK), .I_0_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_0), .I_0_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_1), .I_0_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_0_2), .I_1_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_0), .I_1_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_1), .I_1_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_1_2), .I_2_0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_0), .I_2_1(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_1), .I_2_2(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_O_2_2), .O_0(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_0), .O_1(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_1), .O_2(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_O_2), .valid_down(Map_T_n16_i0_opserialize_tSSeq_3_Int_n3_i6_hasRESETFalse_I_Array_3_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst1_valid_down), .valid_up(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleAppender_tSSeq_3_Int_n2_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_2_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_3_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10(.CLK(CLK), .I_0(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_valid_down), .valid_up(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst11(.CLK(CLK), .I_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst11_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst11_valid_down), .valid_up(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3(.CLK(CLK), .I_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down), .valid_up(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4(.CLK(CLK), .I_0(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_valid_down), .valid_up(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst5(.CLK(CLK), .I_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst5_valid_down), .valid_up(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6(.CLK(CLK), .I_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_valid_down), .valid_up(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst7(.CLK(CLK), .I_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst7_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst7_valid_down), .valid_up(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8(.CLK(CLK), .I_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_valid_down), .valid_up(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down));
Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst9(.CLK(CLK), .I_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_O_0), .O_0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst9_O_0), .valid_down(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst9_valid_down), .valid_up(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_valid_down));
Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .valid_down(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .valid_down(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_O_0), .O_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .valid_down(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down));
Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3(.CLK(CLK), .I_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_0(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .valid_down(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down), .valid_up(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down));
corebit_and and_inst0(.in0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .in1(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .in1(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst9_valid_down), .in1(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst8_valid_down), .out(and_inst10_out));
corebit_and and_inst11(.in0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down), .in1(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .out(and_inst11_out));
corebit_and and_inst12(.in0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down), .in1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst4_valid_down), .out(and_inst12_out));
corebit_and and_inst13(.in0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst11_valid_down), .in1(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst10_valid_down), .out(and_inst13_out));
corebit_and and_inst14(.in0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down), .in1(Map_T_n16_i0_opModule_0_I_Array_3_Array_8_In_Bit_O_Array_1_Array_8_Out_Bit_CLK_In_Clock_valid_up_In_Bit_valid_down_Out_Bit__inst0_valid_down), .out(and_inst14_out));
corebit_and and_inst15(.in0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .in1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst5_valid_down), .out(and_inst15_out));
corebit_and and_inst2(.in0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down), .in1(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .in1(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .in1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst1_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst5_valid_down), .in1(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst4_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down), .in1(FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(Map_T_n16_i0_opMap_T_n1_i8_opsseqTupleCreator_tSSeq_3_Int_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_3_Array_8_In_Bit_I1_Array_3_Array_8_In_Bit_O_Array_2_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst0_valid_down), .in1(Map_T_n16_i0_opMap_T_n1_i8_opRemove_1_S_opstupleToSSeq_tInt_n3_I_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I_Array_1_Array_3_Array_8_In_Bit_O_Array_3_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst2_valid_down), .out(and_inst7_out));
corebit_and and_inst8(.in0(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst7_valid_down), .in1(Shift_t_n16_i0_amt1_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst6_valid_down), .out(and_inst8_out));
corebit_and and_inst9(.in0(Map_T_n16_i0_opMap_T_n1_i8_opNativeMapParallel_n1_opsseqTupleCreator_tInt_I0_Array_8_In_Bit_I1_Array_8_In_Bit_O_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_I0_Array_1_Array_8_In_Bit_I1_Array_1_Array_8_In_Bit_O_Array_1_Array_2_Array_8_Out_Bit_valid_up_In_Bit_valid_down_Out_Bit_CLK_In_Clock__inst3_valid_down), .in1(Shift_t_n16_i0_amt4_tElTSeq_1_8_SSeq_1_Int____hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down), .out(and_inst9_out));
assign O_0 = FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
assign valid_down = FIFO_tTSeq_16_0_TSeq_1_8_SSeq_1_Int____delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
endmodule

